magic
tech sky130B
magscale 1 2
timestamp 1668205333
<< viali >>
rect 1961 57545 1995 57579
rect 3893 57545 3927 57579
rect 5089 57545 5123 57579
rect 6653 57545 6687 57579
rect 8217 57545 8251 57579
rect 9781 57545 9815 57579
rect 11621 57545 11655 57579
rect 12909 57545 12943 57579
rect 14473 57545 14507 57579
rect 16773 57545 16807 57579
rect 17693 57545 17727 57579
rect 19441 57545 19475 57579
rect 20821 57545 20855 57579
rect 22385 57545 22419 57579
rect 24593 57545 24627 57579
rect 25513 57545 25547 57579
rect 27169 57545 27203 57579
rect 28641 57545 28675 57579
rect 30205 57545 30239 57579
rect 32321 57545 32355 57579
rect 33333 57545 33367 57579
rect 34897 57545 34931 57579
rect 36461 57545 36495 57579
rect 38025 57545 38059 57579
rect 40049 57545 40083 57579
rect 41153 57545 41187 57579
rect 42717 57545 42751 57579
rect 44281 57545 44315 57579
rect 45845 57545 45879 57579
rect 47777 57545 47811 57579
rect 2145 57409 2179 57443
rect 4077 57409 4111 57443
rect 5273 57409 5307 57443
rect 6837 57409 6871 57443
rect 8401 57409 8435 57443
rect 9965 57409 9999 57443
rect 11805 57409 11839 57443
rect 13093 57409 13127 57443
rect 14657 57409 14691 57443
rect 16957 57409 16991 57443
rect 17509 57409 17543 57443
rect 19257 57409 19291 57443
rect 20637 57409 20671 57443
rect 22201 57409 22235 57443
rect 24409 57409 24443 57443
rect 25329 57409 25363 57443
rect 26985 57409 27019 57443
rect 28457 57409 28491 57443
rect 30021 57409 30055 57443
rect 32137 57409 32171 57443
rect 33149 57409 33183 57443
rect 34713 57409 34747 57443
rect 36277 57409 36311 57443
rect 37841 57409 37875 57443
rect 39865 57409 39899 57443
rect 40969 57409 41003 57443
rect 42533 57409 42567 57443
rect 44097 57409 44131 57443
rect 45661 57409 45695 57443
rect 47593 57409 47627 57443
rect 48789 57409 48823 57443
rect 50353 57409 50387 57443
rect 51917 57409 51951 57443
rect 53481 57409 53515 57443
rect 56609 57409 56643 57443
rect 57989 57409 58023 57443
rect 55321 57341 55355 57375
rect 2697 57205 2731 57239
rect 18613 57205 18647 57239
rect 20085 57205 20119 57239
rect 18337 57001 18371 57035
rect 19257 57001 19291 57035
rect 57529 57001 57563 57035
rect 18521 56797 18555 56831
rect 19441 56797 19475 56831
rect 25881 56797 25915 56831
rect 58173 56797 58207 56831
rect 17877 56661 17911 56695
rect 20085 56661 20119 56695
rect 20729 56661 20763 56695
rect 22293 56661 22327 56695
rect 25329 56661 25363 56695
rect 26065 56661 26099 56695
rect 26617 56661 26651 56695
rect 42349 56661 42383 56695
rect 13553 56457 13587 56491
rect 15945 56457 15979 56491
rect 17417 56457 17451 56491
rect 17877 56457 17911 56491
rect 18521 56457 18555 56491
rect 19349 56457 19383 56491
rect 19809 56457 19843 56491
rect 21281 56457 21315 56491
rect 22845 56457 22879 56491
rect 26433 56457 26467 56491
rect 27353 56457 27387 56491
rect 29837 56457 29871 56491
rect 32321 56457 32355 56491
rect 34161 56457 34195 56491
rect 36001 56457 36035 56491
rect 45109 56457 45143 56491
rect 45753 56457 45787 56491
rect 13737 56321 13771 56355
rect 16129 56321 16163 56355
rect 16773 56321 16807 56355
rect 17233 56321 17267 56355
rect 18061 56321 18095 56355
rect 18705 56321 18739 56355
rect 19165 56321 19199 56355
rect 19993 56321 20027 56355
rect 20637 56321 20671 56355
rect 21097 56321 21131 56355
rect 22017 56321 22051 56355
rect 22661 56321 22695 56355
rect 23489 56321 23523 56355
rect 23949 56321 23983 56355
rect 24961 56321 24995 56355
rect 25605 56321 25639 56355
rect 26249 56321 26283 56355
rect 27169 56321 27203 56355
rect 27813 56321 27847 56355
rect 29653 56321 29687 56355
rect 30297 56321 30331 56355
rect 30941 56321 30975 56355
rect 31401 56321 31435 56355
rect 32137 56321 32171 56355
rect 32781 56321 32815 56355
rect 33977 56321 34011 56355
rect 34621 56321 34655 56355
rect 35817 56321 35851 56355
rect 36461 56321 36495 56355
rect 44925 56321 44959 56355
rect 45569 56321 45603 56355
rect 46213 56321 46247 56355
rect 58173 56321 58207 56355
rect 20453 56185 20487 56219
rect 22201 56185 22235 56219
rect 24133 56185 24167 56219
rect 25789 56185 25823 56219
rect 14289 56117 14323 56151
rect 25145 56117 25179 56151
rect 31585 56117 31619 56151
rect 44373 56117 44407 56151
rect 16865 55913 16899 55947
rect 18705 55913 18739 55947
rect 19717 55913 19751 55947
rect 26433 55845 26467 55879
rect 20913 55777 20947 55811
rect 17049 55709 17083 55743
rect 18521 55709 18555 55743
rect 19901 55709 19935 55743
rect 26249 55709 26283 55743
rect 26893 55709 26927 55743
rect 16221 55573 16255 55607
rect 18061 55573 18095 55607
rect 20361 55573 20395 55607
rect 22569 55573 22603 55607
rect 24869 55573 24903 55607
rect 25513 55573 25547 55607
rect 19533 55369 19567 55403
rect 17141 55301 17175 55335
rect 18981 55301 19015 55335
rect 58173 55097 58207 55131
rect 58173 53941 58207 53975
rect 58173 52445 58207 52479
rect 58173 51357 58207 51391
rect 58173 49725 58207 49759
rect 58173 48501 58207 48535
rect 58173 47005 58207 47039
rect 58173 45917 58207 45951
rect 58173 44217 58207 44251
rect 58173 43061 58207 43095
rect 13093 42245 13127 42279
rect 12909 42177 12943 42211
rect 14933 42177 14967 42211
rect 15117 42177 15151 42211
rect 13277 41973 13311 42007
rect 15301 41973 15335 42007
rect 15025 41633 15059 41667
rect 13185 41565 13219 41599
rect 13277 41565 13311 41599
rect 13369 41565 13403 41599
rect 13553 41565 13587 41599
rect 14657 41565 14691 41599
rect 15485 41565 15519 41599
rect 15669 41565 15703 41599
rect 15761 41565 15795 41599
rect 15899 41565 15933 41599
rect 16681 41565 16715 41599
rect 58173 41565 58207 41599
rect 12265 41497 12299 41531
rect 12449 41497 12483 41531
rect 14841 41497 14875 41531
rect 16129 41497 16163 41531
rect 19257 41497 19291 41531
rect 19441 41497 19475 41531
rect 12081 41429 12115 41463
rect 12909 41429 12943 41463
rect 14197 41429 14231 41463
rect 19625 41429 19659 41463
rect 20177 41429 20211 41463
rect 23581 41429 23615 41463
rect 21189 41225 21223 41259
rect 16681 41157 16715 41191
rect 19380 41157 19414 41191
rect 20085 41157 20119 41191
rect 21833 41157 21867 41191
rect 9873 41089 9907 41123
rect 9978 41095 10012 41129
rect 10078 41089 10112 41123
rect 10241 41089 10275 41123
rect 13093 41089 13127 41123
rect 13185 41089 13219 41123
rect 13277 41089 13311 41123
rect 13461 41089 13495 41123
rect 15393 41089 15427 41123
rect 15556 41089 15590 41123
rect 15656 41092 15690 41126
rect 15761 41089 15795 41123
rect 19625 41089 19659 41123
rect 20361 41089 20395 41123
rect 20466 41095 20500 41129
rect 20566 41089 20600 41123
rect 20729 41089 20763 41123
rect 22017 41089 22051 41123
rect 22845 41089 22879 41123
rect 23029 41089 23063 41123
rect 23121 41089 23155 41123
rect 23259 41089 23293 41123
rect 10793 40953 10827 40987
rect 13921 40953 13955 40987
rect 16037 40953 16071 40987
rect 23949 40953 23983 40987
rect 9597 40885 9631 40919
rect 12817 40885 12851 40919
rect 18245 40885 18279 40919
rect 22201 40885 22235 40919
rect 23489 40885 23523 40919
rect 11529 40681 11563 40715
rect 18705 40681 18739 40715
rect 24777 40681 24811 40715
rect 5181 40477 5215 40511
rect 10149 40477 10183 40511
rect 10416 40477 10450 40511
rect 11989 40477 12023 40511
rect 12256 40477 12290 40511
rect 14473 40477 14507 40511
rect 17417 40477 17451 40511
rect 18521 40477 18555 40511
rect 19257 40477 19291 40511
rect 19441 40477 19475 40511
rect 19533 40477 19567 40511
rect 19625 40477 19659 40511
rect 20821 40477 20855 40511
rect 22937 40477 22971 40511
rect 23121 40477 23155 40511
rect 23216 40477 23250 40511
rect 23325 40477 23359 40511
rect 30941 40477 30975 40511
rect 58173 40477 58207 40511
rect 5448 40409 5482 40443
rect 14289 40409 14323 40443
rect 17150 40409 17184 40443
rect 18337 40409 18371 40443
rect 21088 40409 21122 40443
rect 24409 40409 24443 40443
rect 24593 40409 24627 40443
rect 31186 40409 31220 40443
rect 6561 40341 6595 40375
rect 7205 40341 7239 40375
rect 13369 40341 13403 40375
rect 14657 40341 14691 40375
rect 16037 40341 16071 40375
rect 19901 40341 19935 40375
rect 22201 40341 22235 40375
rect 23581 40341 23615 40375
rect 32321 40341 32355 40375
rect 3893 40137 3927 40171
rect 10701 40137 10735 40171
rect 14013 40137 14047 40171
rect 21189 40137 21223 40171
rect 21833 40137 21867 40171
rect 22937 40137 22971 40171
rect 25237 40137 25271 40171
rect 28733 40137 28767 40171
rect 4537 40069 4571 40103
rect 20085 40069 20119 40103
rect 23305 40069 23339 40103
rect 24102 40069 24136 40103
rect 2780 40001 2814 40035
rect 4721 40001 4755 40035
rect 6607 40001 6641 40035
rect 6742 40001 6776 40035
rect 6842 40001 6876 40035
rect 7021 40001 7055 40035
rect 7481 40001 7515 40035
rect 7748 40001 7782 40035
rect 9321 40001 9355 40035
rect 9588 40001 9622 40035
rect 11529 40001 11563 40035
rect 11692 40001 11726 40035
rect 11805 40001 11839 40035
rect 11943 40001 11977 40035
rect 15126 40001 15160 40035
rect 22089 40001 22123 40035
rect 22182 40001 22216 40035
rect 22293 40001 22327 40035
rect 22477 40001 22511 40035
rect 23121 40001 23155 40035
rect 27620 40001 27654 40035
rect 2513 39933 2547 39967
rect 15393 39933 15427 39967
rect 18337 39933 18371 39967
rect 23857 39933 23891 39967
rect 27353 39933 27387 39967
rect 5825 39865 5859 39899
rect 20637 39865 20671 39899
rect 4353 39797 4387 39831
rect 5273 39797 5307 39831
rect 6377 39797 6411 39831
rect 8861 39797 8895 39831
rect 12173 39797 12207 39831
rect 12633 39797 12667 39831
rect 17785 39797 17819 39831
rect 3801 39593 3835 39627
rect 5641 39593 5675 39627
rect 11529 39593 11563 39627
rect 14473 39593 14507 39627
rect 19257 39593 19291 39627
rect 30849 39593 30883 39627
rect 6101 39457 6135 39491
rect 13001 39457 13035 39491
rect 32321 39457 32355 39491
rect 4077 39389 4111 39423
rect 4169 39389 4203 39423
rect 4261 39389 4295 39423
rect 4445 39389 4479 39423
rect 4997 39389 5031 39423
rect 5181 39389 5215 39423
rect 5273 39389 5307 39423
rect 5365 39389 5399 39423
rect 6368 39389 6402 39423
rect 9321 39389 9355 39423
rect 12725 39389 12759 39423
rect 14703 39389 14737 39423
rect 14841 39389 14875 39423
rect 14933 39386 14967 39420
rect 15117 39389 15151 39423
rect 18061 39389 18095 39423
rect 20637 39389 20671 39423
rect 24409 39389 24443 39423
rect 27169 39389 27203 39423
rect 31125 39389 31159 39423
rect 31214 39386 31248 39420
rect 31330 39389 31364 39423
rect 31493 39389 31527 39423
rect 9588 39321 9622 39355
rect 11161 39321 11195 39355
rect 11345 39321 11379 39355
rect 17794 39321 17828 39355
rect 20370 39321 20404 39355
rect 24654 39321 24688 39355
rect 27414 39321 27448 39355
rect 31953 39321 31987 39355
rect 32137 39321 32171 39355
rect 7481 39253 7515 39287
rect 10701 39253 10735 39287
rect 12265 39253 12299 39287
rect 15577 39253 15611 39287
rect 16681 39253 16715 39287
rect 18705 39253 18739 39287
rect 25789 39253 25823 39287
rect 28549 39253 28583 39287
rect 29745 39253 29779 39287
rect 30389 39253 30423 39287
rect 6929 39049 6963 39083
rect 7113 38981 7147 39015
rect 3545 38913 3579 38947
rect 4997 38913 5031 38947
rect 6469 38913 6503 38947
rect 7297 38913 7331 38947
rect 9045 38913 9079 38947
rect 13829 38913 13863 38947
rect 27905 38913 27939 38947
rect 30369 38913 30403 38947
rect 3801 38845 3835 38879
rect 5273 38845 5307 38879
rect 13553 38845 13587 38879
rect 30113 38845 30147 38879
rect 58173 38777 58207 38811
rect 2421 38709 2455 38743
rect 4261 38709 4295 38743
rect 10333 38709 10367 38743
rect 11621 38709 11655 38743
rect 29193 38709 29227 38743
rect 31493 38709 31527 38743
rect 6377 38505 6411 38539
rect 10057 38505 10091 38539
rect 12541 38505 12575 38539
rect 27261 38505 27295 38539
rect 28365 38505 28399 38539
rect 9597 38437 9631 38471
rect 8125 38369 8159 38403
rect 11161 38369 11195 38403
rect 20637 38369 20671 38403
rect 32229 38369 32263 38403
rect 32689 38369 32723 38403
rect 2145 38301 2179 38335
rect 2881 38301 2915 38335
rect 2973 38301 3007 38335
rect 3065 38301 3099 38335
rect 3249 38301 3283 38335
rect 6561 38301 6595 38335
rect 8401 38301 8435 38335
rect 9413 38301 9447 38335
rect 10287 38301 10321 38335
rect 10406 38301 10440 38335
rect 10538 38298 10572 38332
rect 10713 38301 10747 38335
rect 11345 38301 11379 38335
rect 12357 38301 12391 38335
rect 13001 38301 13035 38335
rect 13369 38301 13403 38335
rect 27537 38301 27571 38335
rect 27629 38301 27663 38335
rect 27721 38301 27755 38335
rect 27905 38301 27939 38335
rect 28641 38301 28675 38335
rect 28733 38301 28767 38335
rect 28825 38301 28859 38335
rect 29009 38301 29043 38335
rect 30021 38301 30055 38335
rect 1961 38233 1995 38267
rect 5917 38233 5951 38267
rect 6745 38233 6779 38267
rect 9229 38233 9263 38267
rect 11529 38233 11563 38267
rect 13185 38233 13219 38267
rect 13277 38233 13311 38267
rect 20370 38233 20404 38267
rect 30205 38233 30239 38267
rect 31962 38233 31996 38267
rect 32956 38233 32990 38267
rect 1777 38165 1811 38199
rect 2605 38165 2639 38199
rect 4629 38165 4663 38199
rect 13553 38165 13587 38199
rect 19257 38165 19291 38199
rect 26801 38165 26835 38199
rect 30389 38165 30423 38199
rect 30849 38165 30883 38199
rect 34069 38165 34103 38199
rect 4261 37961 4295 37995
rect 5365 37961 5399 37995
rect 9137 37961 9171 37995
rect 10793 37961 10827 37995
rect 13737 37961 13771 37995
rect 28089 37961 28123 37995
rect 28917 37961 28951 37995
rect 29929 37961 29963 37995
rect 31033 37961 31067 37995
rect 33057 37961 33091 37995
rect 5733 37893 5767 37927
rect 11805 37893 11839 37927
rect 13369 37893 13403 37927
rect 13461 37893 13495 37927
rect 19165 37893 19199 37927
rect 19257 37893 19291 37927
rect 26065 37893 26099 37927
rect 28273 37893 28307 37927
rect 29285 37893 29319 37927
rect 2421 37825 2455 37859
rect 2688 37825 2722 37859
rect 4537 37825 4571 37859
rect 4629 37825 4663 37859
rect 4721 37825 4755 37859
rect 4905 37825 4939 37859
rect 5549 37825 5583 37859
rect 9321 37825 9355 37859
rect 11529 37825 11563 37859
rect 11713 37825 11747 37859
rect 11897 37825 11931 37859
rect 13185 37825 13219 37859
rect 13553 37825 13587 37859
rect 17141 37825 17175 37859
rect 17234 37825 17268 37859
rect 17417 37825 17451 37859
rect 17509 37825 17543 37859
rect 17647 37825 17681 37859
rect 18889 37825 18923 37859
rect 19037 37825 19071 37859
rect 19354 37825 19388 37859
rect 19993 37825 20027 37859
rect 20177 37825 20211 37859
rect 20269 37825 20303 37859
rect 20361 37825 20395 37859
rect 21097 37825 21131 37859
rect 24225 37825 24259 37859
rect 24492 37825 24526 37859
rect 28457 37825 28491 37859
rect 29101 37825 29135 37859
rect 30389 37825 30423 37859
rect 30568 37825 30602 37859
rect 30665 37828 30699 37862
rect 30777 37825 30811 37859
rect 32413 37825 32447 37859
rect 32597 37825 32631 37859
rect 32689 37825 32723 37859
rect 32781 37825 32815 37859
rect 34345 37825 34379 37859
rect 34529 37825 34563 37859
rect 34621 37825 34655 37859
rect 34713 37825 34747 37859
rect 6469 37689 6503 37723
rect 19533 37689 19567 37723
rect 3801 37621 3835 37655
rect 12081 37621 12115 37655
rect 17785 37621 17819 37655
rect 20637 37621 20671 37655
rect 22569 37621 22603 37655
rect 23121 37621 23155 37655
rect 25605 37621 25639 37655
rect 31493 37621 31527 37655
rect 33885 37621 33919 37655
rect 34989 37621 35023 37655
rect 58173 37621 58207 37655
rect 20177 37417 20211 37451
rect 26249 37417 26283 37451
rect 33701 37417 33735 37451
rect 5089 37281 5123 37315
rect 13369 37281 13403 37315
rect 6009 37213 6043 37247
rect 7849 37213 7883 37247
rect 8125 37213 8159 37247
rect 8217 37213 8251 37247
rect 15669 37213 15703 37247
rect 18061 37213 18095 37247
rect 18154 37213 18188 37247
rect 18526 37213 18560 37247
rect 19993 37213 20027 37247
rect 21750 37213 21784 37247
rect 22017 37213 22051 37247
rect 22937 37213 22971 37247
rect 23305 37213 23339 37247
rect 24409 37213 24443 37247
rect 26525 37213 26559 37247
rect 26617 37213 26651 37247
rect 26709 37213 26743 37247
rect 26893 37213 26927 37247
rect 27353 37213 27387 37247
rect 35081 37213 35115 37247
rect 35348 37213 35382 37247
rect 6276 37145 6310 37179
rect 8033 37145 8067 37179
rect 13185 37145 13219 37179
rect 15936 37145 15970 37179
rect 18337 37145 18371 37179
rect 18429 37145 18463 37179
rect 19809 37145 19843 37179
rect 23029 37145 23063 37179
rect 23121 37145 23155 37179
rect 24676 37145 24710 37179
rect 31953 37145 31987 37179
rect 32413 37145 32447 37179
rect 7389 37077 7423 37111
rect 8401 37077 8435 37111
rect 11713 37077 11747 37111
rect 12633 37077 12667 37111
rect 17049 37077 17083 37111
rect 18705 37077 18739 37111
rect 20637 37077 20671 37111
rect 22753 37077 22787 37111
rect 25789 37077 25823 37111
rect 28181 37077 28215 37111
rect 29653 37077 29687 37111
rect 36461 37077 36495 37111
rect 12173 36873 12207 36907
rect 15485 36873 15519 36907
rect 16681 36873 16715 36907
rect 18429 36873 18463 36907
rect 30113 36873 30147 36907
rect 32873 36873 32907 36907
rect 35725 36873 35759 36907
rect 6929 36805 6963 36839
rect 7849 36805 7883 36839
rect 19073 36805 19107 36839
rect 23857 36805 23891 36839
rect 25605 36805 25639 36839
rect 27077 36805 27111 36839
rect 33057 36805 33091 36839
rect 6653 36737 6687 36771
rect 6837 36737 6871 36771
rect 7021 36737 7055 36771
rect 8033 36737 8067 36771
rect 12081 36737 12115 36771
rect 14105 36737 14139 36771
rect 14372 36737 14406 36771
rect 16957 36737 16991 36771
rect 17049 36737 17083 36771
rect 17141 36737 17175 36771
rect 17325 36737 17359 36771
rect 17785 36737 17819 36771
rect 17969 36737 18003 36771
rect 18061 36737 18095 36771
rect 18153 36737 18187 36771
rect 18889 36737 18923 36771
rect 22293 36737 22327 36771
rect 22385 36737 22419 36771
rect 22477 36737 22511 36771
rect 22661 36737 22695 36771
rect 26065 36737 26099 36771
rect 26249 36737 26283 36771
rect 27629 36737 27663 36771
rect 27885 36737 27919 36771
rect 29469 36737 29503 36771
rect 29653 36737 29687 36771
rect 29745 36737 29779 36771
rect 29837 36737 29871 36771
rect 31309 36737 31343 36771
rect 33241 36737 33275 36771
rect 34253 36737 34287 36771
rect 34416 36737 34450 36771
rect 34529 36737 34563 36771
rect 34641 36737 34675 36771
rect 35357 36737 35391 36771
rect 35541 36737 35575 36771
rect 13277 36669 13311 36703
rect 13553 36669 13587 36703
rect 19257 36669 19291 36703
rect 31585 36669 31619 36703
rect 7205 36533 7239 36567
rect 7665 36533 7699 36567
rect 19809 36533 19843 36567
rect 22109 36533 22143 36567
rect 23121 36533 23155 36567
rect 26433 36533 26467 36567
rect 29009 36533 29043 36567
rect 33701 36533 33735 36567
rect 34897 36533 34931 36567
rect 5181 36329 5215 36363
rect 7021 36329 7055 36363
rect 9505 36329 9539 36363
rect 13093 36329 13127 36363
rect 14749 36329 14783 36363
rect 16681 36329 16715 36363
rect 18521 36329 18555 36363
rect 24593 36329 24627 36363
rect 26065 36329 26099 36363
rect 27721 36329 27755 36363
rect 29561 36329 29595 36363
rect 34161 36329 34195 36363
rect 34805 36193 34839 36227
rect 3801 36125 3835 36159
rect 7251 36125 7285 36159
rect 7389 36125 7423 36159
rect 7486 36125 7520 36159
rect 7665 36125 7699 36159
rect 9321 36125 9355 36159
rect 9965 36125 9999 36159
rect 14105 36125 14139 36159
rect 14289 36125 14323 36159
rect 14381 36125 14415 36159
rect 14519 36125 14553 36159
rect 15393 36125 15427 36159
rect 16497 36125 16531 36159
rect 24823 36125 24857 36159
rect 24961 36125 24995 36159
rect 25053 36125 25087 36159
rect 25237 36125 25271 36159
rect 25881 36125 25915 36159
rect 27997 36125 28031 36159
rect 28089 36125 28123 36159
rect 28181 36125 28215 36159
rect 28365 36125 28399 36159
rect 29745 36125 29779 36159
rect 31861 36125 31895 36159
rect 32137 36125 32171 36159
rect 33793 36125 33827 36159
rect 35061 36125 35095 36159
rect 58173 36125 58207 36159
rect 4068 36057 4102 36091
rect 10232 36057 10266 36091
rect 11805 36057 11839 36091
rect 15209 36057 15243 36091
rect 15577 36057 15611 36091
rect 16313 36057 16347 36091
rect 25697 36057 25731 36091
rect 28917 36057 28951 36091
rect 29929 36057 29963 36091
rect 33977 36057 34011 36091
rect 6561 35989 6595 36023
rect 11345 35989 11379 36023
rect 17509 35989 17543 36023
rect 22569 35989 22603 36023
rect 23029 35989 23063 36023
rect 27169 35989 27203 36023
rect 30665 35989 30699 36023
rect 31309 35989 31343 36023
rect 36185 35989 36219 36023
rect 13921 35785 13955 35819
rect 27353 35785 27387 35819
rect 28365 35785 28399 35819
rect 4629 35717 4663 35751
rect 11529 35717 11563 35751
rect 14933 35717 14967 35751
rect 18245 35717 18279 35751
rect 23213 35717 23247 35751
rect 28549 35717 28583 35751
rect 4445 35649 4479 35683
rect 7490 35649 7524 35683
rect 7757 35649 7791 35683
rect 9965 35649 9999 35683
rect 10241 35649 10275 35683
rect 11713 35649 11747 35683
rect 13093 35649 13127 35683
rect 18061 35649 18095 35683
rect 23029 35649 23063 35683
rect 23121 35649 23155 35683
rect 23397 35649 23431 35683
rect 28733 35649 28767 35683
rect 30297 35649 30331 35683
rect 30460 35649 30494 35683
rect 30573 35649 30607 35683
rect 30665 35649 30699 35683
rect 8769 35581 8803 35615
rect 9045 35581 9079 35615
rect 13369 35581 13403 35615
rect 29745 35513 29779 35547
rect 4813 35445 4847 35479
rect 6377 35445 6411 35479
rect 11897 35445 11931 35479
rect 17877 35445 17911 35479
rect 22385 35445 22419 35479
rect 22845 35445 22879 35479
rect 24409 35445 24443 35479
rect 25421 35445 25455 35479
rect 30941 35445 30975 35479
rect 4353 35241 4387 35275
rect 7297 35241 7331 35275
rect 18705 35241 18739 35275
rect 30297 35241 30331 35275
rect 9045 35173 9079 35207
rect 25697 35173 25731 35207
rect 6837 35105 6871 35139
rect 9781 35105 9815 35139
rect 32137 35105 32171 35139
rect 4629 35037 4663 35071
rect 4721 35037 4755 35071
rect 4813 35037 4847 35071
rect 4997 35037 5031 35071
rect 7573 35037 7607 35071
rect 7665 35037 7699 35071
rect 7757 35037 7791 35071
rect 7941 35037 7975 35071
rect 9505 35037 9539 35071
rect 10793 35037 10827 35071
rect 10977 35037 11011 35071
rect 11069 35037 11103 35071
rect 11161 35037 11195 35071
rect 12541 35037 12575 35071
rect 12817 35037 12851 35071
rect 12909 35037 12943 35071
rect 17325 35037 17359 35071
rect 21005 35037 21039 35071
rect 21833 35037 21867 35071
rect 21925 35037 21959 35071
rect 22017 35037 22051 35071
rect 22201 35037 22235 35071
rect 24961 35037 24995 35071
rect 27077 35037 27111 35071
rect 31870 35037 31904 35071
rect 58173 35037 58207 35071
rect 6469 34969 6503 35003
rect 6653 34969 6687 35003
rect 11897 34969 11931 35003
rect 12725 34969 12759 35003
rect 17592 34969 17626 35003
rect 24777 34969 24811 35003
rect 26810 34969 26844 35003
rect 29929 34969 29963 35003
rect 30113 34969 30147 35003
rect 5549 34901 5583 34935
rect 11437 34901 11471 34935
rect 13093 34901 13127 34935
rect 19717 34901 19751 34935
rect 21557 34901 21591 34935
rect 25145 34901 25179 34935
rect 30757 34901 30791 34935
rect 3893 34697 3927 34731
rect 8769 34697 8803 34731
rect 10333 34697 10367 34731
rect 12909 34697 12943 34731
rect 16957 34697 16991 34731
rect 17509 34697 17543 34731
rect 19441 34697 19475 34731
rect 25513 34697 25547 34731
rect 32321 34697 32355 34731
rect 4537 34629 4571 34663
rect 8401 34629 8435 34663
rect 13553 34629 13587 34663
rect 13645 34629 13679 34663
rect 19073 34629 19107 34663
rect 19165 34629 19199 34663
rect 22078 34629 22112 34663
rect 34529 34629 34563 34663
rect 2513 34561 2547 34595
rect 2780 34561 2814 34595
rect 4721 34561 4755 34595
rect 8125 34561 8159 34595
rect 8218 34561 8252 34595
rect 8490 34561 8524 34595
rect 8631 34561 8665 34595
rect 9781 34561 9815 34595
rect 10563 34561 10597 34595
rect 10698 34567 10732 34601
rect 10798 34561 10832 34595
rect 10977 34561 11011 34595
rect 11785 34561 11819 34595
rect 13369 34561 13403 34595
rect 13737 34561 13771 34595
rect 17739 34561 17773 34595
rect 17877 34561 17911 34595
rect 17969 34561 18003 34595
rect 18153 34561 18187 34595
rect 18797 34561 18831 34595
rect 18890 34561 18924 34595
rect 19262 34561 19296 34595
rect 19901 34561 19935 34595
rect 20085 34561 20119 34595
rect 20177 34561 20211 34595
rect 20269 34561 20303 34595
rect 21005 34561 21039 34595
rect 21833 34561 21867 34595
rect 24869 34561 24903 34595
rect 25053 34561 25087 34595
rect 25145 34561 25179 34595
rect 25237 34561 25271 34595
rect 25973 34561 26007 34595
rect 31125 34561 31159 34595
rect 32137 34561 32171 34595
rect 7665 34493 7699 34527
rect 11529 34493 11563 34527
rect 20545 34493 20579 34527
rect 29745 34493 29779 34527
rect 30849 34493 30883 34527
rect 13921 34425 13955 34459
rect 4353 34357 4387 34391
rect 9689 34357 9723 34391
rect 23213 34357 23247 34391
rect 2605 34153 2639 34187
rect 9413 34153 9447 34187
rect 10977 34153 11011 34187
rect 11437 34153 11471 34187
rect 11989 34153 12023 34187
rect 15025 34153 15059 34187
rect 20085 34153 20119 34187
rect 22569 34153 22603 34187
rect 27169 34153 27203 34187
rect 14105 34085 14139 34119
rect 20729 34085 20763 34119
rect 5549 34017 5583 34051
rect 16957 34017 16991 34051
rect 30665 34017 30699 34051
rect 2881 33949 2915 33983
rect 2973 33949 3007 33983
rect 3065 33949 3099 33983
rect 3249 33949 3283 33983
rect 4077 33949 4111 33983
rect 4169 33949 4203 33983
rect 4261 33949 4295 33983
rect 4445 33949 4479 33983
rect 10793 33949 10827 33983
rect 14289 33949 14323 33983
rect 17693 33949 17727 33983
rect 17785 33949 17819 33983
rect 17877 33949 17911 33983
rect 18061 33949 18095 33983
rect 19717 33949 19751 33983
rect 19901 33949 19935 33983
rect 21842 33949 21876 33983
rect 22109 33949 22143 33983
rect 24409 33949 24443 33983
rect 24593 33949 24627 33983
rect 24685 33949 24719 33983
rect 24777 33949 24811 33983
rect 27629 33949 27663 33983
rect 29837 33949 29871 33983
rect 30941 33949 30975 33983
rect 31953 33949 31987 33983
rect 33793 33949 33827 33983
rect 33977 33949 34011 33983
rect 34713 33949 34747 33983
rect 34876 33949 34910 33983
rect 34976 33946 35010 33980
rect 35127 33949 35161 33983
rect 2145 33881 2179 33915
rect 4905 33881 4939 33915
rect 9505 33881 9539 33915
rect 10609 33881 10643 33915
rect 14933 33881 14967 33915
rect 16712 33881 16746 33915
rect 17417 33881 17451 33915
rect 22753 33881 22787 33915
rect 22937 33881 22971 33915
rect 23857 33881 23891 33915
rect 27874 33881 27908 33915
rect 30021 33881 30055 33915
rect 32220 33881 32254 33915
rect 34161 33881 34195 33915
rect 3801 33813 3835 33847
rect 15577 33813 15611 33847
rect 25053 33813 25087 33847
rect 29009 33813 29043 33847
rect 30205 33813 30239 33847
rect 33333 33813 33367 33847
rect 35357 33813 35391 33847
rect 4353 33609 4387 33643
rect 8217 33609 8251 33643
rect 17049 33609 17083 33643
rect 19073 33609 19107 33643
rect 27721 33609 27755 33643
rect 12725 33541 12759 33575
rect 16865 33541 16899 33575
rect 17509 33541 17543 33575
rect 18337 33541 18371 33575
rect 23581 33541 23615 33575
rect 23949 33541 23983 33575
rect 29193 33541 29227 33575
rect 34529 33541 34563 33575
rect 36102 33541 36136 33575
rect 2780 33473 2814 33507
rect 4537 33473 4571 33507
rect 4721 33473 4755 33507
rect 6837 33473 6871 33507
rect 7093 33473 7127 33507
rect 12909 33473 12943 33507
rect 16681 33473 16715 33507
rect 18521 33473 18555 33507
rect 19165 33473 19199 33507
rect 23765 33473 23799 33507
rect 24409 33473 24443 33507
rect 24593 33473 24627 33507
rect 24685 33473 24719 33507
rect 24777 33473 24811 33507
rect 27997 33473 28031 33507
rect 28089 33473 28123 33507
rect 28181 33473 28215 33507
rect 28365 33473 28399 33507
rect 29009 33473 29043 33507
rect 30297 33473 30331 33507
rect 30476 33473 30510 33507
rect 30576 33479 30610 33513
rect 30665 33473 30699 33507
rect 33885 33473 33919 33507
rect 34069 33473 34103 33507
rect 34161 33473 34195 33507
rect 34253 33473 34287 33507
rect 36369 33473 36403 33507
rect 2513 33405 2547 33439
rect 14565 33405 14599 33439
rect 14841 33405 14875 33439
rect 18153 33405 18187 33439
rect 25605 33405 25639 33439
rect 28825 33405 28859 33439
rect 32413 33405 32447 33439
rect 32689 33405 32723 33439
rect 3893 33337 3927 33371
rect 25053 33337 25087 33371
rect 58173 33337 58207 33371
rect 19717 33269 19751 33303
rect 27169 33269 27203 33303
rect 29745 33269 29779 33303
rect 30941 33269 30975 33303
rect 34989 33269 35023 33303
rect 6837 33065 6871 33099
rect 23857 33065 23891 33099
rect 25145 33065 25179 33099
rect 29561 33065 29595 33099
rect 31953 33065 31987 33099
rect 34161 33065 34195 33099
rect 34897 33065 34931 33099
rect 18429 32997 18463 33031
rect 19809 32997 19843 33031
rect 33333 32929 33367 32963
rect 7113 32861 7147 32895
rect 7205 32861 7239 32895
rect 7297 32861 7331 32895
rect 7481 32861 7515 32895
rect 8125 32861 8159 32895
rect 14105 32861 14139 32895
rect 16221 32861 16255 32895
rect 16314 32861 16348 32895
rect 16497 32861 16531 32895
rect 16686 32861 16720 32895
rect 17325 32861 17359 32895
rect 17488 32861 17522 32895
rect 17588 32861 17622 32895
rect 17693 32861 17727 32895
rect 23489 32861 23523 32895
rect 26258 32861 26292 32895
rect 26525 32861 26559 32895
rect 29745 32861 29779 32895
rect 29837 32861 29871 32895
rect 30113 32861 30147 32895
rect 32229 32861 32263 32895
rect 32321 32861 32355 32895
rect 32413 32861 32447 32895
rect 32597 32861 32631 32895
rect 33793 32861 33827 32895
rect 33977 32861 34011 32895
rect 36010 32861 36044 32895
rect 36277 32861 36311 32895
rect 7941 32793 7975 32827
rect 8309 32793 8343 32827
rect 14372 32793 14406 32827
rect 16589 32793 16623 32827
rect 18613 32793 18647 32827
rect 19349 32793 19383 32827
rect 23673 32793 23707 32827
rect 28733 32793 28767 32827
rect 29929 32793 29963 32827
rect 30757 32793 30791 32827
rect 3893 32725 3927 32759
rect 6377 32725 6411 32759
rect 15485 32725 15519 32759
rect 16865 32725 16899 32759
rect 17969 32725 18003 32759
rect 27445 32725 27479 32759
rect 30665 32725 30699 32759
rect 31401 32725 31435 32759
rect 8309 32521 8343 32555
rect 14473 32521 14507 32555
rect 18429 32521 18463 32555
rect 20729 32521 20763 32555
rect 24133 32521 24167 32555
rect 29929 32521 29963 32555
rect 36277 32521 36311 32555
rect 10241 32453 10275 32487
rect 12541 32453 12575 32487
rect 15117 32453 15151 32487
rect 16129 32453 16163 32487
rect 19594 32453 19628 32487
rect 25246 32453 25280 32487
rect 28641 32453 28675 32487
rect 32505 32453 32539 32487
rect 2237 32385 2271 32419
rect 2493 32385 2527 32419
rect 6377 32385 6411 32419
rect 6633 32385 6667 32419
rect 9505 32385 9539 32419
rect 10425 32385 10459 32419
rect 12725 32385 12759 32419
rect 13829 32385 13863 32419
rect 14013 32385 14047 32419
rect 14105 32385 14139 32419
rect 14197 32385 14231 32419
rect 14933 32385 14967 32419
rect 15945 32385 15979 32419
rect 17141 32385 17175 32419
rect 19349 32385 19383 32419
rect 22661 32385 22695 32419
rect 23489 32385 23523 32419
rect 25513 32385 25547 32419
rect 28549 32385 28583 32419
rect 28733 32385 28767 32419
rect 28917 32385 28951 32419
rect 29745 32385 29779 32419
rect 30481 32385 30515 32419
rect 32137 32385 32171 32419
rect 32321 32385 32355 32419
rect 34989 32385 35023 32419
rect 9781 32317 9815 32351
rect 15301 32317 15335 32351
rect 21281 32317 21315 32351
rect 22385 32317 22419 32351
rect 23673 32249 23707 32283
rect 34529 32249 34563 32283
rect 3617 32181 3651 32215
rect 7757 32181 7791 32215
rect 10609 32181 10643 32215
rect 12909 32181 12943 32215
rect 28365 32181 28399 32215
rect 58173 32181 58207 32215
rect 2053 31977 2087 32011
rect 7021 31977 7055 32011
rect 17049 31977 17083 32011
rect 28917 31977 28951 32011
rect 29745 31977 29779 32011
rect 35541 31977 35575 32011
rect 10701 31909 10735 31943
rect 14197 31909 14231 31943
rect 21557 31909 21591 31943
rect 9321 31841 9355 31875
rect 11437 31841 11471 31875
rect 17785 31841 17819 31875
rect 23581 31841 23615 31875
rect 24961 31841 24995 31875
rect 36737 31841 36771 31875
rect 37565 31841 37599 31875
rect 2283 31773 2317 31807
rect 2402 31773 2436 31807
rect 2534 31773 2568 31807
rect 2697 31773 2731 31807
rect 5733 31773 5767 31807
rect 8309 31773 8343 31807
rect 9588 31773 9622 31807
rect 11704 31773 11738 31807
rect 17509 31773 17543 31807
rect 22109 31773 22143 31807
rect 23857 31773 23891 31807
rect 25237 31773 25271 31807
rect 30858 31773 30892 31807
rect 31125 31773 31159 31807
rect 36099 31773 36133 31807
rect 36277 31773 36311 31807
rect 36369 31773 36403 31807
rect 36507 31773 36541 31807
rect 37821 31773 37855 31807
rect 7941 31705 7975 31739
rect 8125 31705 8159 31739
rect 22291 31705 22325 31739
rect 3249 31637 3283 31671
rect 12817 31637 12851 31671
rect 22477 31637 22511 31671
rect 38945 31637 38979 31671
rect 2421 31433 2455 31467
rect 5181 31433 5215 31467
rect 5641 31433 5675 31467
rect 9137 31433 9171 31467
rect 9689 31433 9723 31467
rect 10885 31433 10919 31467
rect 12909 31433 12943 31467
rect 30389 31433 30423 31467
rect 36185 31433 36219 31467
rect 2605 31365 2639 31399
rect 8401 31365 8435 31399
rect 8585 31365 8619 31399
rect 23397 31365 23431 31399
rect 31125 31365 31159 31399
rect 36001 31365 36035 31399
rect 2789 31297 2823 31331
rect 5825 31297 5859 31331
rect 6653 31297 6687 31331
rect 7113 31297 7147 31331
rect 7297 31297 7331 31331
rect 7389 31297 7423 31331
rect 7481 31297 7515 31331
rect 9965 31297 9999 31331
rect 10057 31297 10091 31331
rect 10149 31297 10183 31331
rect 10333 31297 10367 31331
rect 11713 31297 11747 31331
rect 11897 31297 11931 31331
rect 13185 31297 13219 31331
rect 13274 31297 13308 31331
rect 13369 31297 13403 31331
rect 13553 31297 13587 31331
rect 15117 31297 15151 31331
rect 15209 31297 15243 31331
rect 15301 31297 15335 31331
rect 15485 31297 15519 31331
rect 19789 31297 19823 31331
rect 22293 31297 22327 31331
rect 22385 31297 22419 31331
rect 22482 31297 22516 31331
rect 22661 31297 22695 31331
rect 23213 31297 23247 31331
rect 30205 31297 30239 31331
rect 31033 31297 31067 31331
rect 31217 31297 31251 31331
rect 31401 31297 31435 31331
rect 32321 31297 32355 31331
rect 35817 31297 35851 31331
rect 19533 31229 19567 31263
rect 30021 31229 30055 31263
rect 32137 31161 32171 31195
rect 7757 31093 7791 31127
rect 11529 31093 11563 31127
rect 12449 31093 12483 31127
rect 14013 31093 14047 31127
rect 14841 31093 14875 31127
rect 16037 31093 16071 31127
rect 18981 31093 19015 31127
rect 20913 31093 20947 31127
rect 22017 31093 22051 31127
rect 23949 31093 23983 31127
rect 25053 31093 25087 31127
rect 29469 31093 29503 31127
rect 30849 31093 30883 31127
rect 5917 30889 5951 30923
rect 6377 30889 6411 30923
rect 8033 30889 8067 30923
rect 11897 30889 11931 30923
rect 29653 30889 29687 30923
rect 39313 30889 39347 30923
rect 9045 30821 9079 30855
rect 14197 30821 14231 30855
rect 24409 30821 24443 30855
rect 14841 30753 14875 30787
rect 25605 30753 25639 30787
rect 27537 30753 27571 30787
rect 32321 30753 32355 30787
rect 37013 30753 37047 30787
rect 37933 30753 37967 30787
rect 2605 30685 2639 30719
rect 5549 30685 5583 30719
rect 6653 30685 6687 30719
rect 6745 30685 6779 30719
rect 6837 30685 6871 30719
rect 7021 30685 7055 30719
rect 8125 30685 8159 30719
rect 12633 30685 12667 30719
rect 12909 30685 12943 30719
rect 13025 30685 13059 30719
rect 15097 30685 15131 30719
rect 16865 30685 16899 30719
rect 17049 30685 17083 30719
rect 19717 30685 19751 30719
rect 20269 30685 20303 30719
rect 20545 30685 20579 30719
rect 21741 30685 21775 30719
rect 22008 30685 22042 30719
rect 24961 30685 24995 30719
rect 25145 30685 25179 30719
rect 25256 30685 25290 30719
rect 25375 30685 25409 30719
rect 27270 30685 27304 30719
rect 30389 30685 30423 30719
rect 30757 30685 30791 30719
rect 31217 30685 31251 30719
rect 31401 30685 31435 30719
rect 31493 30685 31527 30719
rect 31585 30685 31619 30719
rect 35265 30685 35299 30719
rect 35909 30685 35943 30719
rect 36093 30682 36127 30716
rect 36188 30682 36222 30716
rect 36277 30685 36311 30719
rect 58173 30685 58207 30719
rect 2789 30617 2823 30651
rect 5733 30617 5767 30651
rect 10425 30617 10459 30651
rect 12817 30617 12851 30651
rect 16681 30617 16715 30651
rect 18337 30617 18371 30651
rect 18521 30617 18555 30651
rect 30481 30617 30515 30651
rect 30573 30617 30607 30651
rect 31861 30617 31895 30651
rect 32566 30617 32600 30651
rect 35081 30617 35115 30651
rect 35449 30617 35483 30651
rect 36553 30617 36587 30651
rect 38178 30617 38212 30651
rect 2421 30549 2455 30583
rect 13185 30549 13219 30583
rect 16221 30549 16255 30583
rect 17785 30549 17819 30583
rect 18705 30549 18739 30583
rect 23121 30549 23155 30583
rect 23673 30549 23707 30583
rect 26157 30549 26191 30583
rect 30205 30549 30239 30583
rect 33701 30549 33735 30583
rect 11805 30345 11839 30379
rect 17233 30345 17267 30379
rect 19073 30345 19107 30379
rect 19533 30345 19567 30379
rect 35357 30345 35391 30379
rect 37657 30345 37691 30379
rect 4629 30277 4663 30311
rect 15393 30277 15427 30311
rect 15485 30277 15519 30311
rect 21005 30277 21039 30311
rect 22477 30277 22511 30311
rect 24593 30277 24627 30311
rect 32229 30277 32263 30311
rect 32597 30277 32631 30311
rect 33609 30277 33643 30311
rect 33701 30277 33735 30311
rect 34621 30277 34655 30311
rect 37289 30277 37323 30311
rect 2421 30209 2455 30243
rect 2677 30209 2711 30243
rect 4445 30209 4479 30243
rect 7501 30209 7535 30243
rect 7757 30209 7791 30243
rect 11989 30209 12023 30243
rect 15117 30209 15151 30243
rect 15265 30209 15299 30243
rect 15582 30209 15616 30243
rect 17693 30209 17727 30243
rect 17960 30209 17994 30243
rect 19809 30209 19843 30243
rect 19914 30212 19948 30246
rect 20014 30212 20048 30246
rect 20189 30209 20223 30243
rect 20637 30209 20671 30243
rect 20821 30209 20855 30243
rect 22385 30209 22419 30243
rect 22569 30209 22603 30243
rect 22753 30209 22787 30243
rect 24225 30209 24259 30243
rect 24409 30209 24443 30243
rect 25414 30209 25448 30243
rect 26157 30209 26191 30243
rect 28733 30209 28767 30243
rect 28825 30209 28859 30243
rect 28917 30209 28951 30243
rect 29101 30209 29135 30243
rect 30481 30209 30515 30243
rect 32413 30209 32447 30243
rect 33517 30209 33551 30243
rect 33885 30209 33919 30243
rect 34529 30209 34563 30243
rect 34713 30209 34747 30243
rect 34897 30209 34931 30243
rect 35909 30209 35943 30243
rect 36072 30215 36106 30249
rect 36185 30209 36219 30243
rect 36323 30209 36357 30243
rect 37473 30209 37507 30243
rect 12173 30141 12207 30175
rect 30205 30141 30239 30175
rect 3801 30073 3835 30107
rect 25237 30073 25271 30107
rect 25973 30073 26007 30107
rect 31493 30073 31527 30107
rect 4261 30005 4295 30039
rect 6377 30005 6411 30039
rect 10517 30005 10551 30039
rect 12725 30005 12759 30039
rect 15761 30005 15795 30039
rect 22201 30005 22235 30039
rect 26985 30005 27019 30039
rect 27905 30005 27939 30039
rect 28457 30005 28491 30039
rect 33333 30005 33367 30039
rect 34345 30005 34379 30039
rect 36553 30005 36587 30039
rect 2145 29801 2179 29835
rect 9137 29801 9171 29835
rect 11989 29801 12023 29835
rect 15485 29801 15519 29835
rect 18061 29801 18095 29835
rect 19441 29801 19475 29835
rect 20729 29801 20763 29835
rect 21557 29801 21591 29835
rect 23857 29801 23891 29835
rect 29009 29801 29043 29835
rect 30665 29801 30699 29835
rect 34897 29801 34931 29835
rect 16957 29733 16991 29767
rect 20177 29733 20211 29767
rect 37933 29733 37967 29767
rect 9505 29665 9539 29699
rect 9965 29665 9999 29699
rect 27169 29665 27203 29699
rect 35357 29665 35391 29699
rect 35633 29665 35667 29699
rect 2375 29597 2409 29631
rect 2494 29594 2528 29628
rect 2605 29597 2639 29631
rect 2789 29597 2823 29631
rect 4169 29597 4203 29631
rect 4445 29597 4479 29631
rect 4537 29597 4571 29631
rect 9321 29597 9355 29631
rect 10609 29597 10643 29631
rect 15117 29597 15151 29631
rect 15301 29597 15335 29631
rect 18337 29597 18371 29631
rect 18429 29597 18463 29631
rect 18521 29597 18555 29631
rect 18705 29597 18739 29631
rect 20821 29597 20855 29631
rect 21373 29597 21407 29631
rect 22201 29597 22235 29631
rect 22569 29597 22603 29631
rect 24685 29597 24719 29631
rect 24869 29597 24903 29631
rect 24961 29597 24995 29631
rect 25053 29597 25087 29631
rect 28641 29597 28675 29631
rect 28825 29597 28859 29631
rect 29745 29597 29779 29631
rect 29837 29597 29871 29631
rect 30113 29597 30147 29631
rect 30573 29597 30607 29631
rect 30757 29597 30791 29631
rect 31217 29597 31251 29631
rect 33793 29597 33827 29631
rect 33977 29597 34011 29631
rect 34161 29597 34195 29631
rect 34713 29597 34747 29631
rect 39313 29597 39347 29631
rect 58173 29597 58207 29631
rect 4353 29529 4387 29563
rect 10876 29529 10910 29563
rect 17509 29529 17543 29563
rect 19993 29529 20027 29563
rect 22385 29529 22419 29563
rect 22477 29529 22511 29563
rect 25329 29529 25363 29563
rect 26902 29529 26936 29563
rect 29929 29529 29963 29563
rect 33885 29529 33919 29563
rect 39046 29529 39080 29563
rect 4721 29461 4755 29495
rect 7205 29461 7239 29495
rect 14197 29461 14231 29495
rect 22753 29461 22787 29495
rect 25789 29461 25823 29495
rect 29561 29461 29595 29495
rect 33609 29461 33643 29495
rect 36645 29461 36679 29495
rect 10977 29257 11011 29291
rect 18797 29257 18831 29291
rect 20453 29257 20487 29291
rect 21281 29257 21315 29291
rect 24409 29257 24443 29291
rect 24961 29257 24995 29291
rect 29929 29257 29963 29291
rect 31217 29257 31251 29291
rect 36737 29257 36771 29291
rect 38577 29257 38611 29291
rect 4445 29189 4479 29223
rect 5549 29189 5583 29223
rect 14933 29189 14967 29223
rect 24225 29189 24259 29223
rect 35449 29189 35483 29223
rect 35633 29189 35667 29223
rect 39690 29189 39724 29223
rect 3019 29121 3053 29155
rect 3157 29121 3191 29155
rect 3270 29127 3304 29161
rect 3433 29121 3467 29155
rect 4261 29121 4295 29155
rect 4537 29121 4571 29155
rect 4629 29121 4663 29155
rect 5273 29121 5307 29155
rect 5457 29121 5491 29155
rect 5641 29121 5675 29155
rect 7849 29121 7883 29155
rect 8116 29121 8150 29155
rect 10339 29121 10373 29155
rect 10512 29124 10546 29158
rect 10609 29121 10643 29155
rect 10701 29121 10735 29155
rect 13461 29121 13495 29155
rect 13553 29121 13587 29155
rect 13645 29121 13679 29155
rect 13829 29121 13863 29155
rect 15117 29121 15151 29155
rect 19257 29121 19291 29155
rect 19441 29121 19475 29155
rect 19533 29121 19567 29155
rect 19625 29121 19659 29155
rect 22569 29121 22603 29155
rect 24041 29121 24075 29155
rect 25145 29121 25179 29155
rect 25881 29121 25915 29155
rect 28641 29121 28675 29155
rect 31033 29121 31067 29155
rect 33517 29121 33551 29155
rect 35265 29121 35299 29155
rect 36093 29121 36127 29155
rect 36277 29121 36311 29155
rect 36369 29121 36403 29155
rect 36507 29121 36541 29155
rect 30849 29053 30883 29087
rect 33793 29053 33827 29087
rect 39957 29053 39991 29087
rect 4813 28985 4847 29019
rect 13185 28985 13219 29019
rect 14381 28985 14415 29019
rect 18245 28985 18279 29019
rect 19809 28985 19843 29019
rect 22753 28985 22787 29019
rect 25697 28985 25731 29019
rect 28089 28985 28123 29019
rect 2789 28917 2823 28951
rect 5825 28917 5859 28951
rect 9229 28917 9263 28951
rect 9873 28917 9907 28951
rect 15301 28917 15335 28951
rect 16037 28917 16071 28951
rect 26433 28917 26467 28951
rect 2881 28713 2915 28747
rect 9045 28713 9079 28747
rect 13553 28713 13587 28747
rect 14473 28713 14507 28747
rect 19717 28713 19751 28747
rect 20453 28713 20487 28747
rect 24777 28713 24811 28747
rect 26985 28713 27019 28747
rect 29009 28713 29043 28747
rect 31401 28713 31435 28747
rect 8401 28577 8435 28611
rect 30389 28577 30423 28611
rect 33517 28577 33551 28611
rect 8125 28509 8159 28543
rect 8309 28509 8343 28543
rect 9275 28509 9309 28543
rect 9413 28509 9447 28543
rect 9505 28509 9539 28543
rect 9689 28509 9723 28543
rect 12449 28509 12483 28543
rect 12633 28509 12667 28543
rect 12817 28509 12851 28543
rect 14289 28509 14323 28543
rect 14933 28509 14967 28543
rect 15117 28509 15151 28543
rect 15209 28509 15243 28543
rect 15301 28509 15335 28543
rect 21465 28509 21499 28543
rect 21649 28509 21683 28543
rect 21833 28509 21867 28543
rect 24961 28509 24995 28543
rect 26433 28509 26467 28543
rect 27169 28509 27203 28543
rect 27629 28509 27663 28543
rect 27896 28509 27930 28543
rect 30113 28509 30147 28543
rect 33793 28509 33827 28543
rect 34897 28509 34931 28543
rect 34989 28509 35023 28543
rect 35265 28509 35299 28543
rect 36185 28509 36219 28543
rect 36369 28509 36403 28543
rect 36461 28509 36495 28543
rect 36553 28509 36587 28543
rect 38761 28509 38795 28543
rect 7573 28441 7607 28475
rect 12725 28441 12759 28475
rect 14105 28441 14139 28475
rect 16221 28441 16255 28475
rect 16405 28441 16439 28475
rect 21557 28441 21591 28475
rect 23857 28441 23891 28475
rect 35081 28441 35115 28475
rect 36829 28441 36863 28475
rect 38494 28441 38528 28475
rect 3893 28373 3927 28407
rect 10241 28373 10275 28407
rect 10793 28373 10827 28407
rect 13001 28373 13035 28407
rect 15577 28373 15611 28407
rect 21281 28373 21315 28407
rect 25513 28373 25547 28407
rect 29561 28373 29595 28407
rect 34713 28373 34747 28407
rect 37381 28373 37415 28407
rect 3893 28169 3927 28203
rect 8493 28169 8527 28203
rect 9321 28169 9355 28203
rect 11529 28169 11563 28203
rect 14749 28169 14783 28203
rect 23581 28169 23615 28203
rect 24317 28169 24351 28203
rect 36369 28169 36403 28203
rect 2780 28101 2814 28135
rect 7021 28101 7055 28135
rect 7849 28101 7883 28135
rect 8953 28101 8987 28135
rect 9137 28101 9171 28135
rect 13921 28101 13955 28135
rect 22293 28101 22327 28135
rect 34253 28101 34287 28135
rect 36185 28101 36219 28135
rect 6653 28033 6687 28067
rect 6746 28033 6780 28067
rect 6929 28033 6963 28067
rect 7159 28033 7193 28067
rect 8309 28033 8343 28067
rect 8493 28033 8527 28067
rect 11713 28033 11747 28067
rect 13553 28033 13587 28067
rect 13646 28033 13680 28067
rect 13829 28033 13863 28067
rect 14018 28033 14052 28067
rect 15862 28033 15896 28067
rect 16129 28033 16163 28067
rect 18337 28033 18371 28067
rect 19717 28033 19751 28067
rect 24133 28033 24167 28067
rect 30021 28033 30055 28067
rect 30205 28033 30239 28067
rect 31309 28033 31343 28067
rect 34161 28033 34195 28067
rect 34345 28033 34379 28067
rect 34529 28033 34563 28067
rect 36001 28033 36035 28067
rect 2513 27965 2547 27999
rect 10701 27965 10735 27999
rect 10977 27965 11011 27999
rect 11897 27965 11931 27999
rect 18061 27965 18095 27999
rect 19441 27965 19475 27999
rect 31585 27965 31619 27999
rect 32137 27965 32171 27999
rect 7297 27897 7331 27931
rect 12449 27897 12483 27931
rect 22477 27897 22511 27931
rect 58173 27897 58207 27931
rect 14197 27829 14231 27863
rect 16865 27829 16899 27863
rect 24961 27829 24995 27863
rect 29469 27829 29503 27863
rect 30113 27829 30147 27863
rect 33977 27829 34011 27863
rect 11529 27625 11563 27659
rect 13553 27625 13587 27659
rect 36001 27625 36035 27659
rect 5641 27557 5675 27591
rect 10977 27557 11011 27591
rect 15577 27557 15611 27591
rect 18061 27557 18095 27591
rect 20269 27557 20303 27591
rect 9045 27489 9079 27523
rect 9873 27489 9907 27523
rect 12173 27489 12207 27523
rect 30389 27489 30423 27523
rect 4997 27421 5031 27455
rect 5090 27421 5124 27455
rect 5365 27421 5399 27455
rect 5503 27421 5537 27455
rect 7573 27421 7607 27455
rect 9505 27421 9539 27455
rect 9781 27421 9815 27455
rect 12440 27421 12474 27455
rect 16497 27421 16531 27455
rect 16681 27421 16715 27455
rect 17417 27421 17451 27455
rect 17877 27421 17911 27455
rect 20821 27421 20855 27455
rect 25053 27421 25087 27455
rect 25237 27421 25271 27455
rect 25329 27421 25363 27455
rect 25421 27421 25455 27455
rect 26525 27421 26559 27455
rect 30665 27421 30699 27455
rect 31125 27421 31159 27455
rect 31401 27421 31435 27455
rect 32597 27421 32631 27455
rect 32689 27421 32723 27455
rect 32965 27421 32999 27455
rect 33793 27421 33827 27455
rect 5273 27353 5307 27387
rect 7389 27353 7423 27387
rect 10793 27353 10827 27387
rect 11621 27353 11655 27387
rect 14841 27353 14875 27387
rect 15393 27353 15427 27387
rect 16589 27353 16623 27387
rect 22569 27353 22603 27387
rect 25697 27353 25731 27387
rect 26770 27353 26804 27387
rect 29009 27353 29043 27387
rect 32781 27353 32815 27387
rect 33609 27353 33643 27387
rect 3157 27285 3191 27319
rect 3893 27285 3927 27319
rect 7757 27285 7791 27319
rect 24501 27285 24535 27319
rect 27905 27285 27939 27319
rect 32413 27285 32447 27319
rect 33425 27285 33459 27319
rect 6377 27081 6411 27115
rect 9505 27081 9539 27115
rect 30941 27081 30975 27115
rect 5273 27013 5307 27047
rect 7512 27013 7546 27047
rect 8217 27013 8251 27047
rect 9597 27013 9631 27047
rect 29745 27013 29779 27047
rect 35357 27013 35391 27047
rect 2881 26945 2915 26979
rect 2970 26951 3004 26985
rect 3070 26945 3104 26979
rect 3249 26945 3283 26979
rect 3893 26945 3927 26979
rect 4077 26945 4111 26979
rect 4905 26945 4939 26979
rect 4998 26945 5032 26979
rect 5181 26945 5215 26979
rect 5411 26945 5445 26979
rect 8493 26945 8527 26979
rect 8585 26945 8619 26979
rect 8677 26945 8711 26979
rect 8861 26945 8895 26979
rect 10149 26945 10183 26979
rect 11897 26945 11931 26979
rect 13185 26945 13219 26979
rect 17141 26945 17175 26979
rect 17408 26945 17442 26979
rect 18981 26945 19015 26979
rect 19248 26945 19282 26979
rect 21005 26945 21039 26979
rect 21833 26945 21867 26979
rect 22017 26945 22051 26979
rect 23774 26945 23808 26979
rect 24041 26945 24075 26979
rect 25053 26945 25087 26979
rect 25320 26945 25354 26979
rect 28161 26945 28195 26979
rect 29929 26945 29963 26979
rect 32413 26945 32447 26979
rect 32597 26945 32631 26979
rect 32689 26945 32723 26979
rect 32781 26945 32815 26979
rect 33885 26945 33919 26979
rect 34069 26945 34103 26979
rect 34161 26945 34195 26979
rect 34299 26945 34333 26979
rect 34989 26945 35023 26979
rect 35173 26945 35207 26979
rect 38669 26945 38703 26979
rect 39129 26945 39163 26979
rect 3709 26877 3743 26911
rect 7757 26877 7791 26911
rect 10425 26877 10459 26911
rect 11621 26877 11655 26911
rect 12909 26877 12943 26911
rect 27905 26877 27939 26911
rect 20361 26809 20395 26843
rect 2605 26741 2639 26775
rect 5549 26741 5583 26775
rect 18521 26741 18555 26775
rect 21189 26741 21223 26775
rect 22201 26741 22235 26775
rect 22661 26741 22695 26775
rect 26433 26741 26467 26775
rect 29285 26741 29319 26775
rect 33057 26741 33091 26775
rect 34529 26741 34563 26775
rect 40417 26741 40451 26775
rect 58173 26741 58207 26775
rect 9505 26537 9539 26571
rect 11437 26537 11471 26571
rect 17233 26537 17267 26571
rect 18705 26537 18739 26571
rect 22477 26537 22511 26571
rect 25329 26537 25363 26571
rect 26433 26537 26467 26571
rect 29653 26537 29687 26571
rect 30113 26537 30147 26571
rect 7481 26469 7515 26503
rect 32229 26469 32263 26503
rect 34713 26469 34747 26503
rect 37933 26469 37967 26503
rect 10793 26401 10827 26435
rect 12633 26401 12667 26435
rect 21281 26401 21315 26435
rect 33885 26401 33919 26435
rect 2145 26333 2179 26367
rect 2881 26333 2915 26367
rect 2973 26330 3007 26364
rect 3065 26333 3099 26367
rect 3249 26333 3283 26367
rect 3985 26333 4019 26367
rect 4169 26333 4203 26367
rect 6009 26333 6043 26367
rect 6844 26333 6878 26367
rect 6985 26333 7019 26367
rect 7113 26333 7147 26367
rect 7343 26333 7377 26367
rect 8033 26333 8067 26367
rect 9413 26333 9447 26367
rect 9597 26333 9631 26367
rect 10609 26333 10643 26367
rect 12909 26333 12943 26367
rect 16405 26333 16439 26367
rect 16865 26333 16899 26367
rect 17049 26333 17083 26367
rect 18061 26333 18095 26367
rect 18245 26333 18279 26367
rect 18337 26333 18371 26367
rect 18429 26333 18463 26367
rect 19349 26333 19383 26367
rect 21833 26333 21867 26367
rect 21996 26333 22030 26367
rect 22109 26333 22143 26367
rect 22247 26333 22281 26367
rect 24685 26333 24719 26367
rect 24869 26333 24903 26367
rect 24964 26333 24998 26367
rect 25099 26333 25133 26367
rect 25789 26333 25823 26367
rect 25952 26333 25986 26367
rect 26065 26333 26099 26367
rect 26203 26333 26237 26367
rect 27261 26333 27295 26367
rect 32965 26333 32999 26367
rect 33057 26333 33091 26367
rect 33149 26333 33183 26367
rect 33333 26333 33367 26367
rect 35826 26333 35860 26367
rect 36093 26333 36127 26367
rect 39313 26333 39347 26367
rect 40049 26333 40083 26367
rect 2605 26265 2639 26299
rect 3801 26265 3835 26299
rect 4721 26265 4755 26299
rect 6193 26265 6227 26299
rect 7205 26265 7239 26299
rect 11345 26265 11379 26299
rect 13461 26265 13495 26299
rect 20821 26265 20855 26299
rect 26893 26265 26927 26299
rect 27077 26265 27111 26299
rect 39068 26265 39102 26299
rect 39865 26265 39899 26299
rect 6377 26197 6411 26231
rect 32781 26197 32815 26231
rect 40233 26197 40267 26231
rect 40785 26197 40819 26231
rect 3985 25993 4019 26027
rect 7573 25993 7607 26027
rect 9045 25993 9079 26027
rect 10609 25993 10643 26027
rect 13553 25993 13587 26027
rect 17693 25993 17727 26027
rect 18797 25993 18831 26027
rect 25789 25993 25823 26027
rect 26985 25993 27019 26027
rect 34345 25993 34379 26027
rect 2872 25925 2906 25959
rect 8033 25925 8067 25959
rect 10701 25925 10735 25959
rect 18981 25925 19015 25959
rect 21281 25925 21315 25959
rect 25329 25925 25363 25959
rect 26157 25925 26191 25959
rect 27721 25925 27755 25959
rect 33232 25925 33266 25959
rect 39712 25925 39746 25959
rect 41061 25925 41095 25959
rect 6377 25857 6411 25891
rect 6561 25857 6595 25891
rect 6653 25857 6687 25891
rect 6745 25857 6779 25891
rect 13645 25857 13679 25891
rect 14289 25857 14323 25891
rect 15761 25857 15795 25891
rect 16865 25857 16899 25891
rect 17923 25857 17957 25891
rect 18061 25857 18095 25891
rect 18174 25857 18208 25891
rect 18337 25857 18371 25891
rect 19165 25857 19199 25891
rect 19809 25857 19843 25891
rect 19993 25857 20027 25891
rect 20913 25857 20947 25891
rect 21097 25857 21131 25891
rect 21833 25857 21867 25891
rect 21996 25857 22030 25891
rect 22109 25857 22143 25891
rect 22247 25857 22281 25891
rect 23029 25857 23063 25891
rect 25973 25857 26007 25891
rect 29929 25857 29963 25891
rect 30113 25857 30147 25891
rect 40417 25857 40451 25891
rect 40601 25857 40635 25891
rect 40693 25857 40727 25891
rect 40785 25857 40819 25891
rect 2605 25789 2639 25823
rect 9781 25789 9815 25823
rect 15485 25789 15519 25823
rect 19625 25789 19659 25823
rect 32965 25789 32999 25823
rect 39957 25789 39991 25823
rect 14473 25721 14507 25755
rect 38577 25721 38611 25755
rect 7021 25653 7055 25687
rect 12909 25653 12943 25687
rect 16681 25653 16715 25687
rect 22477 25653 22511 25687
rect 29009 25653 29043 25687
rect 30297 25653 30331 25687
rect 37381 25653 37415 25687
rect 7757 25449 7791 25483
rect 8401 25449 8435 25483
rect 25605 25449 25639 25483
rect 31309 25449 31343 25483
rect 39313 25449 39347 25483
rect 39865 25449 39899 25483
rect 12081 25313 12115 25347
rect 37105 25313 37139 25347
rect 4353 25245 4387 25279
rect 6377 25245 6411 25279
rect 6644 25245 6678 25279
rect 9505 25245 9539 25279
rect 9597 25245 9631 25279
rect 9689 25245 9723 25279
rect 9873 25245 9907 25279
rect 12541 25245 12575 25279
rect 13553 25245 13587 25279
rect 18061 25245 18095 25279
rect 18245 25245 18279 25279
rect 18337 25245 18371 25279
rect 18475 25245 18509 25279
rect 23029 25245 23063 25279
rect 25973 25245 26007 25279
rect 29837 25245 29871 25279
rect 29926 25242 29960 25276
rect 30021 25239 30055 25273
rect 30205 25245 30239 25279
rect 32689 25245 32723 25279
rect 37795 25245 37829 25279
rect 37946 25245 37980 25279
rect 38046 25245 38080 25279
rect 38209 25245 38243 25279
rect 38945 25245 38979 25279
rect 40141 25245 40175 25279
rect 40230 25245 40264 25279
rect 40325 25245 40359 25279
rect 40521 25245 40555 25279
rect 58173 25245 58207 25279
rect 5917 25177 5951 25211
rect 10333 25177 10367 25211
rect 15117 25177 15151 25211
rect 15301 25177 15335 25211
rect 16221 25177 16255 25211
rect 16773 25177 16807 25211
rect 16957 25177 16991 25211
rect 22762 25177 22796 25211
rect 25789 25177 25823 25211
rect 32422 25177 32456 25211
rect 36860 25177 36894 25211
rect 37565 25177 37599 25211
rect 39129 25177 39163 25211
rect 9229 25109 9263 25143
rect 14105 25109 14139 25143
rect 14933 25109 14967 25143
rect 17601 25109 17635 25143
rect 18705 25109 18739 25143
rect 19349 25109 19383 25143
rect 21649 25109 21683 25143
rect 28917 25109 28951 25143
rect 29561 25109 29595 25143
rect 30757 25109 30791 25143
rect 35725 25109 35759 25143
rect 40969 25109 41003 25143
rect 3893 24905 3927 24939
rect 6469 24905 6503 24939
rect 8861 24905 8895 24939
rect 22661 24837 22695 24871
rect 2780 24769 2814 24803
rect 9045 24769 9079 24803
rect 9229 24769 9263 24803
rect 9919 24769 9953 24803
rect 10057 24769 10091 24803
rect 10149 24769 10183 24803
rect 10333 24769 10367 24803
rect 13553 24769 13587 24803
rect 13737 24769 13771 24803
rect 14729 24769 14763 24803
rect 16957 24769 16991 24803
rect 18889 24769 18923 24803
rect 19156 24769 19190 24803
rect 22523 24769 22557 24803
rect 22753 24769 22787 24803
rect 22881 24769 22915 24803
rect 23029 24769 23063 24803
rect 24869 24769 24903 24803
rect 25053 24769 25087 24803
rect 25145 24769 25179 24803
rect 25237 24769 25271 24803
rect 29949 24769 29983 24803
rect 30665 24769 30699 24803
rect 30849 24772 30883 24806
rect 30941 24769 30975 24803
rect 31033 24769 31067 24803
rect 32137 24769 32171 24803
rect 33517 24769 33551 24803
rect 33977 24769 34011 24803
rect 37289 24769 37323 24803
rect 37473 24769 37507 24803
rect 39782 24769 39816 24803
rect 40049 24769 40083 24803
rect 2513 24701 2547 24735
rect 12541 24701 12575 24735
rect 14473 24701 14507 24735
rect 18153 24701 18187 24735
rect 18429 24701 18463 24735
rect 30205 24701 30239 24735
rect 31309 24701 31343 24735
rect 35725 24701 35759 24735
rect 37657 24701 37691 24735
rect 24409 24633 24443 24667
rect 9689 24565 9723 24599
rect 10793 24565 10827 24599
rect 12081 24565 12115 24599
rect 13369 24565 13403 24599
rect 15853 24565 15887 24599
rect 16773 24565 16807 24599
rect 20269 24565 20303 24599
rect 22385 24565 22419 24599
rect 25513 24565 25547 24599
rect 28273 24565 28307 24599
rect 28825 24565 28859 24599
rect 38669 24565 38703 24599
rect 14381 24361 14415 24395
rect 15485 24361 15519 24395
rect 19257 24361 19291 24395
rect 24593 24361 24627 24395
rect 28181 24361 28215 24395
rect 30205 24361 30239 24395
rect 30665 24293 30699 24327
rect 10333 24225 10367 24259
rect 18153 24225 18187 24259
rect 10066 24157 10100 24191
rect 11897 24157 11931 24191
rect 11989 24157 12023 24191
rect 12081 24157 12115 24191
rect 12265 24157 12299 24191
rect 13001 24157 13035 24191
rect 13093 24157 13127 24191
rect 13185 24157 13219 24191
rect 13369 24157 13403 24191
rect 14657 24157 14691 24191
rect 14746 24154 14780 24188
rect 14846 24157 14880 24191
rect 15025 24157 15059 24191
rect 18429 24157 18463 24191
rect 19441 24157 19475 24191
rect 20961 24157 20995 24191
rect 21097 24157 21131 24191
rect 21372 24157 21406 24191
rect 21465 24157 21499 24191
rect 22063 24157 22097 24191
rect 22293 24157 22327 24191
rect 22476 24157 22510 24191
rect 22569 24157 22603 24191
rect 24777 24157 24811 24191
rect 24961 24157 24995 24191
rect 25421 24157 25455 24191
rect 28825 24157 28859 24191
rect 29561 24157 29595 24191
rect 29724 24157 29758 24191
rect 29824 24154 29858 24188
rect 29929 24157 29963 24191
rect 40233 24157 40267 24191
rect 41061 24157 41095 24191
rect 58173 24157 58207 24191
rect 7849 24089 7883 24123
rect 19625 24089 19659 24123
rect 21189 24089 21223 24123
rect 22201 24089 22235 24123
rect 25666 24089 25700 24123
rect 27813 24089 27847 24123
rect 27997 24089 28031 24123
rect 28641 24089 28675 24123
rect 40049 24089 40083 24123
rect 40877 24089 40911 24123
rect 8953 24021 8987 24055
rect 11161 24021 11195 24055
rect 11621 24021 11655 24055
rect 12725 24021 12759 24055
rect 16589 24021 16623 24055
rect 20821 24021 20855 24055
rect 21925 24021 21959 24055
rect 26801 24021 26835 24055
rect 29009 24021 29043 24055
rect 40417 24021 40451 24055
rect 41245 24021 41279 24055
rect 10149 23817 10183 23851
rect 12173 23817 12207 23851
rect 14197 23817 14231 23851
rect 14657 23817 14691 23851
rect 18245 23817 18279 23851
rect 28549 23817 28583 23851
rect 32505 23817 32539 23851
rect 22753 23749 22787 23783
rect 24317 23749 24351 23783
rect 24961 23749 24995 23783
rect 33701 23749 33735 23783
rect 36093 23749 36127 23783
rect 2237 23681 2271 23715
rect 2421 23681 2455 23715
rect 7665 23681 7699 23715
rect 8309 23681 8343 23715
rect 8576 23681 8610 23715
rect 10333 23681 10367 23715
rect 10517 23681 10551 23715
rect 11805 23681 11839 23715
rect 11989 23681 12023 23715
rect 12817 23681 12851 23715
rect 13073 23681 13107 23715
rect 18061 23681 18095 23715
rect 22523 23681 22557 23715
rect 22661 23681 22695 23715
rect 22936 23681 22970 23715
rect 23029 23681 23063 23715
rect 25421 23681 25455 23715
rect 25605 23681 25639 23715
rect 25697 23681 25731 23715
rect 25789 23681 25823 23715
rect 29662 23681 29696 23715
rect 29929 23681 29963 23715
rect 33425 23681 33459 23715
rect 36001 23681 36035 23715
rect 36185 23681 36219 23715
rect 36369 23681 36403 23715
rect 39885 23681 39919 23715
rect 40141 23681 40175 23715
rect 40877 23681 40911 23715
rect 40969 23681 41003 23715
rect 41061 23681 41095 23715
rect 41245 23681 41279 23715
rect 7389 23613 7423 23647
rect 33517 23613 33551 23647
rect 40601 23613 40635 23647
rect 22385 23545 22419 23579
rect 33241 23545 33275 23579
rect 35817 23545 35851 23579
rect 2605 23477 2639 23511
rect 9689 23477 9723 23511
rect 26065 23477 26099 23511
rect 33701 23477 33735 23511
rect 38761 23477 38795 23511
rect 8125 23273 8159 23307
rect 12357 23273 12391 23307
rect 16865 23273 16899 23307
rect 21557 23273 21591 23307
rect 22385 23273 22419 23307
rect 29653 23273 29687 23307
rect 39957 23273 39991 23307
rect 41061 23273 41095 23307
rect 15945 23205 15979 23239
rect 39313 23205 39347 23239
rect 7573 23137 7607 23171
rect 14105 23137 14139 23171
rect 22477 23137 22511 23171
rect 25605 23137 25639 23171
rect 34069 23137 34103 23171
rect 35909 23137 35943 23171
rect 2559 23069 2593 23103
rect 2697 23069 2731 23103
rect 2789 23069 2823 23103
rect 2973 23069 3007 23103
rect 7297 23069 7331 23103
rect 10977 23069 11011 23103
rect 11244 23069 11278 23103
rect 12817 23069 12851 23103
rect 13001 23069 13035 23103
rect 13185 23069 13219 23103
rect 14841 23069 14875 23103
rect 15025 23069 15059 23103
rect 15209 23069 15243 23103
rect 22569 23069 22603 23103
rect 25872 23069 25906 23103
rect 40233 23069 40267 23103
rect 40325 23069 40359 23103
rect 40417 23069 40451 23103
rect 40601 23069 40635 23103
rect 15117 23001 15151 23035
rect 19257 23001 19291 23035
rect 19441 23001 19475 23035
rect 24869 23001 24903 23035
rect 31861 23001 31895 23035
rect 32045 23001 32079 23035
rect 33802 23001 33836 23035
rect 36176 23001 36210 23035
rect 2329 22933 2363 22967
rect 3801 22933 3835 22967
rect 15393 22933 15427 22967
rect 19625 22933 19659 22967
rect 22201 22933 22235 22967
rect 23765 22933 23799 22967
rect 24961 22933 24995 22967
rect 26985 22933 27019 22967
rect 32229 22933 32263 22967
rect 32689 22933 32723 22967
rect 35449 22933 35483 22967
rect 37289 22933 37323 22967
rect 1593 22729 1627 22763
rect 8493 22729 8527 22763
rect 9689 22729 9723 22763
rect 15577 22729 15611 22763
rect 16129 22729 16163 22763
rect 18061 22729 18095 22763
rect 25329 22729 25363 22763
rect 25973 22729 26007 22763
rect 33241 22729 33275 22763
rect 33701 22729 33735 22763
rect 36093 22729 36127 22763
rect 2666 22661 2700 22695
rect 4445 22661 4479 22695
rect 5457 22661 5491 22695
rect 5641 22661 5675 22695
rect 11805 22661 11839 22695
rect 14381 22661 14415 22695
rect 14473 22661 14507 22695
rect 26157 22661 26191 22695
rect 27905 22661 27939 22695
rect 31217 22661 31251 22695
rect 34069 22661 34103 22695
rect 35357 22661 35391 22695
rect 37473 22661 37507 22695
rect 39681 22661 39715 22695
rect 1777 22593 1811 22627
rect 1961 22593 1995 22627
rect 2421 22593 2455 22627
rect 4629 22593 4663 22627
rect 6653 22593 6687 22627
rect 6920 22593 6954 22627
rect 8677 22593 8711 22627
rect 9597 22593 9631 22627
rect 11529 22593 11563 22627
rect 11713 22593 11747 22627
rect 11897 22593 11931 22627
rect 14289 22593 14323 22627
rect 14657 22593 14691 22627
rect 18705 22593 18739 22627
rect 18961 22593 18995 22627
rect 20729 22593 20763 22627
rect 20913 22593 20947 22627
rect 22201 22593 22235 22627
rect 24133 22593 24167 22627
rect 25145 22593 25179 22627
rect 26341 22593 26375 22627
rect 28089 22593 28123 22627
rect 31033 22593 31067 22627
rect 31309 22593 31343 22627
rect 31401 22593 31435 22627
rect 32597 22593 32631 22627
rect 32760 22596 32794 22630
rect 32873 22593 32907 22627
rect 33011 22593 33045 22627
rect 33885 22593 33919 22627
rect 33977 22593 34011 22627
rect 34253 22593 34287 22627
rect 35265 22593 35299 22627
rect 35449 22593 35483 22627
rect 35633 22593 35667 22627
rect 36369 22593 36403 22627
rect 36461 22593 36495 22627
rect 36553 22593 36587 22627
rect 36737 22593 36771 22627
rect 37657 22593 37691 22627
rect 39497 22593 39531 22627
rect 16681 22525 16715 22559
rect 16957 22525 16991 22559
rect 22109 22525 22143 22559
rect 23857 22525 23891 22559
rect 37289 22525 37323 22559
rect 3801 22457 3835 22491
rect 8033 22457 8067 22491
rect 20085 22457 20119 22491
rect 58173 22457 58207 22491
rect 4261 22389 4295 22423
rect 5825 22389 5859 22423
rect 10333 22389 10367 22423
rect 12081 22389 12115 22423
rect 14105 22389 14139 22423
rect 20545 22389 20579 22423
rect 20913 22389 20947 22423
rect 21833 22389 21867 22423
rect 22017 22389 22051 22423
rect 22845 22389 22879 22423
rect 28273 22389 28307 22423
rect 31585 22389 31619 22423
rect 35081 22389 35115 22423
rect 39865 22389 39899 22423
rect 3249 22185 3283 22219
rect 8953 22185 8987 22219
rect 14933 22185 14967 22219
rect 18705 22185 18739 22219
rect 19441 22185 19475 22219
rect 22109 22185 22143 22219
rect 24409 22185 24443 22219
rect 29009 22185 29043 22219
rect 32505 22185 32539 22219
rect 33149 22185 33183 22219
rect 16129 22117 16163 22151
rect 6837 22049 6871 22083
rect 12357 22049 12391 22083
rect 1869 21981 1903 22015
rect 3801 21981 3835 22015
rect 6193 21981 6227 22015
rect 6377 21981 6411 22015
rect 6469 21981 6503 22015
rect 6561 21981 6595 22015
rect 7297 21981 7331 22015
rect 7481 21981 7515 22015
rect 7573 21981 7607 22015
rect 7665 21981 7699 22015
rect 9873 21981 9907 22015
rect 10149 21981 10183 22015
rect 10241 21981 10275 22015
rect 11621 21981 11655 22015
rect 12173 21981 12207 22015
rect 16313 21981 16347 22015
rect 16405 21981 16439 22015
rect 17233 21981 17267 22015
rect 17325 21981 17359 22015
rect 17417 21981 17451 22015
rect 17601 21981 17635 22015
rect 18061 21981 18095 22015
rect 18245 21981 18279 22015
rect 18337 21981 18371 22015
rect 18475 21981 18509 22015
rect 19533 21981 19567 22015
rect 19625 21981 19659 22015
rect 23305 21981 23339 22015
rect 23394 21981 23428 22015
rect 23489 21981 23523 22015
rect 23673 21981 23707 22015
rect 27629 21981 27663 22015
rect 31953 21981 31987 22015
rect 32229 21981 32263 22015
rect 32321 21981 32355 22015
rect 33149 21981 33183 22015
rect 33241 21981 33275 22015
rect 33425 21981 33459 22015
rect 36001 21981 36035 22015
rect 36093 21981 36127 22015
rect 36369 21981 36403 22015
rect 39313 21981 39347 22015
rect 40141 21981 40175 22015
rect 40230 21978 40264 22012
rect 40325 21981 40359 22015
rect 40509 21981 40543 22015
rect 2136 21913 2170 21947
rect 4046 21913 4080 21947
rect 10057 21913 10091 21947
rect 20821 21913 20855 21947
rect 27874 21913 27908 21947
rect 32137 21913 32171 21947
rect 36185 21913 36219 21947
rect 5181 21845 5215 21879
rect 7941 21845 7975 21879
rect 10425 21845 10459 21879
rect 15669 21845 15703 21879
rect 16957 21845 16991 21879
rect 19257 21845 19291 21879
rect 20269 21845 20303 21879
rect 23029 21845 23063 21879
rect 26893 21845 26927 21879
rect 32965 21845 32999 21879
rect 35817 21845 35851 21879
rect 39865 21845 39899 21879
rect 2053 21641 2087 21675
rect 3709 21641 3743 21675
rect 6377 21641 6411 21675
rect 27629 21641 27663 21675
rect 29561 21641 29595 21675
rect 32781 21641 32815 21675
rect 4905 21573 4939 21607
rect 7512 21573 7546 21607
rect 8309 21573 8343 21607
rect 10149 21573 10183 21607
rect 15761 21573 15795 21607
rect 16948 21573 16982 21607
rect 21005 21573 21039 21607
rect 23314 21573 23348 21607
rect 33241 21573 33275 21607
rect 39712 21573 39746 21607
rect 2329 21505 2363 21539
rect 2421 21505 2455 21539
rect 2513 21505 2547 21539
rect 2697 21505 2731 21539
rect 3985 21505 4019 21539
rect 4077 21505 4111 21539
rect 4169 21505 4203 21539
rect 4353 21505 4387 21539
rect 9873 21505 9907 21539
rect 10057 21505 10091 21539
rect 10241 21505 10275 21539
rect 15393 21505 15427 21539
rect 15486 21505 15520 21539
rect 15669 21505 15703 21539
rect 15899 21505 15933 21539
rect 16681 21505 16715 21539
rect 21189 21505 21223 21539
rect 27905 21505 27939 21539
rect 27997 21505 28031 21539
rect 28089 21505 28123 21539
rect 28273 21505 28307 21539
rect 28917 21505 28951 21539
rect 29745 21505 29779 21539
rect 30021 21505 30055 21539
rect 32965 21505 32999 21539
rect 7757 21437 7791 21471
rect 23581 21437 23615 21471
rect 29101 21437 29135 21471
rect 29837 21437 29871 21471
rect 33057 21437 33091 21471
rect 39957 21437 39991 21471
rect 16037 21369 16071 21403
rect 20453 21369 20487 21403
rect 3249 21301 3283 21335
rect 10425 21301 10459 21335
rect 14289 21301 14323 21335
rect 18061 21301 18095 21335
rect 22201 21301 22235 21335
rect 27169 21301 27203 21335
rect 29745 21301 29779 21335
rect 32965 21301 32999 21335
rect 35909 21301 35943 21335
rect 38577 21301 38611 21335
rect 58173 21301 58207 21335
rect 6377 21097 6411 21131
rect 10609 21097 10643 21131
rect 15853 21097 15887 21131
rect 17601 21097 17635 21131
rect 22293 21097 22327 21131
rect 6929 21029 6963 21063
rect 8125 21029 8159 21063
rect 11621 21029 11655 21063
rect 12449 21029 12483 21063
rect 20269 21029 20303 21063
rect 14749 20961 14783 20995
rect 29009 20961 29043 20995
rect 6009 20893 6043 20927
rect 6193 20893 6227 20927
rect 11805 20893 11839 20927
rect 13001 20893 13035 20927
rect 14565 20893 14599 20927
rect 17785 20893 17819 20927
rect 22759 20893 22793 20927
rect 22916 20887 22950 20921
rect 23016 20890 23050 20924
rect 23121 20893 23155 20927
rect 24777 20893 24811 20927
rect 26617 20893 26651 20927
rect 27353 20893 27387 20927
rect 8309 20825 8343 20859
rect 9873 20825 9907 20859
rect 10701 20825 10735 20859
rect 13185 20825 13219 20859
rect 17141 20825 17175 20859
rect 17969 20825 18003 20859
rect 20453 20825 20487 20859
rect 21925 20825 21959 20859
rect 22109 20825 22143 20859
rect 24409 20825 24443 20859
rect 24593 20825 24627 20859
rect 26372 20825 26406 20859
rect 27169 20825 27203 20859
rect 30021 20825 30055 20859
rect 13369 20757 13403 20791
rect 23397 20757 23431 20791
rect 25237 20757 25271 20791
rect 27813 20757 27847 20791
rect 28457 20757 28491 20791
rect 30113 20757 30147 20791
rect 32229 20757 32263 20791
rect 7573 20553 7607 20587
rect 11989 20553 12023 20587
rect 14013 20553 14047 20587
rect 16037 20553 16071 20587
rect 16957 20553 16991 20587
rect 22661 20553 22695 20587
rect 26985 20553 27019 20587
rect 29745 20553 29779 20587
rect 30205 20553 30239 20587
rect 37289 20553 37323 20587
rect 38301 20553 38335 20587
rect 19349 20485 19383 20519
rect 26065 20485 26099 20519
rect 30665 20485 30699 20519
rect 33057 20485 33091 20519
rect 34630 20485 34664 20519
rect 40325 20485 40359 20519
rect 4813 20417 4847 20451
rect 6837 20417 6871 20451
rect 7665 20417 7699 20451
rect 12633 20417 12667 20451
rect 12889 20417 12923 20451
rect 15209 20417 15243 20451
rect 17049 20417 17083 20451
rect 17785 20417 17819 20451
rect 17969 20417 18003 20451
rect 19160 20417 19194 20451
rect 19260 20417 19294 20451
rect 19477 20417 19511 20451
rect 19625 20417 19659 20451
rect 20264 20417 20298 20451
rect 20361 20417 20395 20451
rect 20453 20417 20487 20451
rect 20636 20417 20670 20451
rect 20729 20417 20763 20451
rect 22109 20417 22143 20451
rect 23121 20417 23155 20451
rect 23388 20417 23422 20451
rect 25881 20417 25915 20451
rect 27261 20417 27295 20451
rect 27353 20417 27387 20451
rect 27445 20417 27479 20451
rect 27629 20417 27663 20451
rect 29193 20417 29227 20451
rect 29377 20417 29411 20451
rect 29469 20417 29503 20451
rect 29561 20417 29595 20451
rect 30389 20417 30423 20451
rect 32413 20417 32447 20451
rect 32597 20417 32631 20451
rect 32689 20417 32723 20451
rect 32827 20417 32861 20451
rect 34897 20417 34931 20451
rect 36185 20417 36219 20451
rect 37473 20417 37507 20451
rect 37565 20417 37599 20451
rect 37657 20417 37691 20451
rect 37841 20417 37875 20451
rect 39425 20417 39459 20451
rect 40141 20417 40175 20451
rect 15485 20349 15519 20383
rect 30481 20349 30515 20383
rect 35909 20349 35943 20383
rect 39681 20349 39715 20383
rect 18981 20281 19015 20315
rect 8309 20213 8343 20247
rect 17601 20213 17635 20247
rect 17877 20213 17911 20247
rect 20085 20213 20119 20247
rect 24501 20213 24535 20247
rect 26249 20213 26283 20247
rect 28365 20213 28399 20247
rect 30389 20213 30423 20247
rect 33517 20213 33551 20247
rect 40509 20213 40543 20247
rect 7297 20009 7331 20043
rect 12725 20009 12759 20043
rect 15577 20009 15611 20043
rect 21833 20009 21867 20043
rect 33057 20009 33091 20043
rect 37565 20009 37599 20043
rect 40233 20009 40267 20043
rect 4629 19941 4663 19975
rect 14381 19873 14415 19907
rect 22385 19873 22419 19907
rect 29929 19873 29963 19907
rect 36553 19873 36587 19907
rect 2605 19805 2639 19839
rect 4445 19805 4479 19839
rect 9413 19805 9447 19839
rect 11529 19805 11563 19839
rect 11621 19805 11655 19839
rect 11713 19805 11747 19839
rect 11897 19805 11931 19839
rect 13001 19805 13035 19839
rect 13093 19805 13127 19839
rect 13185 19805 13219 19839
rect 13369 19805 13403 19839
rect 14105 19805 14139 19839
rect 15761 19805 15795 19839
rect 15853 19805 15887 19839
rect 19717 19805 19751 19839
rect 19810 19805 19844 19839
rect 19993 19805 20027 19839
rect 20182 19805 20216 19839
rect 21741 19805 21775 19839
rect 21925 19805 21959 19839
rect 29653 19805 29687 19839
rect 32689 19805 32723 19839
rect 32873 19805 32907 19839
rect 36277 19805 36311 19839
rect 37749 19805 37783 19839
rect 37841 19805 37875 19839
rect 38117 19805 38151 19839
rect 40509 19805 40543 19839
rect 40601 19805 40635 19839
rect 40693 19805 40727 19839
rect 40877 19805 40911 19839
rect 58173 19805 58207 19839
rect 6653 19737 6687 19771
rect 7573 19737 7607 19771
rect 9680 19737 9714 19771
rect 11253 19737 11287 19771
rect 20085 19737 20119 19771
rect 27445 19737 27479 19771
rect 37933 19737 37967 19771
rect 2421 19669 2455 19703
rect 5641 19669 5675 19703
rect 6101 19669 6135 19703
rect 8401 19669 8435 19703
rect 10793 19669 10827 19703
rect 20361 19669 20395 19703
rect 26157 19669 26191 19703
rect 27905 19669 27939 19703
rect 39221 19669 39255 19703
rect 5181 19465 5215 19499
rect 8677 19465 8711 19499
rect 11529 19465 11563 19499
rect 14197 19465 14231 19499
rect 14841 19465 14875 19499
rect 25835 19465 25869 19499
rect 26985 19465 27019 19499
rect 29009 19465 29043 19499
rect 32689 19465 32723 19499
rect 36001 19465 36035 19499
rect 41705 19465 41739 19499
rect 7113 19397 7147 19431
rect 22017 19397 22051 19431
rect 27445 19397 27479 19431
rect 28733 19397 28767 19431
rect 36369 19397 36403 19431
rect 4353 19329 4387 19363
rect 5273 19329 5307 19363
rect 8217 19329 8251 19363
rect 9045 19329 9079 19363
rect 11713 19329 11747 19363
rect 11897 19329 11931 19363
rect 14197 19329 14231 19363
rect 14381 19329 14415 19363
rect 15209 19329 15243 19363
rect 16681 19329 16715 19363
rect 16937 19329 16971 19363
rect 22201 19329 22235 19363
rect 27169 19329 27203 19363
rect 28457 19329 28491 19363
rect 28641 19329 28675 19363
rect 28825 19329 28859 19363
rect 29469 19329 29503 19363
rect 30895 19329 30929 19363
rect 31033 19329 31067 19363
rect 31125 19329 31159 19363
rect 31309 19329 31343 19363
rect 33802 19329 33836 19363
rect 34069 19329 34103 19363
rect 36185 19329 36219 19363
rect 36277 19329 36311 19363
rect 36553 19329 36587 19363
rect 37657 19329 37691 19363
rect 38117 19329 38151 19363
rect 40581 19329 40615 19363
rect 5365 19261 5399 19295
rect 6837 19261 6871 19295
rect 8125 19261 8159 19295
rect 8953 19261 8987 19295
rect 15117 19261 15151 19295
rect 25605 19261 25639 19295
rect 27261 19261 27295 19295
rect 29745 19261 29779 19295
rect 39865 19261 39899 19295
rect 40325 19261 40359 19295
rect 2881 19193 2915 19227
rect 9597 19193 9631 19227
rect 27905 19193 27939 19227
rect 4813 19125 4847 19159
rect 7849 19125 7883 19159
rect 8033 19125 8067 19159
rect 8861 19125 8895 19159
rect 10977 19125 11011 19159
rect 12633 19125 12667 19159
rect 15025 19125 15059 19159
rect 15761 19125 15795 19159
rect 18061 19125 18095 19159
rect 21833 19125 21867 19159
rect 27169 19125 27203 19159
rect 30757 19125 30791 19159
rect 3249 18921 3283 18955
rect 6285 18921 6319 18955
rect 12909 18921 12943 18955
rect 14473 18921 14507 18955
rect 16313 18921 16347 18955
rect 21695 18921 21729 18955
rect 25789 18921 25823 18955
rect 30113 18921 30147 18955
rect 30757 18921 30791 18955
rect 32965 18921 32999 18955
rect 40417 18921 40451 18955
rect 5641 18853 5675 18887
rect 31861 18853 31895 18887
rect 36093 18853 36127 18887
rect 4445 18785 4479 18819
rect 8217 18785 8251 18819
rect 10241 18785 10275 18819
rect 21925 18785 21959 18819
rect 23029 18785 23063 18819
rect 23305 18785 23339 18819
rect 24501 18785 24535 18819
rect 41889 18785 41923 18819
rect 1869 18717 1903 18751
rect 4169 18717 4203 18751
rect 12449 18717 12483 18751
rect 15853 18717 15887 18751
rect 16589 18717 16623 18751
rect 16681 18717 16715 18751
rect 16773 18717 16807 18751
rect 16957 18717 16991 18751
rect 17693 18717 17727 18751
rect 17877 18717 17911 18751
rect 17969 18717 18003 18751
rect 18061 18717 18095 18751
rect 19257 18717 19291 18751
rect 25237 18717 25271 18751
rect 25421 18717 25455 18751
rect 25605 18717 25639 18751
rect 29561 18717 29595 18751
rect 29745 18717 29779 18751
rect 29929 18717 29963 18751
rect 30757 18717 30791 18751
rect 30849 18717 30883 18751
rect 31033 18717 31067 18751
rect 32321 18717 32355 18751
rect 32500 18711 32534 18745
rect 32600 18714 32634 18748
rect 32689 18717 32723 18751
rect 36277 18717 36311 18751
rect 36461 18717 36495 18751
rect 36645 18717 36679 18751
rect 39957 18717 39991 18751
rect 40647 18717 40681 18751
rect 40785 18717 40819 18751
rect 40877 18717 40911 18751
rect 41061 18717 41095 18751
rect 41705 18717 41739 18751
rect 58173 18717 58207 18751
rect 2136 18649 2170 18683
rect 5457 18649 5491 18683
rect 6193 18649 6227 18683
rect 7950 18649 7984 18683
rect 10508 18649 10542 18683
rect 12265 18649 12299 18683
rect 18337 18649 18371 18683
rect 19502 18649 19536 18683
rect 25513 18649 25547 18683
rect 26617 18649 26651 18683
rect 27169 18649 27203 18683
rect 29837 18649 29871 18683
rect 36369 18649 36403 18683
rect 41521 18649 41555 18683
rect 3801 18581 3835 18615
rect 4261 18581 4295 18615
rect 6837 18581 6871 18615
rect 11621 18581 11655 18615
rect 12081 18581 12115 18615
rect 20637 18581 20671 18615
rect 27261 18581 27295 18615
rect 30573 18581 30607 18615
rect 2421 18377 2455 18411
rect 4537 18377 4571 18411
rect 10517 18377 10551 18411
rect 11529 18377 11563 18411
rect 26249 18377 26283 18411
rect 29653 18377 29687 18411
rect 32597 18377 32631 18411
rect 38761 18377 38795 18411
rect 6929 18309 6963 18343
rect 8401 18309 8435 18343
rect 9229 18309 9263 18343
rect 13001 18309 13035 18343
rect 17141 18309 17175 18343
rect 18613 18309 18647 18343
rect 18797 18309 18831 18343
rect 23949 18309 23983 18343
rect 30113 18309 30147 18343
rect 32229 18309 32263 18343
rect 32413 18309 32447 18343
rect 33241 18309 33275 18343
rect 34069 18309 34103 18343
rect 39896 18309 39930 18343
rect 40601 18309 40635 18343
rect 2237 18241 2271 18275
rect 3065 18241 3099 18275
rect 3249 18241 3283 18275
rect 3893 18241 3927 18275
rect 4997 18241 5031 18275
rect 7113 18241 7147 18275
rect 7251 18241 7285 18275
rect 7493 18239 7527 18273
rect 7677 18251 7711 18285
rect 8217 18241 8251 18275
rect 11805 18241 11839 18275
rect 11897 18241 11931 18275
rect 11989 18241 12023 18275
rect 12173 18241 12207 18275
rect 13461 18241 13495 18275
rect 13645 18241 13679 18275
rect 13737 18241 13771 18275
rect 13829 18241 13863 18275
rect 17325 18241 17359 18275
rect 17509 18241 17543 18275
rect 18981 18241 19015 18275
rect 20453 18241 20487 18275
rect 21097 18241 21131 18275
rect 25136 18241 25170 18275
rect 29837 18241 29871 18275
rect 33425 18241 33459 18275
rect 33885 18241 33919 18275
rect 37565 18241 37599 18275
rect 40831 18241 40865 18275
rect 40969 18241 41003 18275
rect 41061 18241 41095 18275
rect 41245 18241 41279 18275
rect 41705 18241 41739 18275
rect 2053 18173 2087 18207
rect 2881 18173 2915 18207
rect 7365 18173 7399 18207
rect 18061 18173 18095 18207
rect 20913 18173 20947 18207
rect 21281 18173 21315 18207
rect 24869 18173 24903 18207
rect 29929 18173 29963 18207
rect 37289 18173 37323 18207
rect 40141 18173 40175 18207
rect 5181 18105 5215 18139
rect 20269 18105 20303 18139
rect 22661 18105 22695 18139
rect 34253 18105 34287 18139
rect 3709 18037 3743 18071
rect 5733 18037 5767 18071
rect 6377 18037 6411 18071
rect 14105 18037 14139 18071
rect 19809 18037 19843 18071
rect 30113 18037 30147 18071
rect 33057 18037 33091 18071
rect 36369 18037 36403 18071
rect 5457 17833 5491 17867
rect 9045 17833 9079 17867
rect 10793 17833 10827 17867
rect 13553 17833 13587 17867
rect 21833 17833 21867 17867
rect 25697 17833 25731 17867
rect 30757 17833 30791 17867
rect 36737 17833 36771 17867
rect 40417 17833 40451 17867
rect 4353 17765 4387 17799
rect 24961 17765 24995 17799
rect 38025 17765 38059 17799
rect 5181 17697 5215 17731
rect 15485 17697 15519 17731
rect 23213 17697 23247 17731
rect 40877 17697 40911 17731
rect 5273 17629 5307 17663
rect 12173 17629 12207 17663
rect 12265 17629 12299 17663
rect 12357 17629 12391 17663
rect 12541 17629 12575 17663
rect 13185 17629 13219 17663
rect 15218 17629 15252 17663
rect 21005 17629 21039 17663
rect 21097 17629 21131 17663
rect 21210 17629 21244 17663
rect 21373 17629 21407 17663
rect 22946 17629 22980 17663
rect 24409 17629 24443 17663
rect 24777 17629 24811 17663
rect 25973 17629 26007 17663
rect 26065 17629 26099 17663
rect 26157 17629 26191 17663
rect 26341 17629 26375 17663
rect 30573 17629 30607 17663
rect 32505 17629 32539 17663
rect 32684 17629 32718 17663
rect 32781 17629 32815 17663
rect 32893 17629 32927 17663
rect 35633 17629 35667 17663
rect 35817 17629 35851 17663
rect 35909 17629 35943 17663
rect 36001 17629 36035 17663
rect 36921 17629 36955 17663
rect 37289 17629 37323 17663
rect 40233 17629 40267 17663
rect 13369 17561 13403 17595
rect 20729 17561 20763 17595
rect 24593 17561 24627 17595
rect 24685 17561 24719 17595
rect 37013 17561 37047 17595
rect 37105 17561 37139 17595
rect 37841 17561 37875 17595
rect 40049 17561 40083 17595
rect 4813 17493 4847 17527
rect 5917 17493 5951 17527
rect 7941 17493 7975 17527
rect 11437 17493 11471 17527
rect 11897 17493 11931 17527
rect 14105 17493 14139 17527
rect 20269 17493 20303 17527
rect 26893 17493 26927 17527
rect 31953 17493 31987 17527
rect 33149 17493 33183 17527
rect 35081 17493 35115 17527
rect 36277 17493 36311 17527
rect 4169 17289 4203 17323
rect 12265 17289 12299 17323
rect 13829 17289 13863 17323
rect 19717 17289 19751 17323
rect 25881 17289 25915 17323
rect 34713 17289 34747 17323
rect 37289 17289 37323 17323
rect 3056 17221 3090 17255
rect 11897 17221 11931 17255
rect 14197 17221 14231 17255
rect 17969 17221 18003 17255
rect 26065 17221 26099 17255
rect 33140 17221 33174 17255
rect 2789 17153 2823 17187
rect 5089 17153 5123 17187
rect 8410 17153 8444 17187
rect 8677 17153 8711 17187
rect 12081 17153 12115 17187
rect 13967 17153 14001 17187
rect 14105 17153 14139 17187
rect 14325 17153 14359 17187
rect 14473 17153 14507 17187
rect 15209 17153 15243 17187
rect 18889 17153 18923 17187
rect 20085 17153 20119 17187
rect 23029 17153 23063 17187
rect 23765 17153 23799 17187
rect 24944 17153 24978 17187
rect 25237 17153 25271 17187
rect 26249 17153 26283 17187
rect 26985 17153 27019 17187
rect 27169 17153 27203 17187
rect 32873 17153 32907 17187
rect 35826 17153 35860 17187
rect 36093 17153 36127 17187
rect 37473 17153 37507 17187
rect 37657 17153 37691 17187
rect 39221 17153 39255 17187
rect 4721 17085 4755 17119
rect 5181 17085 5215 17119
rect 14933 17085 14967 17119
rect 19993 17085 20027 17119
rect 22753 17085 22787 17119
rect 23489 17085 23523 17119
rect 25053 17085 25087 17119
rect 30757 17085 30791 17119
rect 31033 17085 31067 17119
rect 39497 17085 39531 17119
rect 16681 17017 16715 17051
rect 17417 17017 17451 17051
rect 24777 17017 24811 17051
rect 27353 17017 27387 17051
rect 34253 17017 34287 17051
rect 58173 17017 58207 17051
rect 5365 16949 5399 16983
rect 7297 16949 7331 16983
rect 19901 16949 19935 16983
rect 21281 16949 21315 16983
rect 25145 16949 25179 16983
rect 27905 16949 27939 16983
rect 8033 16745 8067 16779
rect 14933 16745 14967 16779
rect 20637 16745 20671 16779
rect 25881 16745 25915 16779
rect 38945 16745 38979 16779
rect 40325 16745 40359 16779
rect 21097 16677 21131 16711
rect 37381 16677 37415 16711
rect 5089 16609 5123 16643
rect 5273 16609 5307 16643
rect 7573 16609 7607 16643
rect 7665 16609 7699 16643
rect 8953 16609 8987 16643
rect 12541 16609 12575 16643
rect 19993 16609 20027 16643
rect 22845 16609 22879 16643
rect 27261 16609 27295 16643
rect 36001 16609 36035 16643
rect 2421 16541 2455 16575
rect 4997 16541 5031 16575
rect 7297 16541 7331 16575
rect 7481 16541 7515 16575
rect 7849 16541 7883 16575
rect 15761 16541 15795 16575
rect 15853 16541 15887 16575
rect 15945 16541 15979 16575
rect 16129 16541 16163 16575
rect 16589 16541 16623 16575
rect 16773 16541 16807 16575
rect 16865 16541 16899 16575
rect 16957 16541 16991 16575
rect 18061 16541 18095 16575
rect 18245 16541 18279 16575
rect 18337 16541 18371 16575
rect 18429 16541 18463 16575
rect 22569 16541 22603 16575
rect 27977 16541 28011 16575
rect 28086 16541 28120 16575
rect 28181 16541 28215 16575
rect 28365 16541 28399 16575
rect 31033 16541 31067 16575
rect 32781 16541 32815 16575
rect 32965 16541 32999 16575
rect 33057 16541 33091 16575
rect 33149 16541 33183 16575
rect 36268 16541 36302 16575
rect 27016 16473 27050 16507
rect 27721 16473 27755 16507
rect 30766 16473 30800 16507
rect 32321 16473 32355 16507
rect 33425 16473 33459 16507
rect 40417 16473 40451 16507
rect 2237 16405 2271 16439
rect 4629 16405 4663 16439
rect 9965 16405 9999 16439
rect 10517 16405 10551 16439
rect 11161 16405 11195 16439
rect 13001 16405 13035 16439
rect 15485 16405 15519 16439
rect 17233 16405 17267 16439
rect 18705 16405 18739 16439
rect 19441 16405 19475 16439
rect 22109 16405 22143 16439
rect 29653 16405 29687 16439
rect 3433 16201 3467 16235
rect 4353 16201 4387 16235
rect 5181 16201 5215 16235
rect 10885 16201 10919 16235
rect 12725 16201 12759 16235
rect 16681 16201 16715 16235
rect 17509 16201 17543 16235
rect 19073 16201 19107 16235
rect 20821 16201 20855 16235
rect 27169 16201 27203 16235
rect 37289 16201 37323 16235
rect 4261 16133 4295 16167
rect 11897 16133 11931 16167
rect 16129 16133 16163 16167
rect 17049 16133 17083 16167
rect 17877 16133 17911 16167
rect 19441 16133 19475 16167
rect 37657 16133 37691 16167
rect 2053 16065 2087 16099
rect 2320 16065 2354 16099
rect 10149 16065 10183 16099
rect 10333 16065 10367 16099
rect 10793 16065 10827 16099
rect 10977 16065 11011 16099
rect 11529 16065 11563 16099
rect 11622 16065 11656 16099
rect 11805 16065 11839 16099
rect 12035 16065 12069 16099
rect 12633 16065 12667 16099
rect 12817 16065 12851 16099
rect 14289 16065 14323 16099
rect 16865 16065 16899 16099
rect 17693 16065 17727 16099
rect 19257 16065 19291 16099
rect 20085 16065 20119 16099
rect 20729 16065 20763 16099
rect 20913 16065 20947 16099
rect 23029 16065 23063 16099
rect 27353 16065 27387 16099
rect 29101 16065 29135 16099
rect 29285 16065 29319 16099
rect 30757 16065 30791 16099
rect 31401 16065 31435 16099
rect 34253 16065 34287 16099
rect 37473 16065 37507 16099
rect 37565 16065 37599 16099
rect 37841 16065 37875 16099
rect 39977 16065 40011 16099
rect 40233 16065 40267 16099
rect 4537 15997 4571 16031
rect 9689 15997 9723 16031
rect 14565 15997 14599 16031
rect 19901 15997 19935 16031
rect 23305 15997 23339 16031
rect 26433 15997 26467 16031
rect 27537 15997 27571 16031
rect 30481 15997 30515 16031
rect 32505 15997 32539 16031
rect 35173 15997 35207 16031
rect 35449 15997 35483 16031
rect 10333 15929 10367 15963
rect 13829 15929 13863 15963
rect 31217 15929 31251 15963
rect 38301 15929 38335 15963
rect 3893 15861 3927 15895
rect 7113 15861 7147 15895
rect 12173 15861 12207 15895
rect 20269 15861 20303 15895
rect 22293 15861 22327 15895
rect 29469 15861 29503 15895
rect 38853 15861 38887 15895
rect 58173 15861 58207 15895
rect 2513 15657 2547 15691
rect 6837 15657 6871 15691
rect 7757 15657 7791 15691
rect 9321 15657 9355 15691
rect 12449 15657 12483 15691
rect 14289 15657 14323 15691
rect 21281 15657 21315 15691
rect 22477 15657 22511 15691
rect 23305 15657 23339 15691
rect 27077 15657 27111 15691
rect 29561 15657 29595 15691
rect 32597 15657 32631 15691
rect 36921 15657 36955 15691
rect 41797 15657 41831 15691
rect 7389 15589 7423 15623
rect 9965 15589 9999 15623
rect 6837 15521 6871 15555
rect 11069 15521 11103 15555
rect 19257 15521 19291 15555
rect 23765 15521 23799 15555
rect 35725 15521 35759 15555
rect 40417 15521 40451 15555
rect 2237 15453 2271 15487
rect 2329 15453 2363 15487
rect 6929 15453 6963 15487
rect 7665 15453 7699 15487
rect 7757 15453 7791 15487
rect 9413 15453 9447 15487
rect 9505 15453 9539 15487
rect 10144 15453 10178 15487
rect 10241 15453 10275 15487
rect 10516 15453 10550 15487
rect 10609 15453 10643 15487
rect 11336 15453 11370 15487
rect 12909 15453 12943 15487
rect 13002 15453 13036 15487
rect 13185 15453 13219 15487
rect 13415 15453 13449 15487
rect 14105 15453 14139 15487
rect 14289 15453 14323 15487
rect 15117 15453 15151 15487
rect 15384 15453 15418 15487
rect 19513 15453 19547 15487
rect 21097 15453 21131 15487
rect 21281 15453 21315 15487
rect 22477 15453 22511 15487
rect 22661 15453 22695 15487
rect 23121 15453 23155 15487
rect 23305 15453 23339 15487
rect 24409 15453 24443 15487
rect 26985 15453 27019 15487
rect 27169 15453 27203 15487
rect 30941 15453 30975 15487
rect 31677 15453 31711 15487
rect 31769 15453 31803 15487
rect 31861 15453 31895 15487
rect 32045 15453 32079 15487
rect 33333 15453 33367 15487
rect 33609 15453 33643 15487
rect 35449 15453 35483 15487
rect 37381 15453 37415 15487
rect 38209 15453 38243 15487
rect 38372 15450 38406 15484
rect 38485 15453 38519 15487
rect 38623 15453 38657 15487
rect 40693 15453 40727 15487
rect 41153 15453 41187 15487
rect 41337 15453 41371 15487
rect 41429 15453 41463 15487
rect 41521 15453 41555 15487
rect 10333 15385 10367 15419
rect 13277 15385 13311 15419
rect 27629 15385 27663 15419
rect 30696 15385 30730 15419
rect 31401 15385 31435 15419
rect 37565 15385 37599 15419
rect 37749 15385 37783 15419
rect 6561 15317 6595 15351
rect 9137 15317 9171 15351
rect 13553 15317 13587 15351
rect 16497 15317 16531 15351
rect 18429 15317 18463 15351
rect 20637 15317 20671 15351
rect 21925 15317 21959 15351
rect 38853 15317 38887 15351
rect 7757 15113 7791 15147
rect 18797 15113 18831 15147
rect 24225 15113 24259 15147
rect 25053 15113 25087 15147
rect 28273 15113 28307 15147
rect 29929 15113 29963 15147
rect 37473 15113 37507 15147
rect 40233 15113 40267 15147
rect 8892 15045 8926 15079
rect 9597 15045 9631 15079
rect 14289 15045 14323 15079
rect 17132 15045 17166 15079
rect 19441 15045 19475 15079
rect 22661 15045 22695 15079
rect 39098 15045 39132 15079
rect 2145 14977 2179 15011
rect 3045 14977 3079 15011
rect 5641 14977 5675 15011
rect 6377 14977 6411 15011
rect 6561 14977 6595 15011
rect 6653 14977 6687 15011
rect 6929 14977 6963 15011
rect 9137 14977 9171 15011
rect 9781 14977 9815 15011
rect 10149 14977 10183 15011
rect 10333 14977 10367 15011
rect 14105 14977 14139 15011
rect 18705 14977 18739 15011
rect 18889 14977 18923 15011
rect 20453 14977 20487 15011
rect 22569 14977 22603 15011
rect 22753 14977 22787 15011
rect 23213 14977 23247 15011
rect 23397 14977 23431 15011
rect 27537 14977 27571 15011
rect 27721 14977 27755 15011
rect 30205 14977 30239 15011
rect 30297 14977 30331 15011
rect 30389 14977 30423 15011
rect 30573 14977 30607 15011
rect 35357 14977 35391 15011
rect 36001 14977 36035 15011
rect 37289 14977 37323 15011
rect 37473 14977 37507 15011
rect 37933 14977 37967 15011
rect 40969 14977 41003 15011
rect 1961 14909 1995 14943
rect 2789 14909 2823 14943
rect 5181 14909 5215 14943
rect 5549 14909 5583 14943
rect 6745 14909 6779 14943
rect 9965 14909 9999 14943
rect 10057 14909 10091 14943
rect 16865 14909 16899 14943
rect 20177 14909 20211 14943
rect 35081 14909 35115 14943
rect 35817 14909 35851 14943
rect 36645 14909 36679 14943
rect 38853 14909 38887 14943
rect 18245 14841 18279 14875
rect 23397 14841 23431 14875
rect 2329 14773 2363 14807
rect 4169 14773 4203 14807
rect 5825 14773 5859 14807
rect 7113 14773 7147 14807
rect 14749 14773 14783 14807
rect 22109 14773 22143 14807
rect 27353 14773 27387 14807
rect 29469 14773 29503 14807
rect 31217 14773 31251 14807
rect 33241 14773 33275 14807
rect 36185 14773 36219 14807
rect 2789 14569 2823 14603
rect 10425 14569 10459 14603
rect 16681 14569 16715 14603
rect 18613 14569 18647 14603
rect 20913 14569 20947 14603
rect 23397 14569 23431 14603
rect 24593 14569 24627 14603
rect 30205 14569 30239 14603
rect 40233 14569 40267 14603
rect 4537 14501 4571 14535
rect 6377 14501 6411 14535
rect 22385 14501 22419 14535
rect 40969 14501 41003 14535
rect 4997 14433 5031 14467
rect 5181 14433 5215 14467
rect 17141 14433 17175 14467
rect 19533 14433 19567 14467
rect 24685 14433 24719 14467
rect 28365 14433 28399 14467
rect 33517 14433 33551 14467
rect 33793 14433 33827 14467
rect 34713 14433 34747 14467
rect 36001 14433 36035 14467
rect 2605 14365 2639 14399
rect 7490 14365 7524 14399
rect 7757 14365 7791 14399
rect 10241 14365 10275 14399
rect 10425 14365 10459 14399
rect 11989 14365 12023 14399
rect 16497 14365 16531 14399
rect 16681 14365 16715 14399
rect 19441 14365 19475 14399
rect 19625 14365 19659 14399
rect 20177 14365 20211 14399
rect 20361 14365 20395 14399
rect 20821 14365 20855 14399
rect 21005 14365 21039 14399
rect 21833 14365 21867 14399
rect 22017 14365 22051 14399
rect 22201 14365 22235 14399
rect 22845 14365 22879 14399
rect 23029 14365 23063 14399
rect 23121 14365 23155 14399
rect 23213 14365 23247 14399
rect 24593 14365 24627 14399
rect 24869 14365 24903 14399
rect 26801 14365 26835 14399
rect 27537 14365 27571 14399
rect 27629 14365 27663 14399
rect 27721 14365 27755 14399
rect 27905 14365 27939 14399
rect 28733 14365 28767 14399
rect 29837 14365 29871 14399
rect 34989 14365 35023 14399
rect 36185 14365 36219 14399
rect 37197 14365 37231 14399
rect 40049 14365 40083 14399
rect 40785 14365 40819 14399
rect 58173 14365 58207 14399
rect 22109 14297 22143 14331
rect 26556 14297 26590 14331
rect 27261 14297 27295 14331
rect 28549 14297 28583 14331
rect 30021 14297 30055 14331
rect 39865 14297 39899 14331
rect 4905 14229 4939 14263
rect 5825 14229 5859 14263
rect 9689 14229 9723 14263
rect 10885 14229 10919 14263
rect 12081 14229 12115 14263
rect 15945 14229 15979 14263
rect 24409 14229 24443 14263
rect 25421 14229 25455 14263
rect 36369 14229 36403 14263
rect 38485 14229 38519 14263
rect 2973 14025 3007 14059
rect 19349 14025 19383 14059
rect 20729 14025 20763 14059
rect 22109 14025 22143 14059
rect 23673 14025 23707 14059
rect 24593 14025 24627 14059
rect 25605 14025 25639 14059
rect 26433 14025 26467 14059
rect 28365 14025 28399 14059
rect 22753 13957 22787 13991
rect 22845 13957 22879 13991
rect 24133 13957 24167 13991
rect 36553 13957 36587 13991
rect 39221 13957 39255 13991
rect 3157 13889 3191 13923
rect 7297 13889 7331 13923
rect 14298 13889 14332 13923
rect 14565 13889 14599 13923
rect 22569 13889 22603 13923
rect 22937 13889 22971 13923
rect 23857 13889 23891 13923
rect 24777 13889 24811 13923
rect 25053 13889 25087 13923
rect 26985 13889 27019 13923
rect 27252 13889 27286 13923
rect 30674 13889 30708 13923
rect 30941 13889 30975 13923
rect 33977 13889 34011 13923
rect 34437 13889 34471 13923
rect 34621 13889 34655 13923
rect 35909 13889 35943 13923
rect 36737 13889 36771 13923
rect 38577 13889 38611 13923
rect 23949 13821 23983 13855
rect 24869 13821 24903 13855
rect 35633 13821 35667 13855
rect 38301 13821 38335 13855
rect 23121 13753 23155 13787
rect 29561 13753 29595 13787
rect 34529 13753 34563 13787
rect 7757 13685 7791 13719
rect 13185 13685 13219 13719
rect 18705 13685 18739 13719
rect 19901 13685 19935 13719
rect 23857 13685 23891 13719
rect 24961 13685 24995 13719
rect 36369 13685 36403 13719
rect 39313 13685 39347 13719
rect 14289 13481 14323 13515
rect 27261 13481 27295 13515
rect 29009 13481 29043 13515
rect 30297 13481 30331 13515
rect 34989 13481 35023 13515
rect 36829 13481 36863 13515
rect 19349 13413 19383 13447
rect 22201 13413 22235 13447
rect 23581 13345 23615 13379
rect 28365 13345 28399 13379
rect 34161 13345 34195 13379
rect 35449 13345 35483 13379
rect 37749 13345 37783 13379
rect 5917 13277 5951 13311
rect 7665 13277 7699 13311
rect 9689 13277 9723 13311
rect 13553 13277 13587 13311
rect 14565 13277 14599 13311
rect 14657 13277 14691 13311
rect 14749 13277 14783 13311
rect 14933 13277 14967 13311
rect 17785 13277 17819 13311
rect 19993 13277 20027 13311
rect 23857 13277 23891 13311
rect 24777 13277 24811 13311
rect 27537 13277 27571 13311
rect 27629 13277 27663 13311
rect 27721 13277 27755 13311
rect 27905 13277 27939 13311
rect 29653 13277 29687 13311
rect 29837 13277 29871 13311
rect 29929 13277 29963 13311
rect 30021 13277 30055 13311
rect 30849 13277 30883 13311
rect 38209 13277 38243 13311
rect 38393 13277 38427 13311
rect 38485 13277 38519 13311
rect 38577 13277 38611 13311
rect 39865 13277 39899 13311
rect 58173 13277 58207 13311
rect 9934 13209 9968 13243
rect 17601 13209 17635 13243
rect 20177 13209 20211 13243
rect 24961 13209 24995 13243
rect 25513 13209 25547 13243
rect 31033 13209 31067 13243
rect 33894 13209 33928 13243
rect 35694 13209 35728 13243
rect 37381 13209 37415 13243
rect 37565 13209 37599 13243
rect 8217 13141 8251 13175
rect 11069 13141 11103 13175
rect 17969 13141 18003 13175
rect 18705 13141 18739 13175
rect 21189 13141 21223 13175
rect 26801 13141 26835 13175
rect 32781 13141 32815 13175
rect 38853 13141 38887 13175
rect 4997 12937 5031 12971
rect 6745 12937 6779 12971
rect 10149 12937 10183 12971
rect 14105 12937 14139 12971
rect 15853 12937 15887 12971
rect 20085 12937 20119 12971
rect 23949 12937 23983 12971
rect 29745 12937 29779 12971
rect 30665 12937 30699 12971
rect 32229 12937 32263 12971
rect 33333 12937 33367 12971
rect 35449 12937 35483 12971
rect 39865 12937 39899 12971
rect 9597 12869 9631 12903
rect 20913 12869 20947 12903
rect 26157 12869 26191 12903
rect 29377 12869 29411 12903
rect 29561 12869 29595 12903
rect 38752 12869 38786 12903
rect 2513 12801 2547 12835
rect 5365 12801 5399 12835
rect 11713 12801 11747 12835
rect 12081 12801 12115 12835
rect 12265 12801 12299 12835
rect 14289 12801 14323 12835
rect 14473 12801 14507 12835
rect 14933 12801 14967 12835
rect 15117 12801 15151 12835
rect 18070 12801 18104 12835
rect 18337 12801 18371 12835
rect 19073 12801 19107 12835
rect 19165 12801 19199 12835
rect 19257 12801 19291 12835
rect 19441 12801 19475 12835
rect 19901 12801 19935 12835
rect 20729 12801 20763 12835
rect 24501 12801 24535 12835
rect 26985 12801 27019 12835
rect 32689 12801 32723 12835
rect 32873 12801 32907 12835
rect 32965 12801 32999 12835
rect 33103 12801 33137 12835
rect 35725 12801 35759 12835
rect 35817 12801 35851 12835
rect 35909 12801 35943 12835
rect 36093 12801 36127 12835
rect 37657 12801 37691 12835
rect 38485 12801 38519 12835
rect 2697 12733 2731 12767
rect 3985 12733 4019 12767
rect 4261 12733 4295 12767
rect 5457 12733 5491 12767
rect 5549 12733 5583 12767
rect 6837 12733 6871 12767
rect 6929 12733 6963 12767
rect 11897 12733 11931 12767
rect 11989 12733 12023 12767
rect 21925 12733 21959 12767
rect 22477 12733 22511 12767
rect 34069 12733 34103 12767
rect 34345 12733 34379 12767
rect 12817 12665 12851 12699
rect 16957 12665 16991 12699
rect 2329 12597 2363 12631
rect 6377 12597 6411 12631
rect 8309 12597 8343 12631
rect 11529 12597 11563 12631
rect 15301 12597 15335 12631
rect 18797 12597 18831 12631
rect 21097 12597 21131 12631
rect 37473 12597 37507 12631
rect 9689 12393 9723 12427
rect 10241 12393 10275 12427
rect 13185 12393 13219 12427
rect 22661 12393 22695 12427
rect 32873 12393 32907 12427
rect 33885 12393 33919 12427
rect 36001 12393 36035 12427
rect 35541 12325 35575 12359
rect 3801 12257 3835 12291
rect 5825 12257 5859 12291
rect 6653 12257 6687 12291
rect 6745 12257 6779 12291
rect 7849 12257 7883 12291
rect 21005 12257 21039 12291
rect 21465 12257 21499 12291
rect 30113 12257 30147 12291
rect 40141 12257 40175 12291
rect 1869 12189 1903 12223
rect 2513 12189 2547 12223
rect 2697 12189 2731 12223
rect 2881 12189 2915 12223
rect 6377 12189 6411 12223
rect 6565 12189 6599 12223
rect 6929 12189 6963 12223
rect 7573 12189 7607 12223
rect 8941 12189 8975 12223
rect 9137 12189 9171 12223
rect 9229 12189 9263 12223
rect 9321 12189 9355 12223
rect 9505 12189 9539 12223
rect 12274 12189 12308 12223
rect 12541 12189 12575 12223
rect 13001 12189 13035 12223
rect 14933 12189 14967 12223
rect 15025 12189 15059 12223
rect 15117 12189 15151 12223
rect 15301 12189 15335 12223
rect 18317 12189 18351 12223
rect 18429 12183 18463 12217
rect 18521 12189 18555 12223
rect 18705 12189 18739 12223
rect 19257 12189 19291 12223
rect 19441 12189 19475 12223
rect 20729 12189 20763 12223
rect 21721 12189 21755 12223
rect 21830 12186 21864 12220
rect 21930 12189 21964 12223
rect 22109 12189 22143 12223
rect 25053 12189 25087 12223
rect 28365 12189 28399 12223
rect 30573 12189 30607 12223
rect 30757 12189 30791 12223
rect 30849 12189 30883 12223
rect 30941 12189 30975 12223
rect 35357 12189 35391 12223
rect 38301 12189 38335 12223
rect 38577 12189 38611 12223
rect 39865 12189 39899 12223
rect 4046 12121 4080 12155
rect 15853 12121 15887 12155
rect 18061 12121 18095 12155
rect 19625 12121 19659 12155
rect 25298 12121 25332 12155
rect 27537 12121 27571 12155
rect 28181 12121 28215 12155
rect 32505 12121 32539 12155
rect 32689 12121 32723 12155
rect 2053 12053 2087 12087
rect 5181 12053 5215 12087
rect 7113 12053 7147 12087
rect 11161 12053 11195 12087
rect 14197 12053 14231 12087
rect 14657 12053 14691 12087
rect 17141 12053 17175 12087
rect 26433 12053 26467 12087
rect 27445 12053 27479 12087
rect 31217 12053 31251 12087
rect 5825 11849 5859 11883
rect 14105 11849 14139 11883
rect 17141 11849 17175 11883
rect 19901 11849 19935 11883
rect 23305 11849 23339 11883
rect 25145 11849 25179 11883
rect 28273 11849 28307 11883
rect 30481 11849 30515 11883
rect 35265 11849 35299 11883
rect 39957 11849 39991 11883
rect 6837 11781 6871 11815
rect 8502 11781 8536 11815
rect 21036 11781 21070 11815
rect 24593 11781 24627 11815
rect 35541 11781 35575 11815
rect 40417 11781 40451 11815
rect 40601 11781 40635 11815
rect 2145 11713 2179 11747
rect 2789 11713 2823 11747
rect 3045 11713 3079 11747
rect 5549 11713 5583 11747
rect 8769 11713 8803 11747
rect 12081 11713 12115 11747
rect 13277 11713 13311 11747
rect 13369 11713 13403 11747
rect 13461 11713 13495 11747
rect 13645 11713 13679 11747
rect 15218 11713 15252 11747
rect 15485 11713 15519 11747
rect 18265 11713 18299 11747
rect 18521 11713 18555 11747
rect 19257 11713 19291 11747
rect 22201 11713 22235 11747
rect 22293 11713 22327 11747
rect 22385 11713 22419 11747
rect 22569 11713 22603 11747
rect 25421 11713 25455 11747
rect 25513 11713 25547 11747
rect 25605 11713 25639 11747
rect 25789 11713 25823 11747
rect 28089 11713 28123 11747
rect 30113 11713 30147 11747
rect 30297 11713 30331 11747
rect 30941 11713 30975 11747
rect 31125 11713 31159 11747
rect 31217 11713 31251 11747
rect 31355 11713 31389 11747
rect 32965 11713 32999 11747
rect 35449 11713 35483 11747
rect 35633 11713 35667 11747
rect 35817 11713 35851 11747
rect 38833 11713 38867 11747
rect 5181 11645 5215 11679
rect 5641 11645 5675 11679
rect 12357 11645 12391 11679
rect 21281 11645 21315 11679
rect 32689 11645 32723 11679
rect 38577 11645 38611 11679
rect 2329 11577 2363 11611
rect 7389 11577 7423 11611
rect 58173 11577 58207 11611
rect 4169 11509 4203 11543
rect 13001 11509 13035 11543
rect 16037 11509 16071 11543
rect 19349 11509 19383 11543
rect 21925 11509 21959 11543
rect 24133 11509 24167 11543
rect 31585 11509 31619 11543
rect 40785 11509 40819 11543
rect 15945 11305 15979 11339
rect 18705 11305 18739 11339
rect 19257 11305 19291 11339
rect 20177 11305 20211 11339
rect 25881 11305 25915 11339
rect 32505 11305 32539 11339
rect 38117 11305 38151 11339
rect 38669 11305 38703 11339
rect 15485 11237 15519 11271
rect 21189 11237 21223 11271
rect 6469 11169 6503 11203
rect 14105 11169 14139 11203
rect 21649 11169 21683 11203
rect 23857 11169 23891 11203
rect 36461 11169 36495 11203
rect 6193 11101 6227 11135
rect 10333 11101 10367 11135
rect 14361 11101 14395 11135
rect 16129 11101 16163 11135
rect 16313 11101 16347 11135
rect 20361 11101 20395 11135
rect 21916 11101 21950 11135
rect 23673 11101 23707 11135
rect 24777 11101 24811 11135
rect 24961 11101 24995 11135
rect 25053 11101 25087 11135
rect 25145 11101 25179 11135
rect 26065 11101 26099 11135
rect 28365 11101 28399 11135
rect 31125 11101 31159 11135
rect 35633 11101 35667 11135
rect 35725 11101 35759 11135
rect 35817 11101 35851 11135
rect 36001 11101 36035 11135
rect 36645 11101 36679 11135
rect 37657 11101 37691 11135
rect 38945 11101 38979 11135
rect 39037 11101 39071 11135
rect 39129 11101 39163 11135
rect 39313 11101 39347 11135
rect 10149 11033 10183 11067
rect 21005 11033 21039 11067
rect 26249 11033 26283 11067
rect 28549 11033 28583 11067
rect 31392 11033 31426 11067
rect 34897 11033 34931 11067
rect 36829 11033 36863 11067
rect 9413 10965 9447 10999
rect 23029 10965 23063 10999
rect 23489 10965 23523 10999
rect 25421 10965 25455 10999
rect 30665 10965 30699 10999
rect 35357 10965 35391 10999
rect 6377 10761 6411 10795
rect 8861 10761 8895 10795
rect 12173 10761 12207 10795
rect 22201 10761 22235 10795
rect 27445 10761 27479 10795
rect 31585 10761 31619 10795
rect 36645 10761 36679 10795
rect 38393 10761 38427 10795
rect 9781 10693 9815 10727
rect 17325 10693 17359 10727
rect 22569 10693 22603 10727
rect 25320 10693 25354 10727
rect 28641 10693 28675 10727
rect 33250 10693 33284 10727
rect 5457 10625 5491 10659
rect 6561 10625 6595 10659
rect 7021 10625 7055 10659
rect 11897 10625 11931 10659
rect 17141 10625 17175 10659
rect 22385 10625 22419 10659
rect 23029 10625 23063 10659
rect 23213 10625 23247 10659
rect 24317 10625 24351 10659
rect 25053 10625 25087 10659
rect 27997 10625 28031 10659
rect 31217 10625 31251 10659
rect 31401 10625 31435 10659
rect 35521 10625 35555 10659
rect 37933 10625 37967 10659
rect 39221 10625 39255 10659
rect 39313 10625 39347 10659
rect 39405 10625 39439 10659
rect 39589 10625 39623 10659
rect 6653 10557 6687 10591
rect 8677 10557 8711 10591
rect 9045 10557 9079 10591
rect 11529 10557 11563 10591
rect 11989 10557 12023 10591
rect 24593 10557 24627 10591
rect 33517 10557 33551 10591
rect 35265 10557 35299 10591
rect 5641 10489 5675 10523
rect 23121 10489 23155 10523
rect 9229 10421 9263 10455
rect 18981 10421 19015 10455
rect 20821 10421 20855 10455
rect 26433 10421 26467 10455
rect 28181 10421 28215 10455
rect 29929 10421 29963 10455
rect 32137 10421 32171 10455
rect 34805 10421 34839 10455
rect 38945 10421 38979 10455
rect 58173 10421 58207 10455
rect 16497 10217 16531 10251
rect 22845 10217 22879 10251
rect 25237 10217 25271 10251
rect 28273 10217 28307 10251
rect 29009 10217 29043 10251
rect 38577 10217 38611 10251
rect 4997 10149 5031 10183
rect 9965 10149 9999 10183
rect 5641 10081 5675 10115
rect 10425 10081 10459 10115
rect 10609 10081 10643 10115
rect 2697 10013 2731 10047
rect 2881 10013 2915 10047
rect 6285 10013 6319 10047
rect 8953 10013 8987 10047
rect 24593 10013 24627 10047
rect 25421 10013 25455 10047
rect 27721 10013 27755 10047
rect 27997 10013 28031 10047
rect 28089 10013 28123 10047
rect 29837 10013 29871 10047
rect 29929 10013 29963 10047
rect 30021 10013 30055 10047
rect 30205 10013 30239 10047
rect 36645 10013 36679 10047
rect 37105 10013 37139 10047
rect 5365 9945 5399 9979
rect 6469 9945 6503 9979
rect 16589 9945 16623 9979
rect 25605 9945 25639 9979
rect 27905 9945 27939 9979
rect 2513 9877 2547 9911
rect 5457 9877 5491 9911
rect 9137 9877 9171 9911
rect 10333 9877 10367 9911
rect 11161 9877 11195 9911
rect 24777 9877 24811 9911
rect 29561 9877 29595 9911
rect 1869 9673 1903 9707
rect 8401 9673 8435 9707
rect 10241 9673 10275 9707
rect 29929 9673 29963 9707
rect 2574 9605 2608 9639
rect 4537 9605 4571 9639
rect 7297 9605 7331 9639
rect 9128 9605 9162 9639
rect 20729 9605 20763 9639
rect 22753 9605 22787 9639
rect 25605 9605 25639 9639
rect 25697 9605 25731 9639
rect 29561 9605 29595 9639
rect 31585 9605 31619 9639
rect 35449 9605 35483 9639
rect 37565 9605 37599 9639
rect 37933 9605 37967 9639
rect 38660 9605 38694 9639
rect 1685 9537 1719 9571
rect 4905 9537 4939 9571
rect 8217 9537 8251 9571
rect 13369 9537 13403 9571
rect 14197 9537 14231 9571
rect 18337 9537 18371 9571
rect 22477 9537 22511 9571
rect 22661 9537 22695 9571
rect 22845 9537 22879 9571
rect 25421 9537 25455 9571
rect 25789 9537 25823 9571
rect 29745 9537 29779 9571
rect 32137 9537 32171 9571
rect 32321 9537 32355 9571
rect 32413 9537 32447 9571
rect 32505 9537 32539 9571
rect 35633 9537 35667 9571
rect 37749 9537 37783 9571
rect 2329 9469 2363 9503
rect 4997 9469 5031 9503
rect 8033 9469 8067 9503
rect 8861 9469 8895 9503
rect 13461 9469 13495 9503
rect 13553 9469 13587 9503
rect 28273 9469 28307 9503
rect 28549 9469 28583 9503
rect 30389 9469 30423 9503
rect 38393 9469 38427 9503
rect 3709 9401 3743 9435
rect 23029 9401 23063 9435
rect 25973 9401 26007 9435
rect 39773 9401 39807 9435
rect 5181 9333 5215 9367
rect 6469 9333 6503 9367
rect 7389 9333 7423 9367
rect 10701 9333 10735 9367
rect 12541 9333 12575 9367
rect 13001 9333 13035 9367
rect 14381 9333 14415 9367
rect 15301 9333 15335 9367
rect 15853 9333 15887 9367
rect 16773 9333 16807 9367
rect 17877 9333 17911 9367
rect 18521 9333 18555 9367
rect 32781 9333 32815 9367
rect 35265 9333 35299 9367
rect 7481 9129 7515 9163
rect 10241 9129 10275 9163
rect 20637 9129 20671 9163
rect 28917 9129 28951 9163
rect 32689 9129 32723 9163
rect 33701 9129 33735 9163
rect 36093 9129 36127 9163
rect 4721 9061 4755 9095
rect 13369 9061 13403 9095
rect 16129 9061 16163 9095
rect 18705 9061 18739 9095
rect 2513 8993 2547 9027
rect 5457 8993 5491 9027
rect 9229 8993 9263 9027
rect 9321 8993 9355 9027
rect 13001 8993 13035 9027
rect 15485 8993 15519 9027
rect 17325 8993 17359 9027
rect 21189 8993 21223 9027
rect 21925 8993 21959 9027
rect 22201 8993 22235 9027
rect 34713 8993 34747 9027
rect 2329 8925 2363 8959
rect 5181 8925 5215 8959
rect 6929 8925 6963 8959
rect 8953 8925 8987 8959
rect 9137 8925 9171 8959
rect 9505 8925 9539 8959
rect 11161 8925 11195 8959
rect 11345 8925 11379 8959
rect 11437 8925 11471 8959
rect 11529 8925 11563 8959
rect 11713 8925 11747 8959
rect 13185 8925 13219 8959
rect 15218 8925 15252 8959
rect 15945 8925 15979 8959
rect 19257 8925 19291 8959
rect 21097 8925 21131 8959
rect 21281 8925 21315 8959
rect 28365 8925 28399 8959
rect 28733 8925 28767 8959
rect 32137 8925 32171 8959
rect 32413 8925 32447 8959
rect 32505 8925 32539 8959
rect 33149 8925 33183 8959
rect 33425 8925 33459 8959
rect 33517 8925 33551 8959
rect 37933 8925 37967 8959
rect 58173 8925 58207 8959
rect 4537 8857 4571 8891
rect 17570 8857 17604 8891
rect 19502 8857 19536 8891
rect 28549 8857 28583 8891
rect 28641 8857 28675 8891
rect 29929 8857 29963 8891
rect 32321 8857 32355 8891
rect 33333 8857 33367 8891
rect 34980 8857 35014 8891
rect 37105 8857 37139 8891
rect 37289 8857 37323 8891
rect 38178 8857 38212 8891
rect 1593 8789 1627 8823
rect 2145 8789 2179 8823
rect 3065 8789 3099 8823
rect 3893 8789 3927 8823
rect 6745 8789 6779 8823
rect 8033 8789 8067 8823
rect 9689 8789 9723 8823
rect 11897 8789 11931 8823
rect 14105 8789 14139 8823
rect 16681 8789 16715 8823
rect 23397 8789 23431 8823
rect 31217 8789 31251 8823
rect 37473 8789 37507 8823
rect 39313 8789 39347 8823
rect 1685 8585 1719 8619
rect 7021 8585 7055 8619
rect 12173 8585 12207 8619
rect 17325 8585 17359 8619
rect 19073 8585 19107 8619
rect 27721 8585 27755 8619
rect 29561 8585 29595 8619
rect 32873 8585 32907 8619
rect 34897 8585 34931 8619
rect 38025 8585 38059 8619
rect 2390 8517 2424 8551
rect 9680 8517 9714 8551
rect 11529 8517 11563 8551
rect 13001 8517 13035 8551
rect 16773 8517 16807 8551
rect 19533 8517 19567 8551
rect 19717 8517 19751 8551
rect 27353 8517 27387 8551
rect 30674 8517 30708 8551
rect 32597 8517 32631 8551
rect 1501 8449 1535 8483
rect 6653 8449 6687 8483
rect 6837 8449 6871 8483
rect 7849 8449 7883 8483
rect 9413 8449 9447 8483
rect 11897 8449 11931 8483
rect 14013 8449 14047 8483
rect 14749 8449 14783 8483
rect 17555 8449 17589 8483
rect 17693 8449 17727 8483
rect 17785 8449 17819 8483
rect 17969 8449 18003 8483
rect 18429 8449 18463 8483
rect 18613 8449 18647 8483
rect 18705 8449 18739 8483
rect 18797 8449 18831 8483
rect 19901 8449 19935 8483
rect 21833 8449 21867 8483
rect 22109 8449 22143 8483
rect 23765 8449 23799 8483
rect 23857 8449 23891 8483
rect 23949 8449 23983 8483
rect 24133 8449 24167 8483
rect 27169 8449 27203 8483
rect 27445 8449 27479 8483
rect 27537 8449 27571 8483
rect 28457 8449 28491 8483
rect 32321 8449 32355 8483
rect 32505 8449 32539 8483
rect 32689 8449 32723 8483
rect 35173 8449 35207 8483
rect 35265 8449 35299 8483
rect 35357 8449 35391 8483
rect 35541 8449 35575 8483
rect 37381 8449 37415 8483
rect 37565 8449 37599 8483
rect 37657 8449 37691 8483
rect 37749 8449 37783 8483
rect 2145 8381 2179 8415
rect 4997 8381 5031 8415
rect 5273 8381 5307 8415
rect 7941 8381 7975 8415
rect 8033 8381 8067 8415
rect 11989 8381 12023 8415
rect 16037 8381 16071 8415
rect 21005 8381 21039 8415
rect 28181 8381 28215 8415
rect 30941 8381 30975 8415
rect 34345 8381 34379 8415
rect 7481 8313 7515 8347
rect 8769 8313 8803 8347
rect 10793 8313 10827 8347
rect 13553 8313 13587 8347
rect 15485 8313 15519 8347
rect 3525 8245 3559 8279
rect 3985 8245 4019 8279
rect 14197 8245 14231 8279
rect 14933 8245 14967 8279
rect 23489 8245 23523 8279
rect 2421 8041 2455 8075
rect 5365 8041 5399 8075
rect 7665 8041 7699 8075
rect 18337 8041 18371 8075
rect 24409 8041 24443 8075
rect 26709 8041 26743 8075
rect 29009 8041 29043 8075
rect 31585 8041 31619 8075
rect 37289 8041 37323 8075
rect 11529 7973 11563 8007
rect 2881 7905 2915 7939
rect 3065 7905 3099 7939
rect 4169 7905 4203 7939
rect 4537 7905 4571 7939
rect 19809 7905 19843 7939
rect 2789 7837 2823 7871
rect 4077 7837 4111 7871
rect 6285 7837 6319 7871
rect 6552 7837 6586 7871
rect 8217 7837 8251 7871
rect 13001 7837 13035 7871
rect 15393 7837 15427 7871
rect 23590 7837 23624 7871
rect 23857 7837 23891 7871
rect 25329 7837 25363 7871
rect 28457 7837 28491 7871
rect 28825 7837 28859 7871
rect 31401 7837 31435 7871
rect 35265 7837 35299 7871
rect 35633 7837 35667 7871
rect 58173 7837 58207 7871
rect 5273 7769 5307 7803
rect 10241 7769 10275 7803
rect 15660 7769 15694 7803
rect 17233 7769 17267 7803
rect 17785 7769 17819 7803
rect 18521 7769 18555 7803
rect 18705 7769 18739 7803
rect 19349 7769 19383 7803
rect 24593 7769 24627 7803
rect 24777 7769 24811 7803
rect 25596 7769 25630 7803
rect 28641 7769 28675 7803
rect 28733 7769 28767 7803
rect 31217 7769 31251 7803
rect 35357 7769 35391 7803
rect 35449 7769 35483 7803
rect 1869 7701 1903 7735
rect 3893 7701 3927 7735
rect 9229 7701 9263 7735
rect 9689 7701 9723 7735
rect 13553 7701 13587 7735
rect 14657 7701 14691 7735
rect 16773 7701 16807 7735
rect 20361 7701 20395 7735
rect 21649 7701 21683 7735
rect 22477 7701 22511 7735
rect 35081 7701 35115 7735
rect 10425 7497 10459 7531
rect 15577 7497 15611 7531
rect 23029 7497 23063 7531
rect 25605 7497 25639 7531
rect 28641 7497 28675 7531
rect 32505 7497 32539 7531
rect 35081 7497 35115 7531
rect 36369 7497 36403 7531
rect 38117 7497 38151 7531
rect 7573 7429 7607 7463
rect 12326 7429 12360 7463
rect 16681 7429 16715 7463
rect 16865 7429 16899 7463
rect 22753 7429 22787 7463
rect 26065 7429 26099 7463
rect 26249 7429 26283 7463
rect 30389 7429 30423 7463
rect 33618 7429 33652 7463
rect 35449 7429 35483 7463
rect 38669 7429 38703 7463
rect 3709 7361 3743 7395
rect 3985 7361 4019 7395
rect 4077 7361 4111 7395
rect 4261 7361 4295 7395
rect 5273 7361 5307 7395
rect 6561 7361 6595 7395
rect 6745 7361 6779 7395
rect 6929 7361 6963 7395
rect 7113 7361 7147 7395
rect 7941 7361 7975 7395
rect 8033 7361 8067 7395
rect 12081 7361 12115 7395
rect 14197 7361 14231 7395
rect 14933 7361 14967 7395
rect 15096 7361 15130 7395
rect 15212 7361 15246 7395
rect 15321 7361 15355 7395
rect 17049 7361 17083 7395
rect 17877 7361 17911 7395
rect 19349 7361 19383 7395
rect 20913 7361 20947 7395
rect 21097 7361 21131 7395
rect 21833 7361 21867 7395
rect 22017 7361 22051 7395
rect 22477 7361 22511 7395
rect 22661 7361 22695 7395
rect 22845 7361 22879 7395
rect 23673 7361 23707 7395
rect 23857 7361 23891 7395
rect 24961 7361 24995 7395
rect 25145 7361 25179 7395
rect 25237 7361 25271 7395
rect 25329 7361 25363 7395
rect 27517 7361 27551 7395
rect 30573 7361 30607 7395
rect 35265 7361 35299 7395
rect 35357 7361 35391 7395
rect 35633 7361 35667 7395
rect 38853 7361 38887 7395
rect 3893 7293 3927 7327
rect 6837 7293 6871 7327
rect 18153 7293 18187 7327
rect 26433 7293 26467 7327
rect 27261 7293 27295 7327
rect 33885 7293 33919 7327
rect 1961 7225 1995 7259
rect 3065 7225 3099 7259
rect 6377 7225 6411 7259
rect 8217 7225 8251 7259
rect 10977 7225 11011 7259
rect 16037 7225 16071 7259
rect 19901 7225 19935 7259
rect 24409 7225 24443 7259
rect 2513 7157 2547 7191
rect 3525 7157 3559 7191
rect 5825 7157 5859 7191
rect 8769 7157 8803 7191
rect 9873 7157 9907 7191
rect 11529 7157 11563 7191
rect 13461 7157 13495 7191
rect 14105 7157 14139 7191
rect 19165 7157 19199 7191
rect 20361 7157 20395 7191
rect 21281 7157 21315 7191
rect 21925 7157 21959 7191
rect 23489 7157 23523 7191
rect 30205 7157 30239 7191
rect 39037 7157 39071 7191
rect 4353 6953 4387 6987
rect 31309 6953 31343 6987
rect 36001 6953 36035 6987
rect 39865 6953 39899 6987
rect 13277 6885 13311 6919
rect 2697 6817 2731 6851
rect 6745 6817 6779 6851
rect 10057 6817 10091 6851
rect 11529 6817 11563 6851
rect 15485 6817 15519 6851
rect 21925 6817 21959 6851
rect 24409 6817 24443 6851
rect 25973 6817 26007 6851
rect 26249 6817 26283 6851
rect 28365 6817 28399 6851
rect 29929 6817 29963 6851
rect 2145 6749 2179 6783
rect 4997 6749 5031 6783
rect 5089 6749 5123 6783
rect 6469 6749 6503 6783
rect 7941 6749 7975 6783
rect 8953 6749 8987 6783
rect 9781 6749 9815 6783
rect 9965 6749 9999 6783
rect 10149 6749 10183 6783
rect 10333 6749 10367 6783
rect 10793 6749 10827 6783
rect 11989 6749 12023 6783
rect 12725 6749 12759 6783
rect 14427 6749 14461 6783
rect 14565 6749 14599 6783
rect 14662 6749 14696 6783
rect 14841 6749 14875 6783
rect 16037 6749 16071 6783
rect 16313 6749 16347 6783
rect 21649 6749 21683 6783
rect 23489 6749 23523 6783
rect 23581 6749 23615 6783
rect 23673 6749 23707 6783
rect 23857 6749 23891 6783
rect 24685 6749 24719 6783
rect 24777 6749 24811 6783
rect 24869 6749 24903 6783
rect 25053 6749 25087 6783
rect 27537 6749 27571 6783
rect 27629 6749 27663 6783
rect 27721 6749 27755 6783
rect 27905 6749 27939 6783
rect 28733 6749 28767 6783
rect 33793 6749 33827 6783
rect 35173 6749 35207 6783
rect 35265 6746 35299 6780
rect 35357 6749 35391 6783
rect 35541 6749 35575 6783
rect 36645 6749 36679 6783
rect 36829 6749 36863 6783
rect 36921 6749 36955 6783
rect 37013 6749 37047 6783
rect 37749 6749 37783 6783
rect 38623 6749 38657 6783
rect 38761 6749 38795 6783
rect 38858 6749 38892 6783
rect 39037 6749 39071 6783
rect 1593 6681 1627 6715
rect 13461 6681 13495 6715
rect 19349 6681 19383 6715
rect 27261 6681 27295 6715
rect 28549 6681 28583 6715
rect 30196 6681 30230 6715
rect 33977 6681 34011 6715
rect 34161 6681 34195 6715
rect 3249 6613 3283 6647
rect 3801 6613 3835 6647
rect 6009 6613 6043 6647
rect 8125 6613 8159 6647
rect 9137 6613 9171 6647
rect 9597 6613 9631 6647
rect 12173 6613 12207 6647
rect 14197 6613 14231 6647
rect 17601 6613 17635 6647
rect 18337 6613 18371 6647
rect 19993 6613 20027 6647
rect 20729 6613 20763 6647
rect 23213 6613 23247 6647
rect 34897 6613 34931 6647
rect 37289 6613 37323 6647
rect 38393 6613 38427 6647
rect 15577 6409 15611 6443
rect 23673 6409 23707 6443
rect 27629 6409 27663 6443
rect 30205 6409 30239 6443
rect 37289 6409 37323 6443
rect 39681 6409 39715 6443
rect 3249 6341 3283 6375
rect 4997 6341 5031 6375
rect 9864 6341 9898 6375
rect 19073 6341 19107 6375
rect 19533 6341 19567 6375
rect 23305 6341 23339 6375
rect 23397 6341 23431 6375
rect 30849 6341 30883 6375
rect 34437 6341 34471 6375
rect 36277 6341 36311 6375
rect 36461 6341 36495 6375
rect 37657 6341 37691 6375
rect 38546 6341 38580 6375
rect 2513 6273 2547 6307
rect 5641 6273 5675 6307
rect 5825 6273 5859 6307
rect 6469 6273 6503 6307
rect 6929 6273 6963 6307
rect 7573 6273 7607 6307
rect 8401 6273 8435 6307
rect 9045 6273 9079 6307
rect 9597 6273 9631 6307
rect 13737 6273 13771 6307
rect 14004 6273 14038 6307
rect 15761 6273 15795 6307
rect 15945 6273 15979 6307
rect 16865 6273 16899 6307
rect 17325 6273 17359 6307
rect 19717 6273 19751 6307
rect 23121 6273 23155 6307
rect 23489 6273 23523 6307
rect 24685 6273 24719 6307
rect 26985 6273 27019 6307
rect 29561 6273 29595 6307
rect 29745 6273 29779 6307
rect 29837 6273 29871 6307
rect 29975 6273 30009 6307
rect 31033 6273 31067 6307
rect 35265 6273 35299 6307
rect 35357 6273 35391 6307
rect 35449 6273 35483 6307
rect 35633 6273 35667 6307
rect 37473 6273 37507 6307
rect 38301 6273 38335 6307
rect 21833 6205 21867 6239
rect 22109 6205 22143 6239
rect 24225 6205 24259 6239
rect 29009 6205 29043 6239
rect 36093 6205 36127 6239
rect 7113 6137 7147 6171
rect 10977 6137 11011 6171
rect 27169 6137 27203 6171
rect 58173 6137 58207 6171
rect 1869 6069 1903 6103
rect 2329 6069 2363 6103
rect 5641 6069 5675 6103
rect 7757 6069 7791 6103
rect 8217 6069 8251 6103
rect 8861 6069 8895 6103
rect 11621 6069 11655 6103
rect 12265 6069 12299 6103
rect 13093 6069 13127 6103
rect 15117 6069 15151 6103
rect 19901 6069 19935 6103
rect 20729 6069 20763 6103
rect 21189 6069 21223 6103
rect 26157 6069 26191 6103
rect 30665 6069 30699 6103
rect 34989 6069 35023 6103
rect 5733 5865 5767 5899
rect 12541 5865 12575 5899
rect 18705 5865 18739 5899
rect 20637 5865 20671 5899
rect 22661 5865 22695 5899
rect 24777 5865 24811 5899
rect 29561 5865 29595 5899
rect 32689 5865 32723 5899
rect 36185 5865 36219 5899
rect 38853 5865 38887 5899
rect 3249 5797 3283 5831
rect 7297 5797 7331 5831
rect 10149 5797 10183 5831
rect 11345 5797 11379 5831
rect 16221 5797 16255 5831
rect 4261 5729 4295 5763
rect 4445 5729 4479 5763
rect 5549 5729 5583 5763
rect 9505 5729 9539 5763
rect 17601 5729 17635 5763
rect 19257 5729 19291 5763
rect 23213 5729 23247 5763
rect 25605 5729 25639 5763
rect 1869 5661 1903 5695
rect 2136 5661 2170 5695
rect 5457 5661 5491 5695
rect 6377 5661 6411 5695
rect 8401 5661 8435 5695
rect 10793 5661 10827 5695
rect 11529 5661 11563 5695
rect 12541 5661 12575 5695
rect 12725 5661 12759 5695
rect 13369 5661 13403 5695
rect 14105 5661 14139 5695
rect 15117 5661 15151 5695
rect 15301 5661 15335 5695
rect 15393 5661 15427 5695
rect 15485 5661 15519 5695
rect 18061 5661 18095 5695
rect 18245 5661 18279 5695
rect 18337 5661 18371 5695
rect 18429 5661 18463 5695
rect 22109 5661 22143 5695
rect 22293 5661 22327 5695
rect 22477 5661 22511 5695
rect 24593 5661 24627 5695
rect 25881 5661 25915 5695
rect 30113 5661 30147 5695
rect 30297 5661 30331 5695
rect 30389 5661 30423 5695
rect 30527 5661 30561 5695
rect 31309 5661 31343 5695
rect 34805 5661 34839 5695
rect 37473 5661 37507 5695
rect 37729 5661 37763 5695
rect 4169 5593 4203 5627
rect 6561 5593 6595 5627
rect 7113 5593 7147 5627
rect 16405 5593 16439 5627
rect 16589 5593 16623 5627
rect 19502 5593 19536 5627
rect 22385 5593 22419 5627
rect 24409 5593 24443 5627
rect 30757 5593 30791 5627
rect 31554 5593 31588 5627
rect 35050 5593 35084 5627
rect 3801 5525 3835 5559
rect 5089 5525 5123 5559
rect 11989 5525 12023 5559
rect 15761 5525 15795 5559
rect 21649 5525 21683 5559
rect 23673 5525 23707 5559
rect 26985 5525 27019 5559
rect 2513 5321 2547 5355
rect 4997 5321 5031 5355
rect 5181 5321 5215 5355
rect 6561 5321 6595 5355
rect 12449 5321 12483 5355
rect 19073 5321 19107 5355
rect 23765 5321 23799 5355
rect 25605 5321 25639 5355
rect 35449 5321 35483 5355
rect 1501 5253 1535 5287
rect 19441 5253 19475 5287
rect 24900 5253 24934 5287
rect 27997 5253 28031 5287
rect 33701 5253 33735 5287
rect 34161 5253 34195 5287
rect 2697 5185 2731 5219
rect 2881 5185 2915 5219
rect 4353 5185 4387 5219
rect 5733 5217 5767 5251
rect 6377 5185 6411 5219
rect 6745 5185 6779 5219
rect 6929 5185 6963 5219
rect 7665 5185 7699 5219
rect 8309 5185 8343 5219
rect 9689 5185 9723 5219
rect 11897 5185 11931 5219
rect 12265 5185 12299 5219
rect 15025 5185 15059 5219
rect 17785 5185 17819 5219
rect 17969 5185 18003 5219
rect 18064 5185 18098 5219
rect 18173 5185 18207 5219
rect 19257 5185 19291 5219
rect 25145 5185 25179 5219
rect 28181 5185 28215 5219
rect 3893 5117 3927 5151
rect 5273 5117 5307 5151
rect 7849 5117 7883 5151
rect 11805 5117 11839 5151
rect 54401 5117 54435 5151
rect 5733 5049 5767 5083
rect 8493 5049 8527 5083
rect 10977 5049 11011 5083
rect 13093 5049 13127 5083
rect 18429 5049 18463 5083
rect 55045 5049 55079 5083
rect 2053 4981 2087 5015
rect 4537 4981 4571 5015
rect 6745 4981 6779 5015
rect 7481 4981 7515 5015
rect 10333 4981 10367 5015
rect 12265 4981 12299 5015
rect 13737 4981 13771 5015
rect 14197 4981 14231 5015
rect 14841 4981 14875 5015
rect 15761 4981 15795 5015
rect 17325 4981 17359 5015
rect 20177 4981 20211 5015
rect 21005 4981 21039 5015
rect 21833 4981 21867 5015
rect 22661 4981 22695 5015
rect 27813 4981 27847 5015
rect 53757 4981 53791 5015
rect 58173 4981 58207 5015
rect 3249 4777 3283 4811
rect 6929 4777 6963 4811
rect 7941 4777 7975 4811
rect 8309 4777 8343 4811
rect 8953 4777 8987 4811
rect 9413 4777 9447 4811
rect 10333 4777 10367 4811
rect 11713 4777 11747 4811
rect 11897 4777 11931 4811
rect 22477 4777 22511 4811
rect 2053 4709 2087 4743
rect 6837 4709 6871 4743
rect 10517 4709 10551 4743
rect 11621 4709 11655 4743
rect 17417 4709 17451 4743
rect 26433 4709 26467 4743
rect 52837 4709 52871 4743
rect 55321 4709 55355 4743
rect 6653 4641 6687 4675
rect 9045 4641 9079 4675
rect 10425 4641 10459 4675
rect 11805 4641 11839 4675
rect 12909 4641 12943 4675
rect 16129 4641 16163 4675
rect 18061 4641 18095 4675
rect 23857 4641 23891 4675
rect 31493 4641 31527 4675
rect 54125 4641 54159 4675
rect 55965 4641 55999 4675
rect 3065 4573 3099 4607
rect 3893 4573 3927 4607
rect 4721 4573 4755 4607
rect 4905 4573 4939 4607
rect 6193 4573 6227 4607
rect 6929 4573 6963 4607
rect 7481 4573 7515 4607
rect 7573 4573 7607 4607
rect 8007 4573 8041 4607
rect 8953 4573 8987 4607
rect 9229 4573 9263 4607
rect 10646 4573 10680 4607
rect 11253 4573 11287 4607
rect 13369 4573 13403 4607
rect 14841 4573 14875 4607
rect 15485 4573 15519 4607
rect 16773 4573 16807 4607
rect 18705 4573 18739 4607
rect 19441 4573 19475 4607
rect 20085 4573 20119 4607
rect 20729 4573 20763 4607
rect 21373 4573 21407 4607
rect 22017 4573 22051 4607
rect 23590 4573 23624 4607
rect 24961 4573 24995 4607
rect 27169 4573 27203 4607
rect 27261 4573 27295 4607
rect 27353 4573 27387 4607
rect 27537 4573 27571 4607
rect 30021 4573 30055 4607
rect 30205 4573 30239 4607
rect 30297 4573 30331 4607
rect 30435 4573 30469 4607
rect 31125 4573 31159 4607
rect 31309 4573 31343 4607
rect 52193 4573 52227 4607
rect 53481 4573 53515 4607
rect 1501 4505 1535 4539
rect 10793 4505 10827 4539
rect 25513 4505 25547 4539
rect 2605 4437 2639 4471
rect 4077 4437 4111 4471
rect 4537 4437 4571 4471
rect 5457 4437 5491 4471
rect 6009 4437 6043 4471
rect 13553 4437 13587 4471
rect 14197 4437 14231 4471
rect 24409 4437 24443 4471
rect 26893 4437 26927 4471
rect 30665 4437 30699 4471
rect 6561 4233 6595 4267
rect 8769 4233 8803 4267
rect 9781 4233 9815 4267
rect 29929 4233 29963 4267
rect 4905 4165 4939 4199
rect 6377 4165 6411 4199
rect 7665 4165 7699 4199
rect 2329 4097 2363 4131
rect 2789 4097 2823 4131
rect 3433 4097 3467 4131
rect 4077 4097 4111 4131
rect 5825 4097 5859 4131
rect 8125 4097 8159 4131
rect 8953 4097 8987 4131
rect 9137 4097 9171 4131
rect 9597 4097 9631 4131
rect 10609 4097 10643 4131
rect 11529 4097 11563 4131
rect 16681 4097 16715 4131
rect 16948 4097 16982 4131
rect 19441 4097 19475 4131
rect 19697 4097 19731 4131
rect 34897 4097 34931 4131
rect 35164 4097 35198 4131
rect 54677 4097 54711 4131
rect 7941 4029 7975 4063
rect 12081 4029 12115 4063
rect 12357 4029 12391 4063
rect 14841 4029 14875 4063
rect 52745 4029 52779 4063
rect 55965 4029 55999 4063
rect 2973 3961 3007 3995
rect 10425 3961 10459 3995
rect 11989 3961 12023 3995
rect 14197 3961 14231 3995
rect 15485 3961 15519 3995
rect 20821 3961 20855 3995
rect 26065 3961 26099 3995
rect 1685 3893 1719 3927
rect 2145 3893 2179 3927
rect 3617 3893 3651 3927
rect 4261 3893 4295 3927
rect 4997 3893 5031 3927
rect 5641 3893 5675 3927
rect 6561 3893 6595 3927
rect 6745 3893 6779 3927
rect 7757 3893 7791 3927
rect 8309 3893 8343 3927
rect 8953 3893 8987 3927
rect 11897 3893 11931 3927
rect 13553 3893 13587 3927
rect 16129 3893 16163 3927
rect 18061 3893 18095 3927
rect 18981 3893 19015 3927
rect 22385 3893 22419 3927
rect 23029 3893 23063 3927
rect 23489 3893 23523 3927
rect 24317 3893 24351 3927
rect 25421 3893 25455 3927
rect 36277 3893 36311 3927
rect 51181 3893 51215 3927
rect 51825 3893 51859 3927
rect 53389 3893 53423 3927
rect 54033 3893 54067 3927
rect 55321 3893 55355 3927
rect 58173 3893 58207 3927
rect 3249 3689 3283 3723
rect 5917 3689 5951 3723
rect 6101 3689 6135 3723
rect 8309 3689 8343 3723
rect 9413 3689 9447 3723
rect 10517 3689 10551 3723
rect 12265 3689 12299 3723
rect 16129 3689 16163 3723
rect 17049 3689 17083 3723
rect 17785 3689 17819 3723
rect 18613 3689 18647 3723
rect 21005 3689 21039 3723
rect 27997 3689 28031 3723
rect 32413 3689 32447 3723
rect 3893 3621 3927 3655
rect 8953 3621 8987 3655
rect 9321 3621 9355 3655
rect 13553 3621 13587 3655
rect 14841 3621 14875 3655
rect 20361 3621 20395 3655
rect 21741 3621 21775 3655
rect 46949 3621 46983 3655
rect 52837 3621 52871 3655
rect 55321 3621 55355 3655
rect 5273 3553 5307 3587
rect 6561 3553 6595 3587
rect 6837 3553 6871 3587
rect 9505 3553 9539 3587
rect 9873 3553 9907 3587
rect 14381 3553 14415 3587
rect 19625 3553 19659 3587
rect 26617 3553 26651 3587
rect 31033 3553 31067 3587
rect 51549 3553 51583 3587
rect 53481 3553 53515 3587
rect 56609 3553 56643 3587
rect 1869 3485 1903 3519
rect 8033 3485 8067 3519
rect 10333 3485 10367 3519
rect 11069 3485 11103 3519
rect 12725 3485 12759 3519
rect 13369 3485 13403 3519
rect 15945 3485 15979 3519
rect 16865 3485 16899 3519
rect 17601 3485 17635 3519
rect 18521 3485 18555 3519
rect 21097 3485 21131 3519
rect 21925 3485 21959 3519
rect 23213 3485 23247 3519
rect 23857 3485 23891 3519
rect 24685 3485 24719 3519
rect 25513 3485 25547 3519
rect 26157 3485 26191 3519
rect 26884 3485 26918 3519
rect 28733 3485 28767 3519
rect 31289 3485 31323 3519
rect 34805 3485 34839 3519
rect 35449 3485 35483 3519
rect 36093 3485 36127 3519
rect 36737 3485 36771 3519
rect 37565 3485 37599 3519
rect 38669 3485 38703 3519
rect 40049 3485 40083 3519
rect 40693 3485 40727 3519
rect 41337 3485 41371 3519
rect 42533 3485 42567 3519
rect 43177 3485 43211 3519
rect 45017 3485 45051 3519
rect 45661 3485 45695 3519
rect 46305 3485 46339 3519
rect 47777 3485 47811 3519
rect 48421 3485 48455 3519
rect 50261 3485 50295 3519
rect 50905 3485 50939 3519
rect 52193 3485 52227 3519
rect 54125 3485 54159 3519
rect 55965 3485 55999 3519
rect 57529 3485 57563 3519
rect 58173 3485 58207 3519
rect 2136 3417 2170 3451
rect 5028 3417 5062 3451
rect 5733 3417 5767 3451
rect 14289 3417 14323 3451
rect 14841 3417 14875 3451
rect 15485 3417 15519 3451
rect 20177 3417 20211 3451
rect 5933 3349 5967 3383
rect 11253 3349 11287 3383
rect 12909 3349 12943 3383
rect 14105 3349 14139 3383
rect 22569 3349 22603 3383
rect 3801 3145 3835 3179
rect 8953 3145 8987 3179
rect 11621 3145 11655 3179
rect 14565 3145 14599 3179
rect 15301 3145 15335 3179
rect 15945 3145 15979 3179
rect 17417 3145 17451 3179
rect 18153 3145 18187 3179
rect 19625 3145 19659 3179
rect 20361 3145 20395 3179
rect 22293 3145 22327 3179
rect 23029 3145 23063 3179
rect 2688 3077 2722 3111
rect 18245 3077 18279 3111
rect 18797 3077 18831 3111
rect 18981 3077 19015 3111
rect 20453 3077 20487 3111
rect 21005 3077 21039 3111
rect 21189 3077 21223 3111
rect 22201 3077 22235 3111
rect 1777 3009 1811 3043
rect 2421 3009 2455 3043
rect 5089 3009 5123 3043
rect 5825 3009 5859 3043
rect 8125 3009 8159 3043
rect 9597 3009 9631 3043
rect 9965 3009 9999 3043
rect 10517 3009 10551 3043
rect 10885 3009 10919 3043
rect 11805 3009 11839 3043
rect 12265 3009 12299 3043
rect 14381 3009 14415 3043
rect 15117 3009 15151 3043
rect 16129 3009 16163 3043
rect 17601 3009 17635 3043
rect 19809 3009 19843 3043
rect 22845 3009 22879 3043
rect 54033 3009 54067 3043
rect 54677 3009 54711 3043
rect 55321 3009 55355 3043
rect 6837 2941 6871 2975
rect 7113 2941 7147 2975
rect 8677 2941 8711 2975
rect 13921 2941 13955 2975
rect 23857 2941 23891 2975
rect 25789 2941 25823 2975
rect 33425 2941 33459 2975
rect 39221 2941 39255 2975
rect 43085 2941 43119 2975
rect 55965 2941 55999 2975
rect 56609 2941 56643 2975
rect 4353 2873 4387 2907
rect 8585 2873 8619 2907
rect 13277 2873 13311 2907
rect 16865 2873 16899 2907
rect 34069 2873 34103 2907
rect 35357 2873 35391 2907
rect 37933 2873 37967 2907
rect 39865 2873 39899 2907
rect 41153 2873 41187 2907
rect 43729 2873 43763 2907
rect 45017 2873 45051 2907
rect 45661 2873 45695 2907
rect 48237 2873 48271 2907
rect 49525 2873 49559 2907
rect 50813 2873 50847 2907
rect 52745 2873 52779 2907
rect 57897 2873 57931 2907
rect 1961 2805 1995 2839
rect 4905 2805 4939 2839
rect 5641 2805 5675 2839
rect 8493 2805 8527 2839
rect 12449 2805 12483 2839
rect 24501 2805 24535 2839
rect 25145 2805 25179 2839
rect 26433 2805 26467 2839
rect 27629 2805 27663 2839
rect 28089 2805 28123 2839
rect 28917 2805 28951 2839
rect 29561 2805 29595 2839
rect 30021 2805 30055 2839
rect 30665 2805 30699 2839
rect 32137 2805 32171 2839
rect 32781 2805 32815 2839
rect 34713 2805 34747 2839
rect 36001 2805 36035 2839
rect 37289 2805 37323 2839
rect 38577 2805 38611 2839
rect 40509 2805 40543 2839
rect 42441 2805 42475 2839
rect 44373 2805 44407 2839
rect 46305 2805 46339 2839
rect 47593 2805 47627 2839
rect 48881 2805 48915 2839
rect 50169 2805 50203 2839
rect 51457 2805 51491 2839
rect 53389 2805 53423 2839
rect 10425 2601 10459 2635
rect 12449 2601 12483 2635
rect 13461 2601 13495 2635
rect 14565 2601 14599 2635
rect 17417 2601 17451 2635
rect 55321 2601 55355 2635
rect 2329 2533 2363 2567
rect 3065 2533 3099 2567
rect 11713 2533 11747 2567
rect 15209 2533 15243 2567
rect 16129 2533 16163 2567
rect 18061 2533 18095 2567
rect 19257 2533 19291 2567
rect 20269 2533 20303 2567
rect 21097 2533 21131 2567
rect 22753 2533 22787 2567
rect 23581 2533 23615 2567
rect 25789 2533 25823 2567
rect 27721 2533 27755 2567
rect 36001 2533 36035 2567
rect 39865 2533 39899 2567
rect 43729 2533 43763 2567
rect 47593 2533 47627 2567
rect 51457 2533 51491 2567
rect 54033 2533 54067 2567
rect 5549 2465 5583 2499
rect 7849 2465 7883 2499
rect 9597 2465 9631 2499
rect 32781 2465 32815 2499
rect 34713 2465 34747 2499
rect 37289 2465 37323 2499
rect 40509 2465 40543 2499
rect 42441 2465 42475 2499
rect 45017 2465 45051 2499
rect 48237 2465 48271 2499
rect 50169 2465 50203 2499
rect 52745 2465 52779 2499
rect 57897 2465 57931 2499
rect 1593 2397 1627 2431
rect 2513 2397 2547 2431
rect 3249 2397 3283 2431
rect 4261 2397 4295 2431
rect 5825 2397 5859 2431
rect 6745 2397 6779 2431
rect 8125 2397 8159 2431
rect 11529 2397 11563 2431
rect 12265 2397 12299 2431
rect 13277 2397 13311 2431
rect 14381 2397 14415 2431
rect 15393 2397 15427 2431
rect 15945 2397 15979 2431
rect 16865 2397 16899 2431
rect 18245 2397 18279 2431
rect 21281 2397 21315 2431
rect 22201 2397 22235 2431
rect 22937 2397 22971 2431
rect 23397 2397 23431 2431
rect 24409 2397 24443 2431
rect 25145 2397 25179 2431
rect 26433 2397 26467 2431
rect 28365 2397 28399 2431
rect 29009 2397 29043 2431
rect 30113 2397 30147 2431
rect 30757 2397 30791 2431
rect 31217 2397 31251 2431
rect 32137 2397 32171 2431
rect 33425 2397 33459 2431
rect 35357 2397 35391 2431
rect 37933 2397 37967 2431
rect 38577 2397 38611 2431
rect 41153 2397 41187 2431
rect 43085 2397 43119 2431
rect 45661 2397 45695 2431
rect 46305 2397 46339 2431
rect 48881 2397 48915 2431
rect 50813 2397 50847 2431
rect 53389 2397 53423 2431
rect 55965 2397 55999 2431
rect 56609 2397 56643 2431
rect 10149 2329 10183 2363
rect 17509 2329 17543 2363
rect 19441 2329 19475 2363
rect 20453 2329 20487 2363
rect 1777 2261 1811 2295
rect 4445 2261 4479 2295
rect 6653 2261 6687 2295
rect 22017 2261 22051 2295
rect 26985 2261 27019 2295
<< metal1 >>
rect 5258 57740 5264 57792
rect 5316 57780 5322 57792
rect 18322 57780 18328 57792
rect 5316 57752 18328 57780
rect 5316 57740 5322 57752
rect 18322 57740 18328 57752
rect 18380 57740 18386 57792
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 1762 57536 1768 57588
rect 1820 57576 1826 57588
rect 1949 57579 2007 57585
rect 1949 57576 1961 57579
rect 1820 57548 1961 57576
rect 1820 57536 1826 57548
rect 1949 57545 1961 57548
rect 1995 57545 2007 57579
rect 1949 57539 2007 57545
rect 3326 57536 3332 57588
rect 3384 57576 3390 57588
rect 3881 57579 3939 57585
rect 3881 57576 3893 57579
rect 3384 57548 3893 57576
rect 3384 57536 3390 57548
rect 3881 57545 3893 57548
rect 3927 57545 3939 57579
rect 3881 57539 3939 57545
rect 4890 57536 4896 57588
rect 4948 57576 4954 57588
rect 5077 57579 5135 57585
rect 5077 57576 5089 57579
rect 4948 57548 5089 57576
rect 4948 57536 4954 57548
rect 5077 57545 5089 57548
rect 5123 57545 5135 57579
rect 5077 57539 5135 57545
rect 6454 57536 6460 57588
rect 6512 57576 6518 57588
rect 6641 57579 6699 57585
rect 6641 57576 6653 57579
rect 6512 57548 6653 57576
rect 6512 57536 6518 57548
rect 6641 57545 6653 57548
rect 6687 57545 6699 57579
rect 6641 57539 6699 57545
rect 8018 57536 8024 57588
rect 8076 57576 8082 57588
rect 8205 57579 8263 57585
rect 8205 57576 8217 57579
rect 8076 57548 8217 57576
rect 8076 57536 8082 57548
rect 8205 57545 8217 57548
rect 8251 57545 8263 57579
rect 8205 57539 8263 57545
rect 9674 57536 9680 57588
rect 9732 57576 9738 57588
rect 9769 57579 9827 57585
rect 9769 57576 9781 57579
rect 9732 57548 9781 57576
rect 9732 57536 9738 57548
rect 9769 57545 9781 57548
rect 9815 57545 9827 57579
rect 9769 57539 9827 57545
rect 11146 57536 11152 57588
rect 11204 57576 11210 57588
rect 11609 57579 11667 57585
rect 11609 57576 11621 57579
rect 11204 57548 11621 57576
rect 11204 57536 11210 57548
rect 11609 57545 11621 57548
rect 11655 57545 11667 57579
rect 11609 57539 11667 57545
rect 12710 57536 12716 57588
rect 12768 57576 12774 57588
rect 12897 57579 12955 57585
rect 12897 57576 12909 57579
rect 12768 57548 12909 57576
rect 12768 57536 12774 57548
rect 12897 57545 12909 57548
rect 12943 57545 12955 57579
rect 12897 57539 12955 57545
rect 14274 57536 14280 57588
rect 14332 57576 14338 57588
rect 14461 57579 14519 57585
rect 14461 57576 14473 57579
rect 14332 57548 14473 57576
rect 14332 57536 14338 57548
rect 14461 57545 14473 57548
rect 14507 57545 14519 57579
rect 14461 57539 14519 57545
rect 15838 57536 15844 57588
rect 15896 57576 15902 57588
rect 16761 57579 16819 57585
rect 16761 57576 16773 57579
rect 15896 57548 16773 57576
rect 15896 57536 15902 57548
rect 16761 57545 16773 57548
rect 16807 57545 16819 57579
rect 16761 57539 16819 57545
rect 17402 57536 17408 57588
rect 17460 57576 17466 57588
rect 17681 57579 17739 57585
rect 17681 57576 17693 57579
rect 17460 57548 17693 57576
rect 17460 57536 17466 57548
rect 17681 57545 17693 57548
rect 17727 57545 17739 57579
rect 17681 57539 17739 57545
rect 19334 57536 19340 57588
rect 19392 57576 19398 57588
rect 19429 57579 19487 57585
rect 19429 57576 19441 57579
rect 19392 57548 19441 57576
rect 19392 57536 19398 57548
rect 19429 57545 19441 57548
rect 19475 57545 19487 57579
rect 19429 57539 19487 57545
rect 20714 57536 20720 57588
rect 20772 57576 20778 57588
rect 20809 57579 20867 57585
rect 20809 57576 20821 57579
rect 20772 57548 20821 57576
rect 20772 57536 20778 57548
rect 20809 57545 20821 57548
rect 20855 57545 20867 57579
rect 20809 57539 20867 57545
rect 22094 57536 22100 57588
rect 22152 57576 22158 57588
rect 22373 57579 22431 57585
rect 22373 57576 22385 57579
rect 22152 57548 22385 57576
rect 22152 57536 22158 57548
rect 22373 57545 22385 57548
rect 22419 57545 22431 57579
rect 22373 57539 22431 57545
rect 23658 57536 23664 57588
rect 23716 57576 23722 57588
rect 24581 57579 24639 57585
rect 24581 57576 24593 57579
rect 23716 57548 24593 57576
rect 23716 57536 23722 57548
rect 24581 57545 24593 57548
rect 24627 57545 24639 57579
rect 24581 57539 24639 57545
rect 25222 57536 25228 57588
rect 25280 57576 25286 57588
rect 25501 57579 25559 57585
rect 25501 57576 25513 57579
rect 25280 57548 25513 57576
rect 25280 57536 25286 57548
rect 25501 57545 25513 57548
rect 25547 57545 25559 57579
rect 25501 57539 25559 57545
rect 26786 57536 26792 57588
rect 26844 57576 26850 57588
rect 27157 57579 27215 57585
rect 27157 57576 27169 57579
rect 26844 57548 27169 57576
rect 26844 57536 26850 57548
rect 27157 57545 27169 57548
rect 27203 57545 27215 57579
rect 27157 57539 27215 57545
rect 28350 57536 28356 57588
rect 28408 57576 28414 57588
rect 28629 57579 28687 57585
rect 28629 57576 28641 57579
rect 28408 57548 28641 57576
rect 28408 57536 28414 57548
rect 28629 57545 28641 57548
rect 28675 57545 28687 57579
rect 28629 57539 28687 57545
rect 29914 57536 29920 57588
rect 29972 57576 29978 57588
rect 30193 57579 30251 57585
rect 30193 57576 30205 57579
rect 29972 57548 30205 57576
rect 29972 57536 29978 57548
rect 30193 57545 30205 57548
rect 30239 57545 30251 57579
rect 30193 57539 30251 57545
rect 31478 57536 31484 57588
rect 31536 57576 31542 57588
rect 32309 57579 32367 57585
rect 32309 57576 32321 57579
rect 31536 57548 32321 57576
rect 31536 57536 31542 57548
rect 32309 57545 32321 57548
rect 32355 57545 32367 57579
rect 32309 57539 32367 57545
rect 33134 57536 33140 57588
rect 33192 57576 33198 57588
rect 33321 57579 33379 57585
rect 33321 57576 33333 57579
rect 33192 57548 33333 57576
rect 33192 57536 33198 57548
rect 33321 57545 33333 57548
rect 33367 57545 33379 57579
rect 33321 57539 33379 57545
rect 34606 57536 34612 57588
rect 34664 57576 34670 57588
rect 34885 57579 34943 57585
rect 34885 57576 34897 57579
rect 34664 57548 34897 57576
rect 34664 57536 34670 57548
rect 34885 57545 34897 57548
rect 34931 57545 34943 57579
rect 34885 57539 34943 57545
rect 36170 57536 36176 57588
rect 36228 57576 36234 57588
rect 36449 57579 36507 57585
rect 36449 57576 36461 57579
rect 36228 57548 36461 57576
rect 36228 57536 36234 57548
rect 36449 57545 36461 57548
rect 36495 57545 36507 57579
rect 36449 57539 36507 57545
rect 37734 57536 37740 57588
rect 37792 57576 37798 57588
rect 38013 57579 38071 57585
rect 38013 57576 38025 57579
rect 37792 57548 38025 57576
rect 37792 57536 37798 57548
rect 38013 57545 38025 57548
rect 38059 57545 38071 57579
rect 38013 57539 38071 57545
rect 39298 57536 39304 57588
rect 39356 57576 39362 57588
rect 40037 57579 40095 57585
rect 40037 57576 40049 57579
rect 39356 57548 40049 57576
rect 39356 57536 39362 57548
rect 40037 57545 40049 57548
rect 40083 57545 40095 57579
rect 40037 57539 40095 57545
rect 40862 57536 40868 57588
rect 40920 57576 40926 57588
rect 41141 57579 41199 57585
rect 41141 57576 41153 57579
rect 40920 57548 41153 57576
rect 40920 57536 40926 57548
rect 41141 57545 41153 57548
rect 41187 57545 41199 57579
rect 41141 57539 41199 57545
rect 42426 57536 42432 57588
rect 42484 57576 42490 57588
rect 42705 57579 42763 57585
rect 42705 57576 42717 57579
rect 42484 57548 42717 57576
rect 42484 57536 42490 57548
rect 42705 57545 42717 57548
rect 42751 57545 42763 57579
rect 42705 57539 42763 57545
rect 44174 57536 44180 57588
rect 44232 57576 44238 57588
rect 44269 57579 44327 57585
rect 44269 57576 44281 57579
rect 44232 57548 44281 57576
rect 44232 57536 44238 57548
rect 44269 57545 44281 57548
rect 44315 57545 44327 57579
rect 44269 57539 44327 57545
rect 45554 57536 45560 57588
rect 45612 57576 45618 57588
rect 45833 57579 45891 57585
rect 45833 57576 45845 57579
rect 45612 57548 45845 57576
rect 45612 57536 45618 57548
rect 45833 57545 45845 57548
rect 45879 57545 45891 57579
rect 45833 57539 45891 57545
rect 47118 57536 47124 57588
rect 47176 57576 47182 57588
rect 47765 57579 47823 57585
rect 47765 57576 47777 57579
rect 47176 57548 47777 57576
rect 47176 57536 47182 57548
rect 47765 57545 47777 57548
rect 47811 57545 47823 57579
rect 47765 57539 47823 57545
rect 19150 57508 19156 57520
rect 8404 57480 19156 57508
rect 2133 57443 2191 57449
rect 2133 57409 2145 57443
rect 2179 57440 2191 57443
rect 2682 57440 2688 57452
rect 2179 57412 2688 57440
rect 2179 57409 2191 57412
rect 2133 57403 2191 57409
rect 2682 57400 2688 57412
rect 2740 57400 2746 57452
rect 4062 57440 4068 57452
rect 4023 57412 4068 57440
rect 4062 57400 4068 57412
rect 4120 57400 4126 57452
rect 5258 57440 5264 57452
rect 5219 57412 5264 57440
rect 5258 57400 5264 57412
rect 5316 57400 5322 57452
rect 8404 57449 8432 57480
rect 19150 57468 19156 57480
rect 19208 57468 19214 57520
rect 6825 57443 6883 57449
rect 6825 57409 6837 57443
rect 6871 57409 6883 57443
rect 6825 57403 6883 57409
rect 8389 57443 8447 57449
rect 8389 57409 8401 57443
rect 8435 57409 8447 57443
rect 8389 57403 8447 57409
rect 9953 57443 10011 57449
rect 9953 57409 9965 57443
rect 9999 57409 10011 57443
rect 11790 57440 11796 57452
rect 11751 57412 11796 57440
rect 9953 57403 10011 57409
rect 6840 57372 6868 57403
rect 6840 57344 6914 57372
rect 2682 57236 2688 57248
rect 2643 57208 2688 57236
rect 2682 57196 2688 57208
rect 2740 57196 2746 57248
rect 6886 57236 6914 57344
rect 9968 57304 9996 57403
rect 11790 57400 11796 57412
rect 11848 57400 11854 57452
rect 13078 57440 13084 57452
rect 13039 57412 13084 57440
rect 13078 57400 13084 57412
rect 13136 57400 13142 57452
rect 14645 57443 14703 57449
rect 14645 57409 14657 57443
rect 14691 57440 14703 57443
rect 15930 57440 15936 57452
rect 14691 57412 15936 57440
rect 14691 57409 14703 57412
rect 14645 57403 14703 57409
rect 15930 57400 15936 57412
rect 15988 57400 15994 57452
rect 16942 57440 16948 57452
rect 16903 57412 16948 57440
rect 16942 57400 16948 57412
rect 17000 57400 17006 57452
rect 17494 57440 17500 57452
rect 17455 57412 17500 57440
rect 17494 57400 17500 57412
rect 17552 57400 17558 57452
rect 19242 57440 19248 57452
rect 19203 57412 19248 57440
rect 19242 57400 19248 57412
rect 19300 57400 19306 57452
rect 19334 57400 19340 57452
rect 19392 57440 19398 57452
rect 20625 57443 20683 57449
rect 20625 57440 20637 57443
rect 19392 57412 20637 57440
rect 19392 57400 19398 57412
rect 20625 57409 20637 57412
rect 20671 57409 20683 57443
rect 22186 57440 22192 57452
rect 22147 57412 22192 57440
rect 20625 57403 20683 57409
rect 22186 57400 22192 57412
rect 22244 57400 22250 57452
rect 24394 57440 24400 57452
rect 24355 57412 24400 57440
rect 24394 57400 24400 57412
rect 24452 57400 24458 57452
rect 25314 57440 25320 57452
rect 25275 57412 25320 57440
rect 25314 57400 25320 57412
rect 25372 57400 25378 57452
rect 26970 57440 26976 57452
rect 26931 57412 26976 57440
rect 26970 57400 26976 57412
rect 27028 57400 27034 57452
rect 28442 57440 28448 57452
rect 28403 57412 28448 57440
rect 28442 57400 28448 57412
rect 28500 57400 28506 57452
rect 30006 57440 30012 57452
rect 29967 57412 30012 57440
rect 30006 57400 30012 57412
rect 30064 57400 30070 57452
rect 32125 57443 32183 57449
rect 32125 57440 32137 57443
rect 30116 57412 32137 57440
rect 27614 57332 27620 57384
rect 27672 57372 27678 57384
rect 30116 57372 30144 57412
rect 32125 57409 32137 57412
rect 32171 57409 32183 57443
rect 32125 57403 32183 57409
rect 33137 57443 33195 57449
rect 33137 57409 33149 57443
rect 33183 57409 33195 57443
rect 33137 57403 33195 57409
rect 27672 57344 30144 57372
rect 27672 57332 27678 57344
rect 30374 57332 30380 57384
rect 30432 57372 30438 57384
rect 33152 57372 33180 57403
rect 33226 57400 33232 57452
rect 33284 57440 33290 57452
rect 34701 57443 34759 57449
rect 34701 57440 34713 57443
rect 33284 57412 34713 57440
rect 33284 57400 33290 57412
rect 34701 57409 34713 57412
rect 34747 57409 34759 57443
rect 34701 57403 34759 57409
rect 34790 57400 34796 57452
rect 34848 57440 34854 57452
rect 36265 57443 36323 57449
rect 36265 57440 36277 57443
rect 34848 57412 36277 57440
rect 34848 57400 34854 57412
rect 36265 57409 36277 57412
rect 36311 57409 36323 57443
rect 37826 57440 37832 57452
rect 37787 57412 37832 57440
rect 36265 57403 36323 57409
rect 37826 57400 37832 57412
rect 37884 57400 37890 57452
rect 37918 57400 37924 57452
rect 37976 57440 37982 57452
rect 39853 57443 39911 57449
rect 39853 57440 39865 57443
rect 37976 57412 39865 57440
rect 37976 57400 37982 57412
rect 39853 57409 39865 57412
rect 39899 57409 39911 57443
rect 40954 57440 40960 57452
rect 40915 57412 40960 57440
rect 39853 57403 39911 57409
rect 40954 57400 40960 57412
rect 41012 57400 41018 57452
rect 42334 57400 42340 57452
rect 42392 57440 42398 57452
rect 42521 57443 42579 57449
rect 42521 57440 42533 57443
rect 42392 57412 42533 57440
rect 42392 57400 42398 57412
rect 42521 57409 42533 57412
rect 42567 57409 42579 57443
rect 44082 57440 44088 57452
rect 44043 57412 44088 57440
rect 42521 57403 42579 57409
rect 44082 57400 44088 57412
rect 44140 57400 44146 57452
rect 45646 57440 45652 57452
rect 45607 57412 45652 57440
rect 45646 57400 45652 57412
rect 45704 57400 45710 57452
rect 47578 57440 47584 57452
rect 47539 57412 47584 57440
rect 47578 57400 47584 57412
rect 47636 57400 47642 57452
rect 48682 57400 48688 57452
rect 48740 57440 48746 57452
rect 48777 57443 48835 57449
rect 48777 57440 48789 57443
rect 48740 57412 48789 57440
rect 48740 57400 48746 57412
rect 48777 57409 48789 57412
rect 48823 57409 48835 57443
rect 48777 57403 48835 57409
rect 50154 57400 50160 57452
rect 50212 57440 50218 57452
rect 50341 57443 50399 57449
rect 50341 57440 50353 57443
rect 50212 57412 50353 57440
rect 50212 57400 50218 57412
rect 50341 57409 50353 57412
rect 50387 57409 50399 57443
rect 50341 57403 50399 57409
rect 51810 57400 51816 57452
rect 51868 57440 51874 57452
rect 51905 57443 51963 57449
rect 51905 57440 51917 57443
rect 51868 57412 51917 57440
rect 51868 57400 51874 57412
rect 51905 57409 51917 57412
rect 51951 57409 51963 57443
rect 51905 57403 51963 57409
rect 53374 57400 53380 57452
rect 53432 57440 53438 57452
rect 53469 57443 53527 57449
rect 53469 57440 53481 57443
rect 53432 57412 53481 57440
rect 53432 57400 53438 57412
rect 53469 57409 53481 57412
rect 53515 57409 53527 57443
rect 56594 57440 56600 57452
rect 56555 57412 56600 57440
rect 53469 57403 53527 57409
rect 56594 57400 56600 57412
rect 56652 57400 56658 57452
rect 57977 57443 58035 57449
rect 57977 57409 57989 57443
rect 58023 57440 58035 57443
rect 58066 57440 58072 57452
rect 58023 57412 58072 57440
rect 58023 57409 58035 57412
rect 57977 57403 58035 57409
rect 58066 57400 58072 57412
rect 58124 57400 58130 57452
rect 30432 57344 33180 57372
rect 30432 57332 30438 57344
rect 54938 57332 54944 57384
rect 54996 57372 55002 57384
rect 55309 57375 55367 57381
rect 55309 57372 55321 57375
rect 54996 57344 55321 57372
rect 54996 57332 55002 57344
rect 55309 57341 55321 57344
rect 55355 57341 55367 57375
rect 55309 57335 55367 57341
rect 18414 57304 18420 57316
rect 9968 57276 18420 57304
rect 18414 57264 18420 57276
rect 18472 57264 18478 57316
rect 17862 57236 17868 57248
rect 6886 57208 17868 57236
rect 17862 57196 17868 57208
rect 17920 57196 17926 57248
rect 18506 57196 18512 57248
rect 18564 57236 18570 57248
rect 18601 57239 18659 57245
rect 18601 57236 18613 57239
rect 18564 57208 18613 57236
rect 18564 57196 18570 57208
rect 18601 57205 18613 57208
rect 18647 57205 18659 57239
rect 20070 57236 20076 57248
rect 20031 57208 20076 57236
rect 18601 57199 18659 57205
rect 20070 57196 20076 57208
rect 20128 57196 20134 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 18322 57032 18328 57044
rect 18283 57004 18328 57032
rect 18322 56992 18328 57004
rect 18380 56992 18386 57044
rect 19150 56992 19156 57044
rect 19208 57032 19214 57044
rect 19245 57035 19303 57041
rect 19245 57032 19257 57035
rect 19208 57004 19257 57032
rect 19208 56992 19214 57004
rect 19245 57001 19257 57004
rect 19291 57001 19303 57035
rect 57514 57032 57520 57044
rect 57475 57004 57520 57032
rect 19245 56995 19303 57001
rect 57514 56992 57520 57004
rect 57572 56992 57578 57044
rect 11790 56924 11796 56976
rect 11848 56964 11854 56976
rect 19426 56964 19432 56976
rect 11848 56936 19432 56964
rect 11848 56924 11854 56936
rect 19426 56924 19432 56936
rect 19484 56924 19490 56976
rect 18506 56828 18512 56840
rect 18467 56800 18512 56828
rect 18506 56788 18512 56800
rect 18564 56788 18570 56840
rect 19429 56831 19487 56837
rect 19429 56797 19441 56831
rect 19475 56828 19487 56831
rect 20070 56828 20076 56840
rect 19475 56800 20076 56828
rect 19475 56797 19487 56800
rect 19429 56791 19487 56797
rect 20070 56788 20076 56800
rect 20128 56788 20134 56840
rect 25869 56831 25927 56837
rect 25869 56828 25881 56831
rect 25332 56800 25881 56828
rect 17865 56695 17923 56701
rect 17865 56661 17877 56695
rect 17911 56692 17923 56695
rect 18046 56692 18052 56704
rect 17911 56664 18052 56692
rect 17911 56661 17923 56664
rect 17865 56655 17923 56661
rect 18046 56652 18052 56664
rect 18104 56652 18110 56704
rect 19978 56652 19984 56704
rect 20036 56692 20042 56704
rect 20073 56695 20131 56701
rect 20073 56692 20085 56695
rect 20036 56664 20085 56692
rect 20036 56652 20042 56664
rect 20073 56661 20085 56664
rect 20119 56661 20131 56695
rect 20714 56692 20720 56704
rect 20675 56664 20720 56692
rect 20073 56655 20131 56661
rect 20714 56652 20720 56664
rect 20772 56652 20778 56704
rect 22278 56692 22284 56704
rect 22239 56664 22284 56692
rect 22278 56652 22284 56664
rect 22336 56652 22342 56704
rect 25130 56652 25136 56704
rect 25188 56692 25194 56704
rect 25332 56701 25360 56800
rect 25869 56797 25881 56800
rect 25915 56797 25927 56831
rect 25869 56791 25927 56797
rect 57882 56788 57888 56840
rect 57940 56828 57946 56840
rect 58161 56831 58219 56837
rect 58161 56828 58173 56831
rect 57940 56800 58173 56828
rect 57940 56788 57946 56800
rect 58161 56797 58173 56800
rect 58207 56797 58219 56831
rect 58161 56791 58219 56797
rect 30006 56760 30012 56772
rect 26206 56732 30012 56760
rect 25317 56695 25375 56701
rect 25317 56692 25329 56695
rect 25188 56664 25329 56692
rect 25188 56652 25194 56664
rect 25317 56661 25329 56664
rect 25363 56661 25375 56695
rect 25317 56655 25375 56661
rect 26053 56695 26111 56701
rect 26053 56661 26065 56695
rect 26099 56692 26111 56695
rect 26206 56692 26234 56732
rect 30006 56720 30012 56732
rect 30064 56720 30070 56772
rect 26602 56692 26608 56704
rect 26099 56664 26234 56692
rect 26563 56664 26608 56692
rect 26099 56661 26111 56664
rect 26053 56655 26111 56661
rect 26602 56652 26608 56664
rect 26660 56652 26666 56704
rect 42334 56692 42340 56704
rect 42295 56664 42340 56692
rect 42334 56652 42340 56664
rect 42392 56652 42398 56704
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 13078 56448 13084 56500
rect 13136 56488 13142 56500
rect 13541 56491 13599 56497
rect 13541 56488 13553 56491
rect 13136 56460 13553 56488
rect 13136 56448 13142 56460
rect 13541 56457 13553 56460
rect 13587 56457 13599 56491
rect 15930 56488 15936 56500
rect 15891 56460 15936 56488
rect 13541 56451 13599 56457
rect 15930 56448 15936 56460
rect 15988 56448 15994 56500
rect 17405 56491 17463 56497
rect 17405 56457 17417 56491
rect 17451 56488 17463 56491
rect 17494 56488 17500 56500
rect 17451 56460 17500 56488
rect 17451 56457 17463 56460
rect 17405 56451 17463 56457
rect 17494 56448 17500 56460
rect 17552 56448 17558 56500
rect 17862 56488 17868 56500
rect 17823 56460 17868 56488
rect 17862 56448 17868 56460
rect 17920 56448 17926 56500
rect 18414 56448 18420 56500
rect 18472 56488 18478 56500
rect 18509 56491 18567 56497
rect 18509 56488 18521 56491
rect 18472 56460 18521 56488
rect 18472 56448 18478 56460
rect 18509 56457 18521 56460
rect 18555 56457 18567 56491
rect 19334 56488 19340 56500
rect 19295 56460 19340 56488
rect 18509 56451 18567 56457
rect 19334 56448 19340 56460
rect 19392 56448 19398 56500
rect 19797 56491 19855 56497
rect 19797 56457 19809 56491
rect 19843 56457 19855 56491
rect 19797 56451 19855 56457
rect 21269 56491 21327 56497
rect 21269 56457 21281 56491
rect 21315 56488 21327 56491
rect 22186 56488 22192 56500
rect 21315 56460 22192 56488
rect 21315 56457 21327 56460
rect 21269 56451 21327 56457
rect 18874 56420 18880 56432
rect 18248 56392 18880 56420
rect 13722 56352 13728 56364
rect 13683 56324 13728 56352
rect 13722 56312 13728 56324
rect 13780 56312 13786 56364
rect 16117 56355 16175 56361
rect 16117 56321 16129 56355
rect 16163 56352 16175 56355
rect 16206 56352 16212 56364
rect 16163 56324 16212 56352
rect 16163 56321 16175 56324
rect 16117 56315 16175 56321
rect 16206 56312 16212 56324
rect 16264 56312 16270 56364
rect 16761 56355 16819 56361
rect 16761 56321 16773 56355
rect 16807 56352 16819 56355
rect 17221 56355 17279 56361
rect 17221 56352 17233 56355
rect 16807 56324 17233 56352
rect 16807 56321 16819 56324
rect 16761 56315 16819 56321
rect 17221 56321 17233 56324
rect 17267 56352 17279 56355
rect 17402 56352 17408 56364
rect 17267 56324 17408 56352
rect 17267 56321 17279 56324
rect 17221 56315 17279 56321
rect 17402 56312 17408 56324
rect 17460 56312 17466 56364
rect 18046 56352 18052 56364
rect 17959 56324 18052 56352
rect 18046 56312 18052 56324
rect 18104 56352 18110 56364
rect 18248 56352 18276 56392
rect 18874 56380 18880 56392
rect 18932 56380 18938 56432
rect 18690 56352 18696 56364
rect 18104 56324 18276 56352
rect 18651 56324 18696 56352
rect 18104 56312 18110 56324
rect 18690 56312 18696 56324
rect 18748 56312 18754 56364
rect 18966 56312 18972 56364
rect 19024 56352 19030 56364
rect 19153 56355 19211 56361
rect 19153 56352 19165 56355
rect 19024 56324 19165 56352
rect 19024 56312 19030 56324
rect 19153 56321 19165 56324
rect 19199 56321 19211 56355
rect 19153 56315 19211 56321
rect 2682 56244 2688 56296
rect 2740 56284 2746 56296
rect 19812 56284 19840 56451
rect 22186 56448 22192 56460
rect 22244 56448 22250 56500
rect 22833 56491 22891 56497
rect 22833 56457 22845 56491
rect 22879 56488 22891 56491
rect 24394 56488 24400 56500
rect 22879 56460 24400 56488
rect 22879 56457 22891 56460
rect 22833 56451 22891 56457
rect 24394 56448 24400 56460
rect 24452 56448 24458 56500
rect 26421 56491 26479 56497
rect 26421 56457 26433 56491
rect 26467 56488 26479 56491
rect 26970 56488 26976 56500
rect 26467 56460 26976 56488
rect 26467 56457 26479 56460
rect 26421 56451 26479 56457
rect 26970 56448 26976 56460
rect 27028 56448 27034 56500
rect 27341 56491 27399 56497
rect 27341 56457 27353 56491
rect 27387 56488 27399 56491
rect 27614 56488 27620 56500
rect 27387 56460 27620 56488
rect 27387 56457 27399 56460
rect 27341 56451 27399 56457
rect 27614 56448 27620 56460
rect 27672 56448 27678 56500
rect 29825 56491 29883 56497
rect 29825 56457 29837 56491
rect 29871 56488 29883 56491
rect 30374 56488 30380 56500
rect 29871 56460 30380 56488
rect 29871 56457 29883 56460
rect 29825 56451 29883 56457
rect 30374 56448 30380 56460
rect 30432 56448 30438 56500
rect 32309 56491 32367 56497
rect 32309 56457 32321 56491
rect 32355 56488 32367 56491
rect 33226 56488 33232 56500
rect 32355 56460 33232 56488
rect 32355 56457 32367 56460
rect 32309 56451 32367 56457
rect 33226 56448 33232 56460
rect 33284 56448 33290 56500
rect 34149 56491 34207 56497
rect 34149 56457 34161 56491
rect 34195 56488 34207 56491
rect 34790 56488 34796 56500
rect 34195 56460 34796 56488
rect 34195 56457 34207 56460
rect 34149 56451 34207 56457
rect 34790 56448 34796 56460
rect 34848 56448 34854 56500
rect 35989 56491 36047 56497
rect 35989 56457 36001 56491
rect 36035 56488 36047 56491
rect 37918 56488 37924 56500
rect 36035 56460 37924 56488
rect 36035 56457 36047 56460
rect 35989 56451 36047 56457
rect 37918 56448 37924 56460
rect 37976 56448 37982 56500
rect 45097 56491 45155 56497
rect 45097 56457 45109 56491
rect 45143 56488 45155 56491
rect 45646 56488 45652 56500
rect 45143 56460 45652 56488
rect 45143 56457 45155 56460
rect 45097 56451 45155 56457
rect 45646 56448 45652 56460
rect 45704 56448 45710 56500
rect 45741 56491 45799 56497
rect 45741 56457 45753 56491
rect 45787 56488 45799 56491
rect 47578 56488 47584 56500
rect 45787 56460 47584 56488
rect 45787 56457 45799 56460
rect 45741 56451 45799 56457
rect 47578 56448 47584 56460
rect 47636 56448 47642 56500
rect 42334 56420 42340 56432
rect 30852 56392 42340 56420
rect 19978 56352 19984 56364
rect 19939 56324 19984 56352
rect 19978 56312 19984 56324
rect 20036 56312 20042 56364
rect 20530 56312 20536 56364
rect 20588 56352 20594 56364
rect 20625 56355 20683 56361
rect 20625 56352 20637 56355
rect 20588 56324 20637 56352
rect 20588 56312 20594 56324
rect 20625 56321 20637 56324
rect 20671 56352 20683 56355
rect 20714 56352 20720 56364
rect 20671 56324 20720 56352
rect 20671 56321 20683 56324
rect 20625 56315 20683 56321
rect 20714 56312 20720 56324
rect 20772 56312 20778 56364
rect 21082 56352 21088 56364
rect 21043 56324 21088 56352
rect 21082 56312 21088 56324
rect 21140 56312 21146 56364
rect 21634 56312 21640 56364
rect 21692 56352 21698 56364
rect 22005 56355 22063 56361
rect 22005 56352 22017 56355
rect 21692 56324 22017 56352
rect 21692 56312 21698 56324
rect 22005 56321 22017 56324
rect 22051 56352 22063 56355
rect 22278 56352 22284 56364
rect 22051 56324 22284 56352
rect 22051 56321 22063 56324
rect 22005 56315 22063 56321
rect 22278 56312 22284 56324
rect 22336 56312 22342 56364
rect 22554 56312 22560 56364
rect 22612 56352 22618 56364
rect 22649 56355 22707 56361
rect 22649 56352 22661 56355
rect 22612 56324 22661 56352
rect 22612 56312 22618 56324
rect 22649 56321 22661 56324
rect 22695 56321 22707 56355
rect 22649 56315 22707 56321
rect 23477 56355 23535 56361
rect 23477 56321 23489 56355
rect 23523 56352 23535 56355
rect 23934 56352 23940 56364
rect 23523 56324 23940 56352
rect 23523 56321 23535 56324
rect 23477 56315 23535 56321
rect 23934 56312 23940 56324
rect 23992 56312 23998 56364
rect 24946 56352 24952 56364
rect 24907 56324 24952 56352
rect 24946 56312 24952 56324
rect 25004 56312 25010 56364
rect 25590 56352 25596 56364
rect 25551 56324 25596 56352
rect 25590 56312 25596 56324
rect 25648 56312 25654 56364
rect 26237 56355 26295 56361
rect 26237 56321 26249 56355
rect 26283 56352 26295 56355
rect 26602 56352 26608 56364
rect 26283 56324 26608 56352
rect 26283 56321 26295 56324
rect 26237 56315 26295 56321
rect 26602 56312 26608 56324
rect 26660 56312 26666 56364
rect 27154 56352 27160 56364
rect 27115 56324 27160 56352
rect 27154 56312 27160 56324
rect 27212 56352 27218 56364
rect 27801 56355 27859 56361
rect 27801 56352 27813 56355
rect 27212 56324 27813 56352
rect 27212 56312 27218 56324
rect 27801 56321 27813 56324
rect 27847 56321 27859 56355
rect 29638 56352 29644 56364
rect 29599 56324 29644 56352
rect 27801 56315 27859 56321
rect 29638 56312 29644 56324
rect 29696 56352 29702 56364
rect 30285 56355 30343 56361
rect 30285 56352 30297 56355
rect 29696 56324 30297 56352
rect 29696 56312 29702 56324
rect 30285 56321 30297 56324
rect 30331 56321 30343 56355
rect 30285 56315 30343 56321
rect 30852 56284 30880 56392
rect 42334 56380 42340 56392
rect 42392 56380 42398 56432
rect 30929 56355 30987 56361
rect 30929 56321 30941 56355
rect 30975 56352 30987 56355
rect 31389 56355 31447 56361
rect 31389 56352 31401 56355
rect 30975 56324 31401 56352
rect 30975 56321 30987 56324
rect 30929 56315 30987 56321
rect 31389 56321 31401 56324
rect 31435 56352 31447 56355
rect 31662 56352 31668 56364
rect 31435 56324 31668 56352
rect 31435 56321 31447 56324
rect 31389 56315 31447 56321
rect 31662 56312 31668 56324
rect 31720 56312 31726 56364
rect 32122 56352 32128 56364
rect 32083 56324 32128 56352
rect 32122 56312 32128 56324
rect 32180 56352 32186 56364
rect 32769 56355 32827 56361
rect 32769 56352 32781 56355
rect 32180 56324 32781 56352
rect 32180 56312 32186 56324
rect 32769 56321 32781 56324
rect 32815 56321 32827 56355
rect 33962 56352 33968 56364
rect 33923 56324 33968 56352
rect 32769 56315 32827 56321
rect 33962 56312 33968 56324
rect 34020 56352 34026 56364
rect 34609 56355 34667 56361
rect 34609 56352 34621 56355
rect 34020 56324 34621 56352
rect 34020 56312 34026 56324
rect 34609 56321 34621 56324
rect 34655 56321 34667 56355
rect 35802 56352 35808 56364
rect 35715 56324 35808 56352
rect 34609 56315 34667 56321
rect 35802 56312 35808 56324
rect 35860 56352 35866 56364
rect 36449 56355 36507 56361
rect 36449 56352 36461 56355
rect 35860 56324 36461 56352
rect 35860 56312 35866 56324
rect 36449 56321 36461 56324
rect 36495 56321 36507 56355
rect 44913 56355 44971 56361
rect 44913 56352 44925 56355
rect 36449 56315 36507 56321
rect 44376 56324 44925 56352
rect 2740 56256 19840 56284
rect 22204 56256 30880 56284
rect 2740 56244 2746 56256
rect 4062 56176 4068 56228
rect 4120 56216 4126 56228
rect 22204 56225 22232 56256
rect 20441 56219 20499 56225
rect 20441 56216 20453 56219
rect 4120 56188 20453 56216
rect 4120 56176 4126 56188
rect 20441 56185 20453 56188
rect 20487 56185 20499 56219
rect 20441 56179 20499 56185
rect 22189 56219 22247 56225
rect 22189 56185 22201 56219
rect 22235 56185 22247 56219
rect 22189 56179 22247 56185
rect 24121 56219 24179 56225
rect 24121 56185 24133 56219
rect 24167 56216 24179 56219
rect 25314 56216 25320 56228
rect 24167 56188 25320 56216
rect 24167 56185 24179 56188
rect 24121 56179 24179 56185
rect 25314 56176 25320 56188
rect 25372 56176 25378 56228
rect 25777 56219 25835 56225
rect 25777 56185 25789 56219
rect 25823 56216 25835 56219
rect 40954 56216 40960 56228
rect 25823 56188 40960 56216
rect 25823 56185 25835 56188
rect 25777 56179 25835 56185
rect 40954 56176 40960 56188
rect 41012 56176 41018 56228
rect 44082 56216 44088 56228
rect 41064 56188 44088 56216
rect 13722 56108 13728 56160
rect 13780 56148 13786 56160
rect 14277 56151 14335 56157
rect 14277 56148 14289 56151
rect 13780 56120 14289 56148
rect 13780 56108 13786 56120
rect 14277 56117 14289 56120
rect 14323 56148 14335 56151
rect 18782 56148 18788 56160
rect 14323 56120 18788 56148
rect 14323 56117 14335 56120
rect 14277 56111 14335 56117
rect 18782 56108 18788 56120
rect 18840 56108 18846 56160
rect 25130 56148 25136 56160
rect 25091 56120 25136 56148
rect 25130 56108 25136 56120
rect 25188 56108 25194 56160
rect 31573 56151 31631 56157
rect 31573 56117 31585 56151
rect 31619 56148 31631 56151
rect 41064 56148 41092 56188
rect 44082 56176 44088 56188
rect 44140 56176 44146 56228
rect 31619 56120 41092 56148
rect 31619 56117 31631 56120
rect 31573 56111 31631 56117
rect 42058 56108 42064 56160
rect 42116 56148 42122 56160
rect 44376 56157 44404 56324
rect 44913 56321 44925 56324
rect 44959 56321 44971 56355
rect 44913 56315 44971 56321
rect 45554 56312 45560 56364
rect 45612 56352 45618 56364
rect 46201 56355 46259 56361
rect 46201 56352 46213 56355
rect 45612 56324 46213 56352
rect 45612 56312 45618 56324
rect 46201 56321 46213 56324
rect 46247 56321 46259 56355
rect 46201 56315 46259 56321
rect 58161 56355 58219 56361
rect 58161 56321 58173 56355
rect 58207 56352 58219 56355
rect 58434 56352 58440 56364
rect 58207 56324 58440 56352
rect 58207 56321 58219 56324
rect 58161 56315 58219 56321
rect 58434 56312 58440 56324
rect 58492 56312 58498 56364
rect 44361 56151 44419 56157
rect 44361 56148 44373 56151
rect 42116 56120 44373 56148
rect 42116 56108 42122 56120
rect 44361 56117 44373 56120
rect 44407 56117 44419 56151
rect 44361 56111 44419 56117
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 16853 55947 16911 55953
rect 16853 55913 16865 55947
rect 16899 55944 16911 55947
rect 16942 55944 16948 55956
rect 16899 55916 16948 55944
rect 16899 55913 16911 55916
rect 16853 55907 16911 55913
rect 16942 55904 16948 55916
rect 17000 55904 17006 55956
rect 18693 55947 18751 55953
rect 18693 55913 18705 55947
rect 18739 55944 18751 55947
rect 19242 55944 19248 55956
rect 18739 55916 19248 55944
rect 18739 55913 18751 55916
rect 18693 55907 18751 55913
rect 19242 55904 19248 55916
rect 19300 55904 19306 55956
rect 19426 55904 19432 55956
rect 19484 55944 19490 55956
rect 19705 55947 19763 55953
rect 19705 55944 19717 55947
rect 19484 55916 19717 55944
rect 19484 55904 19490 55916
rect 19705 55913 19717 55916
rect 19751 55913 19763 55947
rect 19705 55907 19763 55913
rect 25130 55904 25136 55956
rect 25188 55944 25194 55956
rect 37826 55944 37832 55956
rect 25188 55916 37832 55944
rect 25188 55904 25194 55916
rect 37826 55904 37832 55916
rect 37884 55904 37890 55956
rect 26421 55879 26479 55885
rect 26421 55845 26433 55879
rect 26467 55876 26479 55879
rect 28442 55876 28448 55888
rect 26467 55848 28448 55876
rect 26467 55845 26479 55848
rect 26421 55839 26479 55845
rect 28442 55836 28448 55848
rect 28500 55836 28506 55888
rect 17310 55768 17316 55820
rect 17368 55808 17374 55820
rect 20901 55811 20959 55817
rect 20901 55808 20913 55811
rect 17368 55780 20913 55808
rect 17368 55768 17374 55780
rect 20901 55777 20913 55780
rect 20947 55808 20959 55811
rect 21082 55808 21088 55820
rect 20947 55780 21088 55808
rect 20947 55777 20959 55780
rect 20901 55771 20959 55777
rect 21082 55768 21088 55780
rect 21140 55768 21146 55820
rect 17037 55743 17095 55749
rect 17037 55709 17049 55743
rect 17083 55740 17095 55743
rect 17126 55740 17132 55752
rect 17083 55712 17132 55740
rect 17083 55709 17095 55712
rect 17037 55703 17095 55709
rect 17126 55700 17132 55712
rect 17184 55700 17190 55752
rect 18509 55743 18567 55749
rect 18509 55740 18521 55743
rect 18064 55712 18521 55740
rect 18064 55616 18092 55712
rect 18509 55709 18521 55712
rect 18555 55709 18567 55743
rect 18509 55703 18567 55709
rect 19889 55743 19947 55749
rect 19889 55709 19901 55743
rect 19935 55740 19947 55743
rect 26237 55743 26295 55749
rect 19935 55712 20392 55740
rect 19935 55709 19947 55712
rect 19889 55703 19947 55709
rect 20364 55616 20392 55712
rect 26237 55709 26249 55743
rect 26283 55740 26295 55743
rect 26326 55740 26332 55752
rect 26283 55712 26332 55740
rect 26283 55709 26295 55712
rect 26237 55703 26295 55709
rect 26326 55700 26332 55712
rect 26384 55740 26390 55752
rect 26881 55743 26939 55749
rect 26881 55740 26893 55743
rect 26384 55712 26893 55740
rect 26384 55700 26390 55712
rect 26881 55709 26893 55712
rect 26927 55709 26939 55743
rect 26881 55703 26939 55709
rect 16206 55604 16212 55616
rect 16167 55576 16212 55604
rect 16206 55564 16212 55576
rect 16264 55564 16270 55616
rect 18046 55604 18052 55616
rect 18007 55576 18052 55604
rect 18046 55564 18052 55576
rect 18104 55564 18110 55616
rect 20346 55604 20352 55616
rect 20307 55576 20352 55604
rect 20346 55564 20352 55576
rect 20404 55564 20410 55616
rect 22554 55604 22560 55616
rect 22515 55576 22560 55604
rect 22554 55564 22560 55576
rect 22612 55564 22618 55616
rect 24857 55607 24915 55613
rect 24857 55573 24869 55607
rect 24903 55604 24915 55607
rect 24946 55604 24952 55616
rect 24903 55576 24952 55604
rect 24903 55573 24915 55576
rect 24857 55567 24915 55573
rect 24946 55564 24952 55576
rect 25004 55564 25010 55616
rect 25501 55607 25559 55613
rect 25501 55573 25513 55607
rect 25547 55604 25559 55607
rect 25590 55604 25596 55616
rect 25547 55576 25596 55604
rect 25547 55573 25559 55576
rect 25501 55567 25559 55573
rect 25590 55564 25596 55576
rect 25648 55604 25654 55616
rect 26142 55604 26148 55616
rect 25648 55576 26148 55604
rect 25648 55564 25654 55576
rect 26142 55564 26148 55576
rect 26200 55564 26206 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 18690 55360 18696 55412
rect 18748 55400 18754 55412
rect 19150 55400 19156 55412
rect 18748 55372 19156 55400
rect 18748 55360 18754 55372
rect 19150 55360 19156 55372
rect 19208 55400 19214 55412
rect 19521 55403 19579 55409
rect 19521 55400 19533 55403
rect 19208 55372 19533 55400
rect 19208 55360 19214 55372
rect 19521 55369 19533 55372
rect 19567 55369 19579 55403
rect 19521 55363 19579 55369
rect 17126 55332 17132 55344
rect 17087 55304 17132 55332
rect 17126 55292 17132 55304
rect 17184 55292 17190 55344
rect 18966 55332 18972 55344
rect 18927 55304 18972 55332
rect 18966 55292 18972 55304
rect 19024 55292 19030 55344
rect 58158 55128 58164 55140
rect 58119 55100 58164 55128
rect 58158 55088 58164 55100
rect 58216 55088 58222 55140
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 57882 53932 57888 53984
rect 57940 53972 57946 53984
rect 58161 53975 58219 53981
rect 58161 53972 58173 53975
rect 57940 53944 58173 53972
rect 57940 53932 57946 53944
rect 58161 53941 58173 53944
rect 58207 53941 58219 53975
rect 58161 53935 58219 53941
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 57882 52436 57888 52488
rect 57940 52476 57946 52488
rect 58161 52479 58219 52485
rect 58161 52476 58173 52479
rect 57940 52448 58173 52476
rect 57940 52436 57946 52448
rect 58161 52445 58173 52448
rect 58207 52445 58219 52479
rect 58161 52439 58219 52445
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 58158 51388 58164 51400
rect 58119 51360 58164 51388
rect 58158 51348 58164 51360
rect 58216 51348 58222 51400
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 58158 49756 58164 49768
rect 58119 49728 58164 49756
rect 58158 49716 58164 49728
rect 58216 49716 58222 49768
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 58158 48532 58164 48544
rect 58119 48504 58164 48532
rect 58158 48492 58164 48504
rect 58216 48492 58222 48544
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 15286 47540 15292 47592
rect 15344 47580 15350 47592
rect 33962 47580 33968 47592
rect 15344 47552 33968 47580
rect 15344 47540 15350 47552
rect 33962 47540 33968 47552
rect 34020 47540 34026 47592
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 58158 47036 58164 47048
rect 58119 47008 58164 47036
rect 58158 46996 58164 47008
rect 58216 46996 58222 47048
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 58158 45948 58164 45960
rect 58119 45920 58164 45948
rect 58158 45908 58164 45920
rect 58216 45908 58222 45960
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 58158 44248 58164 44260
rect 58119 44220 58164 44248
rect 58158 44208 58164 44220
rect 58216 44208 58222 44260
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 58158 43092 58164 43104
rect 58119 43064 58164 43092
rect 58158 43052 58164 43064
rect 58216 43052 58222 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 12802 42236 12808 42288
rect 12860 42276 12866 42288
rect 13081 42279 13139 42285
rect 13081 42276 13093 42279
rect 12860 42248 13093 42276
rect 12860 42236 12866 42248
rect 13081 42245 13093 42248
rect 13127 42245 13139 42279
rect 13081 42239 13139 42245
rect 12897 42211 12955 42217
rect 12897 42177 12909 42211
rect 12943 42208 12955 42211
rect 13814 42208 13820 42220
rect 12943 42180 13820 42208
rect 12943 42177 12955 42180
rect 12897 42171 12955 42177
rect 13814 42168 13820 42180
rect 13872 42168 13878 42220
rect 14918 42208 14924 42220
rect 14879 42180 14924 42208
rect 14918 42168 14924 42180
rect 14976 42168 14982 42220
rect 15105 42211 15163 42217
rect 15105 42177 15117 42211
rect 15151 42208 15163 42211
rect 16666 42208 16672 42220
rect 15151 42180 16672 42208
rect 15151 42177 15163 42180
rect 15105 42171 15163 42177
rect 16666 42168 16672 42180
rect 16724 42168 16730 42220
rect 13265 42007 13323 42013
rect 13265 41973 13277 42007
rect 13311 42004 13323 42007
rect 13354 42004 13360 42016
rect 13311 41976 13360 42004
rect 13311 41973 13323 41976
rect 13265 41967 13323 41973
rect 13354 41964 13360 41976
rect 13412 41964 13418 42016
rect 15289 42007 15347 42013
rect 15289 41973 15301 42007
rect 15335 42004 15347 42007
rect 15562 42004 15568 42016
rect 15335 41976 15568 42004
rect 15335 41973 15347 41976
rect 15289 41967 15347 41973
rect 15562 41964 15568 41976
rect 15620 41964 15626 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 15013 41667 15071 41673
rect 13188 41636 13768 41664
rect 13188 41605 13216 41636
rect 13173 41599 13231 41605
rect 13173 41565 13185 41599
rect 13219 41565 13231 41599
rect 13173 41559 13231 41565
rect 13265 41599 13323 41605
rect 13265 41565 13277 41599
rect 13311 41565 13323 41599
rect 13265 41559 13323 41565
rect 12158 41488 12164 41540
rect 12216 41528 12222 41540
rect 12253 41531 12311 41537
rect 12253 41528 12265 41531
rect 12216 41500 12265 41528
rect 12216 41488 12222 41500
rect 12253 41497 12265 41500
rect 12299 41497 12311 41531
rect 12253 41491 12311 41497
rect 12437 41531 12495 41537
rect 12437 41497 12449 41531
rect 12483 41528 12495 41531
rect 13280 41528 13308 41559
rect 13354 41556 13360 41608
rect 13412 41596 13418 41608
rect 13412 41568 13457 41596
rect 13412 41556 13418 41568
rect 13538 41556 13544 41608
rect 13596 41596 13602 41608
rect 13596 41568 13641 41596
rect 13596 41556 13602 41568
rect 13630 41528 13636 41540
rect 12483 41500 13216 41528
rect 13280 41500 13636 41528
rect 12483 41497 12495 41500
rect 12437 41491 12495 41497
rect 12069 41463 12127 41469
rect 12069 41429 12081 41463
rect 12115 41460 12127 41463
rect 12526 41460 12532 41472
rect 12115 41432 12532 41460
rect 12115 41429 12127 41432
rect 12069 41423 12127 41429
rect 12526 41420 12532 41432
rect 12584 41420 12590 41472
rect 12618 41420 12624 41472
rect 12676 41460 12682 41472
rect 12897 41463 12955 41469
rect 12897 41460 12909 41463
rect 12676 41432 12909 41460
rect 12676 41420 12682 41432
rect 12897 41429 12909 41432
rect 12943 41429 12955 41463
rect 13188 41460 13216 41500
rect 13630 41488 13636 41500
rect 13688 41488 13694 41540
rect 13740 41528 13768 41636
rect 15013 41633 15025 41667
rect 15059 41664 15071 41667
rect 15059 41636 15700 41664
rect 15059 41633 15071 41636
rect 15013 41627 15071 41633
rect 13814 41556 13820 41608
rect 13872 41596 13878 41608
rect 14645 41599 14703 41605
rect 14645 41596 14657 41599
rect 13872 41568 14657 41596
rect 13872 41556 13878 41568
rect 14645 41565 14657 41568
rect 14691 41596 14703 41599
rect 14918 41596 14924 41608
rect 14691 41568 14924 41596
rect 14691 41565 14703 41568
rect 14645 41559 14703 41565
rect 14918 41556 14924 41568
rect 14976 41556 14982 41608
rect 15378 41556 15384 41608
rect 15436 41596 15442 41608
rect 15672 41605 15700 41636
rect 15473 41599 15531 41605
rect 15473 41596 15485 41599
rect 15436 41568 15485 41596
rect 15436 41556 15442 41568
rect 15473 41565 15485 41568
rect 15519 41565 15531 41599
rect 15473 41559 15531 41565
rect 15657 41599 15715 41605
rect 15657 41565 15669 41599
rect 15703 41565 15715 41599
rect 15657 41559 15715 41565
rect 15746 41556 15752 41608
rect 15804 41596 15810 41608
rect 15887 41599 15945 41605
rect 15804 41568 15849 41596
rect 15804 41556 15810 41568
rect 15887 41565 15899 41599
rect 15933 41596 15945 41599
rect 16669 41599 16727 41605
rect 16669 41596 16681 41599
rect 15933 41568 16681 41596
rect 15933 41565 15945 41568
rect 15887 41559 15945 41565
rect 16669 41565 16681 41568
rect 16715 41596 16727 41599
rect 20162 41596 20168 41608
rect 16715 41568 20168 41596
rect 16715 41565 16727 41568
rect 16669 41559 16727 41565
rect 20162 41556 20168 41568
rect 20220 41556 20226 41608
rect 58158 41596 58164 41608
rect 58119 41568 58164 41596
rect 58158 41556 58164 41568
rect 58216 41556 58222 41608
rect 14829 41531 14887 41537
rect 13740 41500 14228 41528
rect 13814 41460 13820 41472
rect 13188 41432 13820 41460
rect 12897 41423 12955 41429
rect 13814 41420 13820 41432
rect 13872 41420 13878 41472
rect 14200 41469 14228 41500
rect 14829 41497 14841 41531
rect 14875 41528 14887 41531
rect 15194 41528 15200 41540
rect 14875 41500 15200 41528
rect 14875 41497 14887 41500
rect 14829 41491 14887 41497
rect 15194 41488 15200 41500
rect 15252 41488 15258 41540
rect 16117 41531 16175 41537
rect 16117 41497 16129 41531
rect 16163 41528 16175 41531
rect 16758 41528 16764 41540
rect 16163 41500 16764 41528
rect 16163 41497 16175 41500
rect 16117 41491 16175 41497
rect 16758 41488 16764 41500
rect 16816 41488 16822 41540
rect 18414 41488 18420 41540
rect 18472 41528 18478 41540
rect 19245 41531 19303 41537
rect 19245 41528 19257 41531
rect 18472 41500 19257 41528
rect 18472 41488 18478 41500
rect 19245 41497 19257 41500
rect 19291 41497 19303 41531
rect 19426 41528 19432 41540
rect 19387 41500 19432 41528
rect 19245 41491 19303 41497
rect 19426 41488 19432 41500
rect 19484 41488 19490 41540
rect 14185 41463 14243 41469
rect 14185 41429 14197 41463
rect 14231 41460 14243 41463
rect 17678 41460 17684 41472
rect 14231 41432 17684 41460
rect 14231 41429 14243 41432
rect 14185 41423 14243 41429
rect 17678 41420 17684 41432
rect 17736 41420 17742 41472
rect 19334 41420 19340 41472
rect 19392 41460 19398 41472
rect 19613 41463 19671 41469
rect 19613 41460 19625 41463
rect 19392 41432 19625 41460
rect 19392 41420 19398 41432
rect 19613 41429 19625 41432
rect 19659 41429 19671 41463
rect 19613 41423 19671 41429
rect 20165 41463 20223 41469
rect 20165 41429 20177 41463
rect 20211 41460 20223 41463
rect 20254 41460 20260 41472
rect 20211 41432 20260 41460
rect 20211 41429 20223 41432
rect 20165 41423 20223 41429
rect 20254 41420 20260 41432
rect 20312 41460 20318 41472
rect 20714 41460 20720 41472
rect 20312 41432 20720 41460
rect 20312 41420 20318 41432
rect 20714 41420 20720 41432
rect 20772 41420 20778 41472
rect 23474 41420 23480 41472
rect 23532 41460 23538 41472
rect 23569 41463 23627 41469
rect 23569 41460 23581 41463
rect 23532 41432 23581 41460
rect 23532 41420 23538 41432
rect 23569 41429 23581 41432
rect 23615 41429 23627 41463
rect 23569 41423 23627 41429
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 10410 41256 10416 41268
rect 9968 41228 10416 41256
rect 9968 41135 9996 41228
rect 10410 41216 10416 41228
rect 10468 41256 10474 41268
rect 11790 41256 11796 41268
rect 10468 41228 11796 41256
rect 10468 41216 10474 41228
rect 11790 41216 11796 41228
rect 11848 41216 11854 41268
rect 15562 41256 15568 41268
rect 15488 41228 15568 41256
rect 12526 41148 12532 41200
rect 12584 41188 12590 41200
rect 12584 41160 13308 41188
rect 12584 41148 12590 41160
rect 9858 41120 9864 41132
rect 9819 41092 9864 41120
rect 9858 41080 9864 41092
rect 9916 41080 9922 41132
rect 9966 41129 10024 41135
rect 9966 41095 9978 41129
rect 10012 41095 10024 41129
rect 10066 41123 10124 41129
rect 10066 41120 10078 41123
rect 9966 41089 10024 41095
rect 10060 41089 10078 41120
rect 10112 41089 10124 41123
rect 10060 41083 10124 41089
rect 10229 41123 10287 41129
rect 10229 41089 10241 41123
rect 10275 41120 10287 41123
rect 10962 41120 10968 41132
rect 10275 41092 10968 41120
rect 10275 41089 10287 41092
rect 10229 41083 10287 41089
rect 9674 40944 9680 40996
rect 9732 40984 9738 40996
rect 10060 40984 10088 41083
rect 10962 41080 10968 41092
rect 11020 41080 11026 41132
rect 13280 41129 13308 41160
rect 13081 41123 13139 41129
rect 13081 41089 13093 41123
rect 13127 41089 13139 41123
rect 13081 41083 13139 41089
rect 13173 41123 13231 41129
rect 13173 41089 13185 41123
rect 13219 41089 13231 41123
rect 13173 41083 13231 41089
rect 13265 41123 13323 41129
rect 13265 41089 13277 41123
rect 13311 41089 13323 41123
rect 13446 41120 13452 41132
rect 13407 41092 13452 41120
rect 13265 41083 13323 41089
rect 9732 40956 10088 40984
rect 10781 40987 10839 40993
rect 9732 40944 9738 40956
rect 10781 40953 10793 40987
rect 10827 40984 10839 40987
rect 13096 40984 13124 41083
rect 13188 41052 13216 41083
rect 13446 41080 13452 41092
rect 13504 41120 13510 41132
rect 15378 41120 15384 41132
rect 13504 41092 15384 41120
rect 13504 41080 13510 41092
rect 15378 41080 15384 41092
rect 15436 41080 15442 41132
rect 15488 41120 15516 41228
rect 15562 41216 15568 41228
rect 15620 41216 15626 41268
rect 21177 41259 21235 41265
rect 21177 41256 21189 41259
rect 16684 41228 21189 41256
rect 16684 41197 16712 41228
rect 16669 41191 16727 41197
rect 16669 41188 16681 41191
rect 15764 41160 16681 41188
rect 15544 41123 15602 41129
rect 15544 41120 15556 41123
rect 15488 41092 15556 41120
rect 15544 41089 15556 41092
rect 15590 41089 15602 41123
rect 15544 41083 15602 41089
rect 15644 41126 15702 41132
rect 15764 41129 15792 41160
rect 16669 41157 16681 41160
rect 16715 41157 16727 41191
rect 16669 41151 16727 41157
rect 19368 41191 19426 41197
rect 19368 41157 19380 41191
rect 19414 41188 19426 41191
rect 20073 41191 20131 41197
rect 20073 41188 20085 41191
rect 19414 41160 20085 41188
rect 19414 41157 19426 41160
rect 19368 41151 19426 41157
rect 20073 41157 20085 41160
rect 20119 41157 20131 41191
rect 20073 41151 20131 41157
rect 15644 41092 15656 41126
rect 15690 41092 15702 41126
rect 15644 41086 15702 41092
rect 15749 41123 15807 41129
rect 15749 41089 15761 41123
rect 15795 41089 15807 41123
rect 13630 41052 13636 41064
rect 13188 41024 13636 41052
rect 13630 41012 13636 41024
rect 13688 41052 13694 41064
rect 13688 41024 15516 41052
rect 13688 41012 13694 41024
rect 13906 40984 13912 40996
rect 10827 40956 13032 40984
rect 13096 40956 13912 40984
rect 10827 40953 10839 40956
rect 10781 40947 10839 40953
rect 8294 40876 8300 40928
rect 8352 40916 8358 40928
rect 9585 40919 9643 40925
rect 9585 40916 9597 40919
rect 8352 40888 9597 40916
rect 8352 40876 8358 40888
rect 9585 40885 9597 40888
rect 9631 40885 9643 40919
rect 9585 40879 9643 40885
rect 9858 40876 9864 40928
rect 9916 40916 9922 40928
rect 10796 40916 10824 40947
rect 9916 40888 10824 40916
rect 9916 40876 9922 40888
rect 11422 40876 11428 40928
rect 11480 40916 11486 40928
rect 12805 40919 12863 40925
rect 12805 40916 12817 40919
rect 11480 40888 12817 40916
rect 11480 40876 11486 40888
rect 12805 40885 12817 40888
rect 12851 40885 12863 40919
rect 13004 40916 13032 40956
rect 13906 40944 13912 40956
rect 13964 40944 13970 40996
rect 15488 40984 15516 41024
rect 15672 40984 15700 41086
rect 15749 41083 15807 41089
rect 19518 41080 19524 41132
rect 19576 41120 19582 41132
rect 20364 41129 20392 41228
rect 21177 41225 21189 41228
rect 21223 41256 21235 41259
rect 25314 41256 25320 41268
rect 21223 41228 25320 41256
rect 21223 41225 21235 41228
rect 21177 41219 21235 41225
rect 25314 41216 25320 41228
rect 25372 41216 25378 41268
rect 21821 41191 21879 41197
rect 21821 41157 21833 41191
rect 21867 41188 21879 41191
rect 23382 41188 23388 41200
rect 21867 41160 23388 41188
rect 21867 41157 21879 41160
rect 21821 41151 21879 41157
rect 23382 41148 23388 41160
rect 23440 41188 23446 41200
rect 24394 41188 24400 41200
rect 23440 41160 24400 41188
rect 23440 41148 23446 41160
rect 24394 41148 24400 41160
rect 24452 41148 24458 41200
rect 20454 41129 20512 41135
rect 19613 41123 19671 41129
rect 19613 41120 19625 41123
rect 19576 41092 19625 41120
rect 19576 41080 19582 41092
rect 19613 41089 19625 41092
rect 19659 41089 19671 41123
rect 19613 41083 19671 41089
rect 20349 41123 20407 41129
rect 20349 41089 20361 41123
rect 20395 41089 20407 41123
rect 20454 41120 20466 41129
rect 20349 41083 20407 41089
rect 20453 41095 20466 41120
rect 20500 41095 20512 41129
rect 20453 41089 20512 41095
rect 20554 41123 20612 41129
rect 20554 41089 20566 41123
rect 20600 41120 20612 41123
rect 20600 41092 20668 41120
rect 20600 41089 20612 41092
rect 20453 40996 20481 41089
rect 20554 41083 20612 41089
rect 20640 40996 20668 41092
rect 20714 41080 20720 41132
rect 20772 41120 20778 41132
rect 22005 41123 22063 41129
rect 20772 41092 20817 41120
rect 20772 41080 20778 41092
rect 22005 41089 22017 41123
rect 22051 41120 22063 41123
rect 22186 41120 22192 41132
rect 22051 41092 22192 41120
rect 22051 41089 22063 41092
rect 22005 41083 22063 41089
rect 22186 41080 22192 41092
rect 22244 41080 22250 41132
rect 22833 41123 22891 41129
rect 22833 41089 22845 41123
rect 22879 41089 22891 41123
rect 23014 41120 23020 41132
rect 22975 41092 23020 41120
rect 22833 41083 22891 41089
rect 22848 41052 22876 41083
rect 23014 41080 23020 41092
rect 23072 41080 23078 41132
rect 23106 41080 23112 41132
rect 23164 41120 23170 41132
rect 23247 41123 23305 41129
rect 23164 41092 23209 41120
rect 23164 41080 23170 41092
rect 23247 41089 23259 41123
rect 23293 41120 23305 41123
rect 23658 41120 23664 41132
rect 23293 41092 23664 41120
rect 23293 41089 23305 41092
rect 23247 41083 23305 41089
rect 23658 41080 23664 41092
rect 23716 41080 23722 41132
rect 22922 41052 22928 41064
rect 22848 41024 22928 41052
rect 22922 41012 22928 41024
rect 22980 41012 22986 41064
rect 15746 40984 15752 40996
rect 15488 40956 15752 40984
rect 15746 40944 15752 40956
rect 15804 40944 15810 40996
rect 16025 40987 16083 40993
rect 16025 40953 16037 40987
rect 16071 40984 16083 40987
rect 17770 40984 17776 40996
rect 16071 40956 17776 40984
rect 16071 40953 16083 40956
rect 16025 40947 16083 40953
rect 17770 40944 17776 40956
rect 17828 40944 17834 40996
rect 20438 40944 20444 40996
rect 20496 40944 20502 40996
rect 20622 40944 20628 40996
rect 20680 40944 20686 40996
rect 23290 40984 23296 40996
rect 22112 40956 23296 40984
rect 15010 40916 15016 40928
rect 13004 40888 15016 40916
rect 12805 40879 12863 40885
rect 15010 40876 15016 40888
rect 15068 40876 15074 40928
rect 17494 40876 17500 40928
rect 17552 40916 17558 40928
rect 18233 40919 18291 40925
rect 18233 40916 18245 40919
rect 17552 40888 18245 40916
rect 17552 40876 17558 40888
rect 18233 40885 18245 40888
rect 18279 40885 18291 40919
rect 18233 40879 18291 40885
rect 18598 40876 18604 40928
rect 18656 40916 18662 40928
rect 22112 40916 22140 40956
rect 23290 40944 23296 40956
rect 23348 40984 23354 40996
rect 23937 40987 23995 40993
rect 23937 40984 23949 40987
rect 23348 40956 23949 40984
rect 23348 40944 23354 40956
rect 23937 40953 23949 40956
rect 23983 40953 23995 40987
rect 23937 40947 23995 40953
rect 18656 40888 22140 40916
rect 22189 40919 22247 40925
rect 18656 40876 18662 40888
rect 22189 40885 22201 40919
rect 22235 40916 22247 40919
rect 22278 40916 22284 40928
rect 22235 40888 22284 40916
rect 22235 40885 22247 40888
rect 22189 40879 22247 40885
rect 22278 40876 22284 40888
rect 22336 40876 22342 40928
rect 23474 40916 23480 40928
rect 23435 40888 23480 40916
rect 23474 40876 23480 40888
rect 23532 40876 23538 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 11517 40715 11575 40721
rect 11517 40681 11529 40715
rect 11563 40712 11575 40715
rect 12158 40712 12164 40724
rect 11563 40684 12164 40712
rect 11563 40681 11575 40684
rect 11517 40675 11575 40681
rect 12158 40672 12164 40684
rect 12216 40672 12222 40724
rect 18693 40715 18751 40721
rect 18693 40681 18705 40715
rect 18739 40712 18751 40715
rect 20622 40712 20628 40724
rect 18739 40684 20628 40712
rect 18739 40681 18751 40684
rect 18693 40675 18751 40681
rect 20622 40672 20628 40684
rect 20680 40672 20686 40724
rect 23014 40672 23020 40724
rect 23072 40712 23078 40724
rect 24765 40715 24823 40721
rect 24765 40712 24777 40715
rect 23072 40684 24777 40712
rect 23072 40672 23078 40684
rect 24765 40681 24777 40684
rect 24811 40681 24823 40715
rect 24765 40675 24823 40681
rect 22094 40604 22100 40656
rect 22152 40644 22158 40656
rect 23106 40644 23112 40656
rect 22152 40616 23112 40644
rect 22152 40604 22158 40616
rect 23106 40604 23112 40616
rect 23164 40604 23170 40656
rect 20254 40576 20260 40588
rect 19260 40548 20260 40576
rect 5169 40511 5227 40517
rect 5169 40477 5181 40511
rect 5215 40508 5227 40511
rect 5258 40508 5264 40520
rect 5215 40480 5264 40508
rect 5215 40477 5227 40480
rect 5169 40471 5227 40477
rect 5258 40468 5264 40480
rect 5316 40468 5322 40520
rect 9858 40468 9864 40520
rect 9916 40508 9922 40520
rect 10137 40511 10195 40517
rect 10137 40508 10149 40511
rect 9916 40480 10149 40508
rect 9916 40468 9922 40480
rect 10137 40477 10149 40480
rect 10183 40477 10195 40511
rect 10137 40471 10195 40477
rect 10404 40511 10462 40517
rect 10404 40477 10416 40511
rect 10450 40508 10462 40511
rect 11422 40508 11428 40520
rect 10450 40480 11428 40508
rect 10450 40477 10462 40480
rect 10404 40471 10462 40477
rect 11422 40468 11428 40480
rect 11480 40468 11486 40520
rect 11977 40511 12035 40517
rect 11977 40477 11989 40511
rect 12023 40508 12035 40511
rect 12244 40511 12302 40517
rect 12023 40480 12112 40508
rect 12023 40477 12035 40480
rect 11977 40471 12035 40477
rect 5436 40443 5494 40449
rect 5436 40409 5448 40443
rect 5482 40440 5494 40443
rect 5626 40440 5632 40452
rect 5482 40412 5632 40440
rect 5482 40409 5494 40412
rect 5436 40403 5494 40409
rect 5626 40400 5632 40412
rect 5684 40400 5690 40452
rect 6454 40400 6460 40452
rect 6512 40440 6518 40452
rect 6512 40412 7236 40440
rect 6512 40400 6518 40412
rect 6546 40372 6552 40384
rect 6507 40344 6552 40372
rect 6546 40332 6552 40344
rect 6604 40332 6610 40384
rect 7208 40381 7236 40412
rect 7193 40375 7251 40381
rect 7193 40341 7205 40375
rect 7239 40372 7251 40375
rect 7558 40372 7564 40384
rect 7239 40344 7564 40372
rect 7239 40341 7251 40344
rect 7193 40335 7251 40341
rect 7558 40332 7564 40344
rect 7616 40332 7622 40384
rect 12084 40372 12112 40480
rect 12244 40477 12256 40511
rect 12290 40508 12302 40511
rect 12618 40508 12624 40520
rect 12290 40480 12624 40508
rect 12290 40477 12302 40480
rect 12244 40471 12302 40477
rect 12618 40468 12624 40480
rect 12676 40468 12682 40520
rect 13722 40468 13728 40520
rect 13780 40508 13786 40520
rect 14461 40511 14519 40517
rect 14461 40508 14473 40511
rect 13780 40480 14473 40508
rect 13780 40468 13786 40480
rect 14461 40477 14473 40480
rect 14507 40477 14519 40511
rect 14461 40471 14519 40477
rect 16574 40468 16580 40520
rect 16632 40508 16638 40520
rect 17405 40511 17463 40517
rect 17405 40508 17417 40511
rect 16632 40480 17417 40508
rect 16632 40468 16638 40480
rect 17405 40477 17417 40480
rect 17451 40477 17463 40511
rect 17405 40471 17463 40477
rect 17494 40468 17500 40520
rect 17552 40508 17558 40520
rect 19260 40517 19288 40548
rect 20254 40536 20260 40548
rect 20312 40536 20318 40588
rect 23124 40576 23152 40604
rect 23124 40548 23244 40576
rect 18509 40511 18567 40517
rect 18509 40508 18521 40511
rect 17552 40480 18521 40508
rect 17552 40468 17558 40480
rect 18509 40477 18521 40480
rect 18555 40477 18567 40511
rect 18509 40471 18567 40477
rect 19245 40511 19303 40517
rect 19245 40477 19257 40511
rect 19291 40477 19303 40511
rect 19245 40471 19303 40477
rect 19334 40468 19340 40520
rect 19392 40508 19398 40520
rect 19429 40511 19487 40517
rect 19429 40508 19441 40511
rect 19392 40480 19441 40508
rect 19392 40468 19398 40480
rect 19429 40477 19441 40480
rect 19475 40477 19487 40511
rect 19429 40471 19487 40477
rect 19521 40511 19579 40517
rect 19521 40477 19533 40511
rect 19567 40477 19579 40511
rect 19521 40471 19579 40477
rect 19613 40511 19671 40517
rect 19613 40477 19625 40511
rect 19659 40508 19671 40511
rect 20070 40508 20076 40520
rect 19659 40480 20076 40508
rect 19659 40477 19671 40480
rect 19613 40471 19671 40477
rect 13814 40400 13820 40452
rect 13872 40440 13878 40452
rect 14274 40440 14280 40452
rect 13872 40412 14280 40440
rect 13872 40400 13878 40412
rect 14274 40400 14280 40412
rect 14332 40400 14338 40452
rect 16758 40400 16764 40452
rect 16816 40440 16822 40452
rect 17138 40443 17196 40449
rect 17138 40440 17150 40443
rect 16816 40412 17150 40440
rect 16816 40400 16822 40412
rect 17138 40409 17150 40412
rect 17184 40409 17196 40443
rect 17138 40403 17196 40409
rect 18325 40443 18383 40449
rect 18325 40409 18337 40443
rect 18371 40440 18383 40443
rect 18414 40440 18420 40452
rect 18371 40412 18420 40440
rect 18371 40409 18383 40412
rect 18325 40403 18383 40409
rect 18414 40400 18420 40412
rect 18472 40400 18478 40452
rect 19536 40440 19564 40471
rect 20070 40468 20076 40480
rect 20128 40468 20134 40520
rect 20622 40468 20628 40520
rect 20680 40508 20686 40520
rect 20809 40511 20867 40517
rect 20809 40508 20821 40511
rect 20680 40480 20821 40508
rect 20680 40468 20686 40480
rect 20809 40477 20821 40480
rect 20855 40477 20867 40511
rect 22922 40508 22928 40520
rect 22883 40480 22928 40508
rect 20809 40471 20867 40477
rect 22922 40468 22928 40480
rect 22980 40468 22986 40520
rect 23216 40517 23244 40548
rect 23109 40511 23167 40517
rect 23109 40477 23121 40511
rect 23155 40477 23167 40511
rect 23109 40471 23167 40477
rect 23204 40511 23262 40517
rect 23204 40477 23216 40511
rect 23250 40477 23262 40511
rect 23204 40471 23262 40477
rect 20438 40440 20444 40452
rect 19536 40412 20444 40440
rect 20438 40400 20444 40412
rect 20496 40400 20502 40452
rect 21076 40443 21134 40449
rect 21076 40409 21088 40443
rect 21122 40440 21134 40443
rect 21818 40440 21824 40452
rect 21122 40412 21824 40440
rect 21122 40409 21134 40412
rect 21076 40403 21134 40409
rect 21818 40400 21824 40412
rect 21876 40400 21882 40452
rect 23014 40400 23020 40452
rect 23072 40440 23078 40452
rect 23124 40440 23152 40471
rect 23290 40468 23296 40520
rect 23348 40517 23354 40520
rect 23348 40511 23371 40517
rect 23359 40477 23371 40511
rect 23348 40471 23371 40477
rect 30929 40511 30987 40517
rect 30929 40477 30941 40511
rect 30975 40508 30987 40511
rect 32214 40508 32220 40520
rect 30975 40480 32220 40508
rect 30975 40477 30987 40480
rect 30929 40471 30987 40477
rect 23348 40468 23354 40471
rect 32214 40468 32220 40480
rect 32272 40468 32278 40520
rect 58158 40508 58164 40520
rect 58119 40480 58164 40508
rect 58158 40468 58164 40480
rect 58216 40468 58222 40520
rect 24394 40440 24400 40452
rect 23072 40412 23152 40440
rect 24355 40412 24400 40440
rect 23072 40400 23078 40412
rect 24394 40400 24400 40412
rect 24452 40400 24458 40452
rect 24581 40443 24639 40449
rect 24581 40409 24593 40443
rect 24627 40440 24639 40443
rect 24854 40440 24860 40452
rect 24627 40412 24860 40440
rect 24627 40409 24639 40412
rect 24581 40403 24639 40409
rect 24854 40400 24860 40412
rect 24912 40400 24918 40452
rect 30834 40400 30840 40452
rect 30892 40440 30898 40452
rect 31174 40443 31232 40449
rect 31174 40440 31186 40443
rect 30892 40412 31186 40440
rect 30892 40400 30898 40412
rect 31174 40409 31186 40412
rect 31220 40409 31232 40443
rect 31174 40403 31232 40409
rect 12342 40372 12348 40384
rect 12084 40344 12348 40372
rect 12342 40332 12348 40344
rect 12400 40332 12406 40384
rect 12802 40332 12808 40384
rect 12860 40372 12866 40384
rect 13357 40375 13415 40381
rect 13357 40372 13369 40375
rect 12860 40344 13369 40372
rect 12860 40332 12866 40344
rect 13357 40341 13369 40344
rect 13403 40341 13415 40375
rect 13357 40335 13415 40341
rect 14645 40375 14703 40381
rect 14645 40341 14657 40375
rect 14691 40372 14703 40375
rect 14918 40372 14924 40384
rect 14691 40344 14924 40372
rect 14691 40341 14703 40344
rect 14645 40335 14703 40341
rect 14918 40332 14924 40344
rect 14976 40332 14982 40384
rect 15194 40332 15200 40384
rect 15252 40372 15258 40384
rect 16022 40372 16028 40384
rect 15252 40344 16028 40372
rect 15252 40332 15258 40344
rect 16022 40332 16028 40344
rect 16080 40332 16086 40384
rect 19889 40375 19947 40381
rect 19889 40341 19901 40375
rect 19935 40372 19947 40375
rect 20346 40372 20352 40384
rect 19935 40344 20352 40372
rect 19935 40341 19947 40344
rect 19889 40335 19947 40341
rect 20346 40332 20352 40344
rect 20404 40332 20410 40384
rect 22186 40372 22192 40384
rect 22099 40344 22192 40372
rect 22186 40332 22192 40344
rect 22244 40372 22250 40384
rect 22646 40372 22652 40384
rect 22244 40344 22652 40372
rect 22244 40332 22250 40344
rect 22646 40332 22652 40344
rect 22704 40332 22710 40384
rect 23566 40372 23572 40384
rect 23527 40344 23572 40372
rect 23566 40332 23572 40344
rect 23624 40332 23630 40384
rect 32030 40332 32036 40384
rect 32088 40372 32094 40384
rect 32309 40375 32367 40381
rect 32309 40372 32321 40375
rect 32088 40344 32321 40372
rect 32088 40332 32094 40344
rect 32309 40341 32321 40344
rect 32355 40341 32367 40375
rect 32309 40335 32367 40341
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 3881 40171 3939 40177
rect 3881 40137 3893 40171
rect 3927 40137 3939 40171
rect 3881 40131 3939 40137
rect 3896 40100 3924 40131
rect 4982 40128 4988 40180
rect 5040 40168 5046 40180
rect 10689 40171 10747 40177
rect 5040 40140 7052 40168
rect 5040 40128 5046 40140
rect 4525 40103 4583 40109
rect 4525 40100 4537 40103
rect 3896 40072 4537 40100
rect 4525 40069 4537 40072
rect 4571 40100 4583 40103
rect 5534 40100 5540 40112
rect 4571 40072 5540 40100
rect 4571 40069 4583 40072
rect 4525 40063 4583 40069
rect 5534 40060 5540 40072
rect 5592 40060 5598 40112
rect 2768 40035 2826 40041
rect 2768 40001 2780 40035
rect 2814 40032 2826 40035
rect 3786 40032 3792 40044
rect 2814 40004 3792 40032
rect 2814 40001 2826 40004
rect 2768 39995 2826 40001
rect 3786 39992 3792 40004
rect 3844 39992 3850 40044
rect 4709 40035 4767 40041
rect 4709 40001 4721 40035
rect 4755 40032 4767 40035
rect 4798 40032 4804 40044
rect 4755 40004 4804 40032
rect 4755 40001 4767 40004
rect 4709 39995 4767 40001
rect 4798 39992 4804 40004
rect 4856 39992 4862 40044
rect 6454 39992 6460 40044
rect 6512 40032 6518 40044
rect 6595 40035 6653 40041
rect 6595 40032 6607 40035
rect 6512 40004 6607 40032
rect 6512 39992 6518 40004
rect 6595 40001 6607 40004
rect 6641 40001 6653 40035
rect 6595 39995 6653 40001
rect 6730 40035 6788 40041
rect 6730 40001 6742 40035
rect 6776 40001 6788 40035
rect 6730 39995 6788 40001
rect 2498 39964 2504 39976
rect 2459 39936 2504 39964
rect 2498 39924 2504 39936
rect 2556 39924 2562 39976
rect 6748 39908 6776 39995
rect 6822 39992 6828 40044
rect 6880 40041 6886 40044
rect 7024 40041 7052 40140
rect 10689 40137 10701 40171
rect 10735 40168 10747 40171
rect 11330 40168 11336 40180
rect 10735 40140 11336 40168
rect 10735 40137 10747 40140
rect 10689 40131 10747 40137
rect 11330 40128 11336 40140
rect 11388 40128 11394 40180
rect 13722 40128 13728 40180
rect 13780 40168 13786 40180
rect 14001 40171 14059 40177
rect 14001 40168 14013 40171
rect 13780 40140 14013 40168
rect 13780 40128 13786 40140
rect 14001 40137 14013 40140
rect 14047 40137 14059 40171
rect 14001 40131 14059 40137
rect 15010 40128 15016 40180
rect 15068 40168 15074 40180
rect 21177 40171 21235 40177
rect 21177 40168 21189 40171
rect 15068 40140 21189 40168
rect 15068 40128 15074 40140
rect 21177 40137 21189 40140
rect 21223 40168 21235 40171
rect 21450 40168 21456 40180
rect 21223 40140 21456 40168
rect 21223 40137 21235 40140
rect 21177 40131 21235 40137
rect 21450 40128 21456 40140
rect 21508 40128 21514 40180
rect 21818 40168 21824 40180
rect 21779 40140 21824 40168
rect 21818 40128 21824 40140
rect 21876 40128 21882 40180
rect 22094 40128 22100 40180
rect 22152 40168 22158 40180
rect 22925 40171 22983 40177
rect 22152 40140 22232 40168
rect 22152 40128 22158 40140
rect 9858 40100 9864 40112
rect 9508 40072 9864 40100
rect 7742 40041 7748 40044
rect 6880 40032 6888 40041
rect 7009 40035 7067 40041
rect 6880 40004 6925 40032
rect 6880 39995 6888 40004
rect 7009 40001 7021 40035
rect 7055 40001 7067 40035
rect 7009 39995 7067 40001
rect 7469 40035 7527 40041
rect 7469 40001 7481 40035
rect 7515 40001 7527 40035
rect 7736 40032 7748 40041
rect 7703 40004 7748 40032
rect 7469 39995 7527 40001
rect 7736 39995 7748 40004
rect 6880 39992 6886 39995
rect 5810 39896 5816 39908
rect 5723 39868 5816 39896
rect 5810 39856 5816 39868
rect 5868 39896 5874 39908
rect 6638 39896 6644 39908
rect 5868 39868 6644 39896
rect 5868 39856 5874 39868
rect 6638 39856 6644 39868
rect 6696 39856 6702 39908
rect 6730 39856 6736 39908
rect 6788 39856 6794 39908
rect 4341 39831 4399 39837
rect 4341 39797 4353 39831
rect 4387 39828 4399 39831
rect 4614 39828 4620 39840
rect 4387 39800 4620 39828
rect 4387 39797 4399 39800
rect 4341 39791 4399 39797
rect 4614 39788 4620 39800
rect 4672 39788 4678 39840
rect 5258 39828 5264 39840
rect 5219 39800 5264 39828
rect 5258 39788 5264 39800
rect 5316 39788 5322 39840
rect 6362 39828 6368 39840
rect 6323 39800 6368 39828
rect 6362 39788 6368 39800
rect 6420 39788 6426 39840
rect 7484 39828 7512 39995
rect 7742 39992 7748 39995
rect 7800 39992 7806 40044
rect 9309 40035 9367 40041
rect 9309 40001 9321 40035
rect 9355 40032 9367 40035
rect 9508 40032 9536 40072
rect 9858 40060 9864 40072
rect 9916 40060 9922 40112
rect 18414 40060 18420 40112
rect 18472 40100 18478 40112
rect 19242 40100 19248 40112
rect 18472 40072 19248 40100
rect 18472 40060 18478 40072
rect 19242 40060 19248 40072
rect 19300 40060 19306 40112
rect 20073 40103 20131 40109
rect 20073 40069 20085 40103
rect 20119 40069 20131 40103
rect 20073 40063 20131 40069
rect 9355 40004 9536 40032
rect 9576 40035 9634 40041
rect 9355 40001 9367 40004
rect 9309 39995 9367 40001
rect 9576 40001 9588 40035
rect 9622 40032 9634 40035
rect 9622 40004 10916 40032
rect 9622 40001 9634 40004
rect 9576 39995 9634 40001
rect 9324 39896 9352 39995
rect 8404 39868 9352 39896
rect 8404 39828 8432 39868
rect 8846 39828 8852 39840
rect 7484 39800 8432 39828
rect 8807 39800 8852 39828
rect 8846 39788 8852 39800
rect 8904 39788 8910 39840
rect 10888 39828 10916 40004
rect 10962 39992 10968 40044
rect 11020 40032 11026 40044
rect 11517 40035 11575 40041
rect 11517 40032 11529 40035
rect 11020 40004 11529 40032
rect 11020 39992 11026 40004
rect 11517 40001 11529 40004
rect 11563 40001 11575 40035
rect 11680 40035 11738 40041
rect 11680 40032 11692 40035
rect 11517 39995 11575 40001
rect 11624 40004 11692 40032
rect 11514 39856 11520 39908
rect 11572 39896 11578 39908
rect 11624 39896 11652 40004
rect 11680 40001 11692 40004
rect 11726 40001 11738 40035
rect 11680 39995 11738 40001
rect 11790 39992 11796 40044
rect 11848 40032 11854 40044
rect 11931 40035 11989 40041
rect 11848 40004 11893 40032
rect 11848 39992 11854 40004
rect 11931 40001 11943 40035
rect 11977 40032 11989 40035
rect 12618 40032 12624 40044
rect 11977 40004 12624 40032
rect 11977 40001 11989 40004
rect 11931 39995 11989 40001
rect 12618 39992 12624 40004
rect 12676 39992 12682 40044
rect 14550 39992 14556 40044
rect 14608 40032 14614 40044
rect 15114 40035 15172 40041
rect 15114 40032 15126 40035
rect 14608 40004 15126 40032
rect 14608 39992 14614 40004
rect 15114 40001 15126 40004
rect 15160 40001 15172 40035
rect 20088 40032 20116 40063
rect 15114 39995 15172 40001
rect 17788 40004 20116 40032
rect 15381 39967 15439 39973
rect 15381 39933 15393 39967
rect 15427 39964 15439 39967
rect 15654 39964 15660 39976
rect 15427 39936 15660 39964
rect 15427 39933 15439 39936
rect 15381 39927 15439 39933
rect 15654 39924 15660 39936
rect 15712 39964 15718 39976
rect 16482 39964 16488 39976
rect 15712 39936 16488 39964
rect 15712 39924 15718 39936
rect 16482 39924 16488 39936
rect 16540 39924 16546 39976
rect 11572 39868 11652 39896
rect 11572 39856 11578 39868
rect 11790 39856 11796 39908
rect 11848 39896 11854 39908
rect 11848 39868 14504 39896
rect 11848 39856 11854 39868
rect 12161 39831 12219 39837
rect 12161 39828 12173 39831
rect 10888 39800 12173 39828
rect 12161 39797 12173 39800
rect 12207 39797 12219 39831
rect 12618 39828 12624 39840
rect 12579 39800 12624 39828
rect 12161 39791 12219 39797
rect 12618 39788 12624 39800
rect 12676 39788 12682 39840
rect 14476 39828 14504 39868
rect 17788 39837 17816 40004
rect 21450 39992 21456 40044
rect 21508 40032 21514 40044
rect 22204 40041 22232 40140
rect 22925 40137 22937 40171
rect 22971 40168 22983 40171
rect 23014 40168 23020 40180
rect 22971 40140 23020 40168
rect 22971 40137 22983 40140
rect 22925 40131 22983 40137
rect 23014 40128 23020 40140
rect 23072 40128 23078 40180
rect 23382 40168 23388 40180
rect 23308 40140 23388 40168
rect 23308 40109 23336 40140
rect 23382 40128 23388 40140
rect 23440 40128 23446 40180
rect 23750 40128 23756 40180
rect 23808 40168 23814 40180
rect 25225 40171 25283 40177
rect 25225 40168 25237 40171
rect 23808 40140 25237 40168
rect 23808 40128 23814 40140
rect 25225 40137 25237 40140
rect 25271 40137 25283 40171
rect 25225 40131 25283 40137
rect 28721 40171 28779 40177
rect 28721 40137 28733 40171
rect 28767 40168 28779 40171
rect 29178 40168 29184 40180
rect 28767 40140 29184 40168
rect 28767 40137 28779 40140
rect 28721 40131 28779 40137
rect 29178 40128 29184 40140
rect 29236 40128 29242 40180
rect 23293 40103 23351 40109
rect 23293 40069 23305 40103
rect 23339 40069 23351 40103
rect 23293 40063 23351 40069
rect 23566 40060 23572 40112
rect 23624 40100 23630 40112
rect 24090 40103 24148 40109
rect 24090 40100 24102 40103
rect 23624 40072 24102 40100
rect 23624 40060 23630 40072
rect 24090 40069 24102 40072
rect 24136 40069 24148 40103
rect 24090 40063 24148 40069
rect 22077 40035 22135 40041
rect 21928 40032 22048 40035
rect 22077 40032 22089 40035
rect 21508 40007 22089 40032
rect 21508 40004 21956 40007
rect 22020 40004 22089 40007
rect 21508 39992 21514 40004
rect 22077 40001 22089 40004
rect 22123 40001 22135 40035
rect 22077 39995 22135 40001
rect 22170 40035 22232 40041
rect 22170 40001 22182 40035
rect 22216 40004 22232 40035
rect 22216 40001 22228 40004
rect 22170 39995 22228 40001
rect 22278 39992 22284 40044
rect 22336 40032 22342 40044
rect 22465 40035 22523 40041
rect 22336 40004 22381 40032
rect 22336 39992 22342 40004
rect 22465 40001 22477 40035
rect 22511 40032 22523 40035
rect 22922 40032 22928 40044
rect 22511 40004 22928 40032
rect 22511 40001 22523 40004
rect 22465 39995 22523 40001
rect 18322 39964 18328 39976
rect 18283 39936 18328 39964
rect 18322 39924 18328 39936
rect 18380 39964 18386 39976
rect 19426 39964 19432 39976
rect 18380 39936 19432 39964
rect 18380 39924 18386 39936
rect 19426 39924 19432 39936
rect 19484 39924 19490 39976
rect 22480 39964 22508 39995
rect 22922 39992 22928 40004
rect 22980 39992 22986 40044
rect 23109 40035 23167 40041
rect 23109 40001 23121 40035
rect 23155 40001 23167 40035
rect 23109 39995 23167 40001
rect 22204 39936 22508 39964
rect 22204 39908 22232 39936
rect 20070 39856 20076 39908
rect 20128 39896 20134 39908
rect 20625 39899 20683 39905
rect 20625 39896 20637 39899
rect 20128 39868 20637 39896
rect 20128 39856 20134 39868
rect 20625 39865 20637 39868
rect 20671 39896 20683 39899
rect 20671 39868 22094 39896
rect 20671 39865 20683 39868
rect 20625 39859 20683 39865
rect 17773 39831 17831 39837
rect 17773 39828 17785 39831
rect 14476 39800 17785 39828
rect 17773 39797 17785 39800
rect 17819 39797 17831 39831
rect 22066 39828 22094 39868
rect 22186 39856 22192 39908
rect 22244 39856 22250 39908
rect 23124 39896 23152 39995
rect 23382 39992 23388 40044
rect 23440 40032 23446 40044
rect 23658 40032 23664 40044
rect 23440 40004 23664 40032
rect 23440 39992 23446 40004
rect 23658 39992 23664 40004
rect 23716 39992 23722 40044
rect 27608 40035 27666 40041
rect 27608 40001 27620 40035
rect 27654 40032 27666 40035
rect 28350 40032 28356 40044
rect 27654 40004 28356 40032
rect 27654 40001 27666 40004
rect 27608 39995 27666 40001
rect 28350 39992 28356 40004
rect 28408 39992 28414 40044
rect 23842 39964 23848 39976
rect 23803 39936 23848 39964
rect 23842 39924 23848 39936
rect 23900 39924 23906 39976
rect 27341 39967 27399 39973
rect 27341 39933 27353 39967
rect 27387 39933 27399 39967
rect 27341 39927 27399 39933
rect 23198 39896 23204 39908
rect 23111 39868 23204 39896
rect 23198 39856 23204 39868
rect 23256 39896 23262 39908
rect 23750 39896 23756 39908
rect 23256 39868 23756 39896
rect 23256 39856 23262 39868
rect 23750 39856 23756 39868
rect 23808 39856 23814 39908
rect 25222 39828 25228 39840
rect 22066 39800 25228 39828
rect 17773 39791 17831 39797
rect 25222 39788 25228 39800
rect 25280 39788 25286 39840
rect 27356 39828 27384 39927
rect 27614 39828 27620 39840
rect 27356 39800 27620 39828
rect 27614 39788 27620 39800
rect 27672 39788 27678 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 3786 39624 3792 39636
rect 3747 39596 3792 39624
rect 3786 39584 3792 39596
rect 3844 39584 3850 39636
rect 4614 39584 4620 39636
rect 4672 39584 4678 39636
rect 5626 39624 5632 39636
rect 5587 39596 5632 39624
rect 5626 39584 5632 39596
rect 5684 39584 5690 39636
rect 6730 39624 6736 39636
rect 5736 39596 6736 39624
rect 4632 39556 4660 39584
rect 5350 39556 5356 39568
rect 4264 39528 4660 39556
rect 5263 39528 5356 39556
rect 4264 39429 4292 39528
rect 5276 39488 5304 39528
rect 5350 39516 5356 39528
rect 5408 39556 5414 39568
rect 5736 39556 5764 39596
rect 6730 39584 6736 39596
rect 6788 39584 6794 39636
rect 11514 39624 11520 39636
rect 11475 39596 11520 39624
rect 11514 39584 11520 39596
rect 11572 39584 11578 39636
rect 14461 39627 14519 39633
rect 14461 39593 14473 39627
rect 14507 39624 14519 39627
rect 14550 39624 14556 39636
rect 14507 39596 14556 39624
rect 14507 39593 14519 39596
rect 14461 39587 14519 39593
rect 14550 39584 14556 39596
rect 14608 39584 14614 39636
rect 19245 39627 19303 39633
rect 19245 39593 19257 39627
rect 19291 39624 19303 39627
rect 19334 39624 19340 39636
rect 19291 39596 19340 39624
rect 19291 39593 19303 39596
rect 19245 39587 19303 39593
rect 19334 39584 19340 39596
rect 19392 39584 19398 39636
rect 30834 39624 30840 39636
rect 30795 39596 30840 39624
rect 30834 39584 30840 39596
rect 30892 39584 30898 39636
rect 5408 39528 5764 39556
rect 5408 39516 5414 39528
rect 4356 39460 5304 39488
rect 4065 39423 4123 39429
rect 4065 39389 4077 39423
rect 4111 39389 4123 39423
rect 4065 39383 4123 39389
rect 4157 39423 4215 39429
rect 4157 39389 4169 39423
rect 4203 39389 4215 39423
rect 4157 39383 4215 39389
rect 4249 39423 4307 39429
rect 4249 39389 4261 39423
rect 4295 39389 4307 39423
rect 4249 39383 4307 39389
rect 4080 39284 4108 39383
rect 4172 39352 4200 39383
rect 4356 39352 4384 39460
rect 4433 39423 4491 39429
rect 4433 39389 4445 39423
rect 4479 39420 4491 39423
rect 4982 39420 4988 39432
rect 4479 39392 4988 39420
rect 4479 39389 4491 39392
rect 4433 39383 4491 39389
rect 4982 39380 4988 39392
rect 5040 39380 5046 39432
rect 5276 39429 5304 39460
rect 5442 39448 5448 39500
rect 5500 39488 5506 39500
rect 6089 39491 6147 39497
rect 6089 39488 6101 39491
rect 5500 39460 6101 39488
rect 5500 39448 5506 39460
rect 6089 39457 6101 39460
rect 6135 39457 6147 39491
rect 6089 39451 6147 39457
rect 12989 39491 13047 39497
rect 12989 39457 13001 39491
rect 13035 39488 13047 39491
rect 13446 39488 13452 39500
rect 13035 39460 13452 39488
rect 13035 39457 13047 39460
rect 12989 39451 13047 39457
rect 13446 39448 13452 39460
rect 13504 39488 13510 39500
rect 32309 39491 32367 39497
rect 32309 39488 32321 39491
rect 13504 39460 15148 39488
rect 13504 39448 13510 39460
rect 5169 39423 5227 39429
rect 5169 39389 5181 39423
rect 5215 39389 5227 39423
rect 5169 39383 5227 39389
rect 5261 39423 5319 39429
rect 5261 39389 5273 39423
rect 5307 39389 5319 39423
rect 5261 39383 5319 39389
rect 5353 39423 5411 39429
rect 5353 39389 5365 39423
rect 5399 39417 5411 39423
rect 5810 39420 5816 39432
rect 5460 39417 5816 39420
rect 5399 39392 5816 39417
rect 5399 39389 5488 39392
rect 5353 39383 5411 39389
rect 4172 39324 4384 39352
rect 5184 39352 5212 39383
rect 5810 39380 5816 39392
rect 5868 39380 5874 39432
rect 6362 39429 6368 39432
rect 6356 39420 6368 39429
rect 6323 39392 6368 39420
rect 6356 39383 6368 39392
rect 6362 39380 6368 39383
rect 6420 39380 6426 39432
rect 9309 39423 9367 39429
rect 9309 39389 9321 39423
rect 9355 39420 9367 39423
rect 9858 39420 9864 39432
rect 9355 39392 9864 39420
rect 9355 39389 9367 39392
rect 9309 39383 9367 39389
rect 9858 39380 9864 39392
rect 9916 39380 9922 39432
rect 12713 39423 12771 39429
rect 12713 39389 12725 39423
rect 12759 39389 12771 39423
rect 12713 39383 12771 39389
rect 6270 39352 6276 39364
rect 5184 39324 6276 39352
rect 6270 39312 6276 39324
rect 6328 39312 6334 39364
rect 9576 39355 9634 39361
rect 9576 39321 9588 39355
rect 9622 39352 9634 39355
rect 10042 39352 10048 39364
rect 9622 39324 10048 39352
rect 9622 39321 9634 39324
rect 9576 39315 9634 39321
rect 10042 39312 10048 39324
rect 10100 39312 10106 39364
rect 11146 39352 11152 39364
rect 11107 39324 11152 39352
rect 11146 39312 11152 39324
rect 11204 39312 11210 39364
rect 11330 39312 11336 39364
rect 11388 39352 11394 39364
rect 11974 39352 11980 39364
rect 11388 39324 11980 39352
rect 11388 39312 11394 39324
rect 11974 39312 11980 39324
rect 12032 39312 12038 39364
rect 12728 39296 12756 39383
rect 14550 39380 14556 39432
rect 14608 39414 14614 39432
rect 14691 39423 14749 39429
rect 14691 39414 14703 39423
rect 14608 39389 14703 39414
rect 14737 39420 14749 39423
rect 14829 39423 14887 39429
rect 14737 39389 14780 39420
rect 14608 39386 14780 39389
rect 14829 39389 14841 39423
rect 14875 39389 14887 39423
rect 14608 39380 14614 39386
rect 14691 39383 14749 39386
rect 14829 39383 14887 39389
rect 13630 39312 13636 39364
rect 13688 39352 13694 39364
rect 14844 39352 14872 39383
rect 14918 39380 14924 39432
rect 14976 39417 14982 39432
rect 15120 39429 15148 39460
rect 31404 39460 32321 39488
rect 15105 39423 15163 39429
rect 14976 39389 15018 39417
rect 15105 39389 15117 39423
rect 15151 39389 15163 39423
rect 14976 39380 14982 39389
rect 15105 39383 15163 39389
rect 16482 39380 16488 39432
rect 16540 39420 16546 39432
rect 18049 39423 18107 39429
rect 18049 39420 18061 39423
rect 16540 39392 18061 39420
rect 16540 39380 16546 39392
rect 18049 39389 18061 39392
rect 18095 39420 18107 39423
rect 18322 39420 18328 39432
rect 18095 39392 18328 39420
rect 18095 39389 18107 39392
rect 18049 39383 18107 39389
rect 18322 39380 18328 39392
rect 18380 39380 18386 39432
rect 19426 39380 19432 39432
rect 19484 39420 19490 39432
rect 20622 39420 20628 39432
rect 19484 39392 20628 39420
rect 19484 39380 19490 39392
rect 20622 39380 20628 39392
rect 20680 39380 20686 39432
rect 23842 39380 23848 39432
rect 23900 39420 23906 39432
rect 24394 39420 24400 39432
rect 23900 39392 24400 39420
rect 23900 39380 23906 39392
rect 24394 39380 24400 39392
rect 24452 39380 24458 39432
rect 27157 39423 27215 39429
rect 27157 39389 27169 39423
rect 27203 39420 27215 39423
rect 31113 39423 31171 39429
rect 27203 39392 27660 39420
rect 31113 39417 31125 39423
rect 27203 39389 27215 39392
rect 27157 39383 27215 39389
rect 27632 39364 27660 39392
rect 31036 39389 31125 39417
rect 31159 39389 31171 39423
rect 13688 39324 14872 39352
rect 15580 39324 17724 39352
rect 13688 39312 13694 39324
rect 5258 39284 5264 39296
rect 4080 39256 5264 39284
rect 5258 39244 5264 39256
rect 5316 39244 5322 39296
rect 7098 39244 7104 39296
rect 7156 39284 7162 39296
rect 7469 39287 7527 39293
rect 7469 39284 7481 39287
rect 7156 39256 7481 39284
rect 7156 39244 7162 39256
rect 7469 39253 7481 39256
rect 7515 39284 7527 39287
rect 8110 39284 8116 39296
rect 7515 39256 8116 39284
rect 7515 39253 7527 39256
rect 7469 39247 7527 39253
rect 8110 39244 8116 39256
rect 8168 39244 8174 39296
rect 10689 39287 10747 39293
rect 10689 39253 10701 39287
rect 10735 39284 10747 39287
rect 11238 39284 11244 39296
rect 10735 39256 11244 39284
rect 10735 39253 10747 39256
rect 10689 39247 10747 39253
rect 11238 39244 11244 39256
rect 11296 39244 11302 39296
rect 12253 39287 12311 39293
rect 12253 39253 12265 39287
rect 12299 39284 12311 39287
rect 12710 39284 12716 39296
rect 12299 39256 12716 39284
rect 12299 39253 12311 39256
rect 12253 39247 12311 39253
rect 12710 39244 12716 39256
rect 12768 39244 12774 39296
rect 14550 39244 14556 39296
rect 14608 39284 14614 39296
rect 15580 39293 15608 39324
rect 15565 39287 15623 39293
rect 15565 39284 15577 39287
rect 14608 39256 15577 39284
rect 14608 39244 14614 39256
rect 15565 39253 15577 39256
rect 15611 39253 15623 39287
rect 16666 39284 16672 39296
rect 16627 39256 16672 39284
rect 15565 39247 15623 39253
rect 16666 39244 16672 39256
rect 16724 39244 16730 39296
rect 17696 39284 17724 39324
rect 17770 39312 17776 39364
rect 17828 39361 17834 39364
rect 17828 39352 17840 39361
rect 20254 39352 20260 39364
rect 17828 39324 17873 39352
rect 18616 39324 20260 39352
rect 17828 39315 17840 39324
rect 17828 39312 17834 39315
rect 18616 39284 18644 39324
rect 20254 39312 20260 39324
rect 20312 39312 20318 39364
rect 20346 39312 20352 39364
rect 20404 39361 20410 39364
rect 20404 39352 20416 39361
rect 20404 39324 20449 39352
rect 20404 39315 20416 39324
rect 20404 39312 20410 39315
rect 23474 39312 23480 39364
rect 23532 39352 23538 39364
rect 24642 39355 24700 39361
rect 24642 39352 24654 39355
rect 23532 39324 24654 39352
rect 23532 39312 23538 39324
rect 24642 39321 24654 39324
rect 24688 39321 24700 39355
rect 24642 39315 24700 39321
rect 27246 39312 27252 39364
rect 27304 39352 27310 39364
rect 27402 39355 27460 39361
rect 27402 39352 27414 39355
rect 27304 39324 27414 39352
rect 27304 39312 27310 39324
rect 27402 39321 27414 39324
rect 27448 39321 27460 39355
rect 27402 39315 27460 39321
rect 27614 39312 27620 39364
rect 27672 39312 27678 39364
rect 31036 39352 31064 39389
rect 31113 39383 31171 39389
rect 31202 39420 31260 39426
rect 31202 39386 31214 39420
rect 31248 39386 31260 39420
rect 31202 39380 31260 39386
rect 31318 39423 31376 39429
rect 31318 39389 31330 39423
rect 31364 39420 31376 39423
rect 31404 39420 31432 39460
rect 32309 39457 32321 39460
rect 32355 39457 32367 39491
rect 32309 39451 32367 39457
rect 31364 39392 31432 39420
rect 31481 39423 31539 39429
rect 31364 39389 31376 39392
rect 31318 39383 31376 39389
rect 31481 39389 31493 39423
rect 31527 39420 31539 39423
rect 31570 39420 31576 39432
rect 31527 39392 31576 39420
rect 31527 39389 31539 39392
rect 31481 39383 31539 39389
rect 31570 39380 31576 39392
rect 31628 39380 31634 39432
rect 31217 39352 31245 39380
rect 30392 39324 31064 39352
rect 31128 39324 31245 39352
rect 31941 39355 31999 39361
rect 30392 39296 30420 39324
rect 31128 39296 31156 39324
rect 31941 39321 31953 39355
rect 31987 39321 31999 39355
rect 31941 39315 31999 39321
rect 17696 39256 18644 39284
rect 18693 39287 18751 39293
rect 18693 39253 18705 39287
rect 18739 39284 18751 39287
rect 20070 39284 20076 39296
rect 18739 39256 20076 39284
rect 18739 39253 18751 39256
rect 18693 39247 18751 39253
rect 20070 39244 20076 39256
rect 20128 39244 20134 39296
rect 24854 39244 24860 39296
rect 24912 39284 24918 39296
rect 25777 39287 25835 39293
rect 25777 39284 25789 39287
rect 24912 39256 25789 39284
rect 24912 39244 24918 39256
rect 25777 39253 25789 39256
rect 25823 39253 25835 39287
rect 25777 39247 25835 39253
rect 28537 39287 28595 39293
rect 28537 39253 28549 39287
rect 28583 39284 28595 39287
rect 28810 39284 28816 39296
rect 28583 39256 28816 39284
rect 28583 39253 28595 39256
rect 28537 39247 28595 39253
rect 28810 39244 28816 39256
rect 28868 39244 28874 39296
rect 28994 39244 29000 39296
rect 29052 39284 29058 39296
rect 29733 39287 29791 39293
rect 29733 39284 29745 39287
rect 29052 39256 29745 39284
rect 29052 39244 29058 39256
rect 29733 39253 29745 39256
rect 29779 39253 29791 39287
rect 30374 39284 30380 39296
rect 30335 39256 30380 39284
rect 29733 39247 29791 39253
rect 30374 39244 30380 39256
rect 30432 39244 30438 39296
rect 31110 39244 31116 39296
rect 31168 39244 31174 39296
rect 31478 39244 31484 39296
rect 31536 39284 31542 39296
rect 31956 39284 31984 39315
rect 32030 39312 32036 39364
rect 32088 39352 32094 39364
rect 32125 39355 32183 39361
rect 32125 39352 32137 39355
rect 32088 39324 32137 39352
rect 32088 39312 32094 39324
rect 32125 39321 32137 39324
rect 32171 39321 32183 39355
rect 32125 39315 32183 39321
rect 31536 39256 31984 39284
rect 31536 39244 31542 39256
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 6822 39040 6828 39092
rect 6880 39080 6886 39092
rect 6917 39083 6975 39089
rect 6917 39080 6929 39083
rect 6880 39052 6929 39080
rect 6880 39040 6886 39052
rect 6917 39049 6929 39052
rect 6963 39049 6975 39083
rect 6917 39043 6975 39049
rect 8386 39040 8392 39092
rect 8444 39080 8450 39092
rect 8444 39052 12434 39080
rect 8444 39040 8450 39052
rect 5442 39012 5448 39024
rect 4632 38984 5448 39012
rect 3533 38947 3591 38953
rect 3533 38913 3545 38947
rect 3579 38944 3591 38947
rect 4154 38944 4160 38956
rect 3579 38916 4160 38944
rect 3579 38913 3591 38916
rect 3533 38907 3591 38913
rect 4154 38904 4160 38916
rect 4212 38904 4218 38956
rect 4632 38888 4660 38984
rect 5442 38972 5448 38984
rect 5500 38972 5506 39024
rect 7098 39012 7104 39024
rect 7059 38984 7104 39012
rect 7098 38972 7104 38984
rect 7156 38972 7162 39024
rect 7208 38984 11744 39012
rect 4985 38947 5043 38953
rect 4985 38913 4997 38947
rect 5031 38944 5043 38947
rect 6457 38947 6515 38953
rect 6457 38944 6469 38947
rect 5031 38916 6469 38944
rect 5031 38913 5043 38916
rect 4985 38907 5043 38913
rect 6457 38913 6469 38916
rect 6503 38944 6515 38947
rect 7208 38944 7236 38984
rect 6503 38916 7236 38944
rect 7285 38947 7343 38953
rect 6503 38913 6515 38916
rect 6457 38907 6515 38913
rect 7285 38913 7297 38947
rect 7331 38913 7343 38947
rect 7285 38907 7343 38913
rect 9033 38947 9091 38953
rect 9033 38913 9045 38947
rect 9079 38944 9091 38947
rect 9079 38916 11652 38944
rect 9079 38913 9091 38916
rect 9033 38907 9091 38913
rect 3789 38879 3847 38885
rect 3789 38845 3801 38879
rect 3835 38876 3847 38879
rect 4614 38876 4620 38888
rect 3835 38848 4620 38876
rect 3835 38845 3847 38848
rect 3789 38839 3847 38845
rect 4614 38836 4620 38848
rect 4672 38836 4678 38888
rect 5074 38836 5080 38888
rect 5132 38876 5138 38888
rect 5261 38879 5319 38885
rect 5261 38876 5273 38879
rect 5132 38848 5273 38876
rect 5132 38836 5138 38848
rect 5261 38845 5273 38848
rect 5307 38845 5319 38879
rect 5261 38839 5319 38845
rect 6822 38836 6828 38888
rect 6880 38876 6886 38888
rect 7300 38876 7328 38907
rect 6880 38848 7328 38876
rect 6880 38836 6886 38848
rect 1946 38700 1952 38752
rect 2004 38740 2010 38752
rect 2409 38743 2467 38749
rect 2409 38740 2421 38743
rect 2004 38712 2421 38740
rect 2004 38700 2010 38712
rect 2409 38709 2421 38712
rect 2455 38709 2467 38743
rect 2409 38703 2467 38709
rect 3970 38700 3976 38752
rect 4028 38740 4034 38752
rect 4249 38743 4307 38749
rect 4249 38740 4261 38743
rect 4028 38712 4261 38740
rect 4028 38700 4034 38712
rect 4249 38709 4261 38712
rect 4295 38709 4307 38743
rect 4249 38703 4307 38709
rect 9858 38700 9864 38752
rect 9916 38740 9922 38752
rect 11624 38749 11652 38916
rect 11716 38808 11744 38984
rect 12406 38876 12434 39052
rect 13630 38904 13636 38956
rect 13688 38944 13694 38956
rect 13817 38947 13875 38953
rect 13817 38944 13829 38947
rect 13688 38916 13829 38944
rect 13688 38904 13694 38916
rect 13817 38913 13829 38916
rect 13863 38913 13875 38947
rect 13817 38907 13875 38913
rect 27893 38947 27951 38953
rect 27893 38913 27905 38947
rect 27939 38944 27951 38947
rect 28994 38944 29000 38956
rect 27939 38916 29000 38944
rect 27939 38913 27951 38916
rect 27893 38907 27951 38913
rect 28994 38904 29000 38916
rect 29052 38904 29058 38956
rect 30190 38904 30196 38956
rect 30248 38944 30254 38956
rect 30357 38947 30415 38953
rect 30357 38944 30369 38947
rect 30248 38916 30369 38944
rect 30248 38904 30254 38916
rect 30357 38913 30369 38916
rect 30403 38913 30415 38947
rect 30357 38907 30415 38913
rect 13541 38879 13599 38885
rect 13541 38876 13553 38879
rect 12406 38848 13553 38876
rect 13541 38845 13553 38848
rect 13587 38845 13599 38879
rect 30101 38879 30159 38885
rect 30101 38876 30113 38879
rect 13541 38839 13599 38845
rect 29196 38848 30113 38876
rect 12710 38808 12716 38820
rect 11716 38780 12716 38808
rect 12710 38768 12716 38780
rect 12768 38768 12774 38820
rect 10321 38743 10379 38749
rect 10321 38740 10333 38743
rect 9916 38712 10333 38740
rect 9916 38700 9922 38712
rect 10321 38709 10333 38712
rect 10367 38709 10379 38743
rect 10321 38703 10379 38709
rect 11609 38743 11667 38749
rect 11609 38709 11621 38743
rect 11655 38740 11667 38743
rect 11790 38740 11796 38752
rect 11655 38712 11796 38740
rect 11655 38709 11667 38712
rect 11609 38703 11667 38709
rect 11790 38700 11796 38712
rect 11848 38700 11854 38752
rect 23382 38700 23388 38752
rect 23440 38740 23446 38752
rect 26970 38740 26976 38752
rect 23440 38712 26976 38740
rect 23440 38700 23446 38712
rect 26970 38700 26976 38712
rect 27028 38700 27034 38752
rect 27614 38700 27620 38752
rect 27672 38740 27678 38752
rect 29196 38749 29224 38848
rect 30101 38845 30113 38848
rect 30147 38845 30159 38879
rect 30101 38839 30159 38845
rect 58158 38808 58164 38820
rect 58119 38780 58164 38808
rect 58158 38768 58164 38780
rect 58216 38768 58222 38820
rect 29181 38743 29239 38749
rect 29181 38740 29193 38743
rect 27672 38712 29193 38740
rect 27672 38700 27678 38712
rect 29181 38709 29193 38712
rect 29227 38709 29239 38743
rect 29181 38703 29239 38709
rect 29730 38700 29736 38752
rect 29788 38740 29794 38752
rect 31481 38743 31539 38749
rect 31481 38740 31493 38743
rect 29788 38712 31493 38740
rect 29788 38700 29794 38712
rect 31481 38709 31493 38712
rect 31527 38709 31539 38743
rect 31481 38703 31539 38709
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 4798 38536 4804 38548
rect 2148 38508 4804 38536
rect 2148 38341 2176 38508
rect 4798 38496 4804 38508
rect 4856 38496 4862 38548
rect 6270 38496 6276 38548
rect 6328 38536 6334 38548
rect 6365 38539 6423 38545
rect 6365 38536 6377 38539
rect 6328 38508 6377 38536
rect 6328 38496 6334 38508
rect 6365 38505 6377 38508
rect 6411 38505 6423 38539
rect 10042 38536 10048 38548
rect 10003 38508 10048 38536
rect 6365 38499 6423 38505
rect 10042 38496 10048 38508
rect 10100 38496 10106 38548
rect 12529 38539 12587 38545
rect 12529 38505 12541 38539
rect 12575 38536 12587 38539
rect 14274 38536 14280 38548
rect 12575 38508 14280 38536
rect 12575 38505 12587 38508
rect 12529 38499 12587 38505
rect 14274 38496 14280 38508
rect 14332 38496 14338 38548
rect 23382 38536 23388 38548
rect 18156 38508 23388 38536
rect 18156 38480 18184 38508
rect 23382 38496 23388 38508
rect 23440 38496 23446 38548
rect 27246 38536 27252 38548
rect 27207 38508 27252 38536
rect 27246 38496 27252 38508
rect 27304 38496 27310 38548
rect 28350 38536 28356 38548
rect 28311 38508 28356 38536
rect 28350 38496 28356 38508
rect 28408 38496 28414 38548
rect 9585 38471 9643 38477
rect 9585 38437 9597 38471
rect 9631 38468 9643 38471
rect 9674 38468 9680 38480
rect 9631 38440 9680 38468
rect 9631 38437 9643 38440
rect 9585 38431 9643 38437
rect 9674 38428 9680 38440
rect 9732 38428 9738 38480
rect 10410 38428 10416 38480
rect 10468 38428 10474 38480
rect 12618 38428 12624 38480
rect 12676 38468 12682 38480
rect 18138 38468 18144 38480
rect 12676 38440 18144 38468
rect 12676 38428 12682 38440
rect 18138 38428 18144 38440
rect 18196 38428 18202 38480
rect 3970 38400 3976 38412
rect 2884 38372 3976 38400
rect 2884 38344 2912 38372
rect 3970 38360 3976 38372
rect 4028 38360 4034 38412
rect 4430 38360 4436 38412
rect 4488 38400 4494 38412
rect 5350 38400 5356 38412
rect 4488 38372 5356 38400
rect 4488 38360 4494 38372
rect 5350 38360 5356 38372
rect 5408 38400 5414 38412
rect 8113 38403 8171 38409
rect 8113 38400 8125 38403
rect 5408 38372 8125 38400
rect 5408 38360 5414 38372
rect 8113 38369 8125 38372
rect 8159 38369 8171 38403
rect 8113 38363 8171 38369
rect 2133 38335 2191 38341
rect 2133 38301 2145 38335
rect 2179 38301 2191 38335
rect 2866 38332 2872 38344
rect 2779 38304 2872 38332
rect 2133 38295 2191 38301
rect 2866 38292 2872 38304
rect 2924 38292 2930 38344
rect 2961 38335 3019 38341
rect 2961 38301 2973 38335
rect 3007 38301 3019 38335
rect 2961 38295 3019 38301
rect 3053 38335 3111 38341
rect 3053 38301 3065 38335
rect 3099 38301 3111 38335
rect 3053 38295 3111 38301
rect 3237 38335 3295 38341
rect 3237 38301 3249 38335
rect 3283 38332 3295 38335
rect 5074 38332 5080 38344
rect 3283 38304 5080 38332
rect 3283 38301 3295 38304
rect 3237 38295 3295 38301
rect 1946 38264 1952 38276
rect 1907 38236 1952 38264
rect 1946 38224 1952 38236
rect 2004 38224 2010 38276
rect 1762 38196 1768 38208
rect 1723 38168 1768 38196
rect 1762 38156 1768 38168
rect 1820 38156 1826 38208
rect 2593 38199 2651 38205
rect 2593 38165 2605 38199
rect 2639 38196 2651 38199
rect 2682 38196 2688 38208
rect 2639 38168 2688 38196
rect 2639 38165 2651 38168
rect 2593 38159 2651 38165
rect 2682 38156 2688 38168
rect 2740 38156 2746 38208
rect 2976 38196 3004 38295
rect 3068 38264 3096 38295
rect 5074 38292 5080 38304
rect 5132 38292 5138 38344
rect 6546 38332 6552 38344
rect 6507 38304 6552 38332
rect 6546 38292 6552 38304
rect 6604 38292 6610 38344
rect 8386 38332 8392 38344
rect 8347 38304 8392 38332
rect 8386 38292 8392 38304
rect 8444 38292 8450 38344
rect 8846 38292 8852 38344
rect 8904 38332 8910 38344
rect 9398 38332 9404 38344
rect 8904 38304 9404 38332
rect 8904 38292 8910 38304
rect 9398 38292 9404 38304
rect 9456 38292 9462 38344
rect 10226 38292 10232 38344
rect 10284 38341 10290 38344
rect 10425 38341 10453 38428
rect 11149 38403 11207 38409
rect 11149 38400 11161 38403
rect 10284 38335 10333 38341
rect 10284 38301 10287 38335
rect 10321 38301 10333 38335
rect 10284 38295 10333 38301
rect 10394 38335 10453 38341
rect 10541 38372 11161 38400
rect 10541 38338 10569 38372
rect 11149 38369 11161 38372
rect 11195 38369 11207 38403
rect 20622 38400 20628 38412
rect 11149 38363 11207 38369
rect 11348 38372 13032 38400
rect 20583 38372 20628 38400
rect 10394 38301 10406 38335
rect 10440 38304 10453 38335
rect 10526 38332 10584 38338
rect 10440 38301 10452 38304
rect 10394 38295 10452 38301
rect 10526 38298 10538 38332
rect 10572 38298 10584 38332
rect 10284 38292 10290 38295
rect 10526 38292 10584 38298
rect 10701 38335 10759 38341
rect 10701 38301 10713 38335
rect 10747 38332 10759 38335
rect 10962 38332 10968 38344
rect 10747 38304 10968 38332
rect 10747 38301 10759 38304
rect 10701 38295 10759 38301
rect 10962 38292 10968 38304
rect 11020 38292 11026 38344
rect 11238 38292 11244 38344
rect 11296 38332 11302 38344
rect 11348 38341 11376 38372
rect 11333 38335 11391 38341
rect 11333 38332 11345 38335
rect 11296 38304 11345 38332
rect 11296 38292 11302 38304
rect 11333 38301 11345 38304
rect 11379 38301 11391 38335
rect 11333 38295 11391 38301
rect 12345 38335 12403 38341
rect 12345 38301 12357 38335
rect 12391 38332 12403 38335
rect 12618 38332 12624 38344
rect 12391 38304 12624 38332
rect 12391 38301 12403 38304
rect 12345 38295 12403 38301
rect 12618 38292 12624 38304
rect 12676 38292 12682 38344
rect 13004 38341 13032 38372
rect 20622 38360 20628 38372
rect 20680 38360 20686 38412
rect 31110 38400 31116 38412
rect 27632 38372 31116 38400
rect 12989 38335 13047 38341
rect 12989 38301 13001 38335
rect 13035 38301 13047 38335
rect 13354 38332 13360 38344
rect 13315 38304 13360 38332
rect 12989 38295 13047 38301
rect 13354 38292 13360 38304
rect 13412 38292 13418 38344
rect 27632 38341 27660 38372
rect 27525 38335 27583 38341
rect 27525 38332 27537 38335
rect 27080 38304 27537 38332
rect 5350 38264 5356 38276
rect 3068 38236 5356 38264
rect 5350 38224 5356 38236
rect 5408 38224 5414 38276
rect 5902 38264 5908 38276
rect 5863 38236 5908 38264
rect 5902 38224 5908 38236
rect 5960 38224 5966 38276
rect 6730 38264 6736 38276
rect 6691 38236 6736 38264
rect 6730 38224 6736 38236
rect 6788 38224 6794 38276
rect 9217 38267 9275 38273
rect 9217 38233 9229 38267
rect 9263 38233 9275 38267
rect 9217 38227 9275 38233
rect 4430 38196 4436 38208
rect 2976 38168 4436 38196
rect 4430 38156 4436 38168
rect 4488 38156 4494 38208
rect 4614 38196 4620 38208
rect 4575 38168 4620 38196
rect 4614 38156 4620 38168
rect 4672 38156 4678 38208
rect 9232 38196 9260 38227
rect 11146 38224 11152 38276
rect 11204 38264 11210 38276
rect 11514 38264 11520 38276
rect 11204 38236 11520 38264
rect 11204 38224 11210 38236
rect 11514 38224 11520 38236
rect 11572 38224 11578 38276
rect 13170 38264 13176 38276
rect 13131 38236 13176 38264
rect 13170 38224 13176 38236
rect 13228 38224 13234 38276
rect 13265 38267 13323 38273
rect 13265 38233 13277 38267
rect 13311 38264 13323 38267
rect 16666 38264 16672 38276
rect 13311 38236 16672 38264
rect 13311 38233 13323 38236
rect 13265 38227 13323 38233
rect 16666 38224 16672 38236
rect 16724 38224 16730 38276
rect 19426 38224 19432 38276
rect 19484 38264 19490 38276
rect 20358 38267 20416 38273
rect 20358 38264 20370 38267
rect 19484 38236 20370 38264
rect 19484 38224 19490 38236
rect 20358 38233 20370 38236
rect 20404 38233 20416 38267
rect 20358 38227 20416 38233
rect 9490 38196 9496 38208
rect 9232 38168 9496 38196
rect 9490 38156 9496 38168
rect 9548 38196 9554 38208
rect 11164 38196 11192 38224
rect 27080 38208 27108 38304
rect 27525 38301 27537 38304
rect 27571 38301 27583 38335
rect 27525 38295 27583 38301
rect 27617 38335 27675 38341
rect 27617 38301 27629 38335
rect 27663 38301 27675 38335
rect 27617 38295 27675 38301
rect 27706 38292 27712 38344
rect 27764 38332 27770 38344
rect 27893 38335 27951 38341
rect 27764 38304 27809 38332
rect 27764 38292 27770 38304
rect 27893 38301 27905 38335
rect 27939 38301 27951 38335
rect 27893 38295 27951 38301
rect 27908 38264 27936 38295
rect 27982 38292 27988 38344
rect 28040 38332 28046 38344
rect 28736 38341 28764 38372
rect 31110 38360 31116 38372
rect 31168 38360 31174 38412
rect 32214 38400 32220 38412
rect 32175 38372 32220 38400
rect 32214 38360 32220 38372
rect 32272 38400 32278 38412
rect 32674 38400 32680 38412
rect 32272 38372 32680 38400
rect 32272 38360 32278 38372
rect 32674 38360 32680 38372
rect 32732 38360 32738 38412
rect 28629 38335 28687 38341
rect 28629 38332 28641 38335
rect 28040 38304 28641 38332
rect 28040 38292 28046 38304
rect 28629 38301 28641 38304
rect 28675 38301 28687 38335
rect 28629 38295 28687 38301
rect 28721 38335 28779 38341
rect 28721 38301 28733 38335
rect 28767 38301 28779 38335
rect 28721 38295 28779 38301
rect 28813 38335 28871 38341
rect 28813 38301 28825 38335
rect 28859 38332 28871 38335
rect 28902 38332 28908 38344
rect 28859 38304 28908 38332
rect 28859 38301 28871 38304
rect 28813 38295 28871 38301
rect 28902 38292 28908 38304
rect 28960 38292 28966 38344
rect 28997 38335 29055 38341
rect 28997 38301 29009 38335
rect 29043 38301 29055 38335
rect 28997 38295 29055 38301
rect 29012 38264 29040 38295
rect 29270 38292 29276 38344
rect 29328 38332 29334 38344
rect 30009 38335 30067 38341
rect 30009 38332 30021 38335
rect 29328 38304 30021 38332
rect 29328 38292 29334 38304
rect 30009 38301 30021 38304
rect 30055 38332 30067 38335
rect 30742 38332 30748 38344
rect 30055 38304 30748 38332
rect 30055 38301 30067 38304
rect 30009 38295 30067 38301
rect 30742 38292 30748 38304
rect 30800 38332 30806 38344
rect 31478 38332 31484 38344
rect 30800 38304 31484 38332
rect 30800 38292 30806 38304
rect 31478 38292 31484 38304
rect 31536 38292 31542 38344
rect 30098 38264 30104 38276
rect 27908 38236 30104 38264
rect 30098 38224 30104 38236
rect 30156 38224 30162 38276
rect 30193 38267 30251 38273
rect 30193 38233 30205 38267
rect 30239 38264 30251 38267
rect 30239 38236 30880 38264
rect 30239 38233 30251 38236
rect 30193 38227 30251 38233
rect 9548 38168 11192 38196
rect 13541 38199 13599 38205
rect 9548 38156 9554 38168
rect 13541 38165 13553 38199
rect 13587 38196 13599 38199
rect 17126 38196 17132 38208
rect 13587 38168 17132 38196
rect 13587 38165 13599 38168
rect 13541 38159 13599 38165
rect 17126 38156 17132 38168
rect 17184 38156 17190 38208
rect 19058 38156 19064 38208
rect 19116 38196 19122 38208
rect 19245 38199 19303 38205
rect 19245 38196 19257 38199
rect 19116 38168 19257 38196
rect 19116 38156 19122 38168
rect 19245 38165 19257 38168
rect 19291 38165 19303 38199
rect 19245 38159 19303 38165
rect 26789 38199 26847 38205
rect 26789 38165 26801 38199
rect 26835 38196 26847 38199
rect 27062 38196 27068 38208
rect 26835 38168 27068 38196
rect 26835 38165 26847 38168
rect 26789 38159 26847 38165
rect 27062 38156 27068 38168
rect 27120 38156 27126 38208
rect 30377 38199 30435 38205
rect 30377 38165 30389 38199
rect 30423 38196 30435 38199
rect 30466 38196 30472 38208
rect 30423 38168 30472 38196
rect 30423 38165 30435 38168
rect 30377 38159 30435 38165
rect 30466 38156 30472 38168
rect 30524 38156 30530 38208
rect 30852 38205 30880 38236
rect 31018 38224 31024 38276
rect 31076 38264 31082 38276
rect 31950 38267 32008 38273
rect 31950 38264 31962 38267
rect 31076 38236 31962 38264
rect 31076 38224 31082 38236
rect 31950 38233 31962 38236
rect 31996 38233 32008 38267
rect 31950 38227 32008 38233
rect 32944 38267 33002 38273
rect 32944 38233 32956 38267
rect 32990 38264 33002 38267
rect 33042 38264 33048 38276
rect 32990 38236 33048 38264
rect 32990 38233 33002 38236
rect 32944 38227 33002 38233
rect 33042 38224 33048 38236
rect 33100 38224 33106 38276
rect 30837 38199 30895 38205
rect 30837 38165 30849 38199
rect 30883 38196 30895 38199
rect 31386 38196 31392 38208
rect 30883 38168 31392 38196
rect 30883 38165 30895 38168
rect 30837 38159 30895 38165
rect 31386 38156 31392 38168
rect 31444 38156 31450 38208
rect 33870 38156 33876 38208
rect 33928 38196 33934 38208
rect 34057 38199 34115 38205
rect 34057 38196 34069 38199
rect 33928 38168 34069 38196
rect 33928 38156 33934 38168
rect 34057 38165 34069 38168
rect 34103 38165 34115 38199
rect 34057 38159 34115 38165
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 4154 37952 4160 38004
rect 4212 37992 4218 38004
rect 4249 37995 4307 38001
rect 4249 37992 4261 37995
rect 4212 37964 4261 37992
rect 4212 37952 4218 37964
rect 4249 37961 4261 37964
rect 4295 37961 4307 37995
rect 5350 37992 5356 38004
rect 5311 37964 5356 37992
rect 4249 37955 4307 37961
rect 5350 37952 5356 37964
rect 5408 37952 5414 38004
rect 6730 37992 6736 38004
rect 5736 37964 6736 37992
rect 1762 37884 1768 37936
rect 1820 37924 1826 37936
rect 1820 37896 4752 37924
rect 1820 37884 1826 37896
rect 2409 37859 2467 37865
rect 2409 37825 2421 37859
rect 2455 37856 2467 37859
rect 2498 37856 2504 37868
rect 2455 37828 2504 37856
rect 2455 37825 2467 37828
rect 2409 37819 2467 37825
rect 2498 37816 2504 37828
rect 2556 37816 2562 37868
rect 2682 37865 2688 37868
rect 2676 37856 2688 37865
rect 2643 37828 2688 37856
rect 2676 37819 2688 37828
rect 2682 37816 2688 37819
rect 2740 37816 2746 37868
rect 4724 37865 4752 37896
rect 4798 37884 4804 37936
rect 4856 37924 4862 37936
rect 5736 37933 5764 37964
rect 6730 37952 6736 37964
rect 6788 37992 6794 38004
rect 9125 37995 9183 38001
rect 9125 37992 9137 37995
rect 6788 37964 9137 37992
rect 6788 37952 6794 37964
rect 9125 37961 9137 37964
rect 9171 37961 9183 37995
rect 9125 37955 9183 37961
rect 10226 37952 10232 38004
rect 10284 37992 10290 38004
rect 10778 37992 10784 38004
rect 10284 37964 10784 37992
rect 10284 37952 10290 37964
rect 10778 37952 10784 37964
rect 10836 37952 10842 38004
rect 13170 37992 13176 38004
rect 11716 37964 13176 37992
rect 5721 37927 5779 37933
rect 5721 37924 5733 37927
rect 4856 37896 5733 37924
rect 4856 37884 4862 37896
rect 5721 37893 5733 37896
rect 5767 37893 5779 37927
rect 5721 37887 5779 37893
rect 4525 37859 4583 37865
rect 4525 37856 4537 37859
rect 4356 37828 4537 37856
rect 4356 37720 4384 37828
rect 4525 37825 4537 37828
rect 4571 37825 4583 37859
rect 4525 37819 4583 37825
rect 4617 37859 4675 37865
rect 4617 37825 4629 37859
rect 4663 37825 4675 37859
rect 4617 37819 4675 37825
rect 4709 37859 4767 37865
rect 4709 37825 4721 37859
rect 4755 37825 4767 37859
rect 4709 37819 4767 37825
rect 4893 37859 4951 37865
rect 4893 37825 4905 37859
rect 4939 37856 4951 37859
rect 5074 37856 5080 37868
rect 4939 37828 5080 37856
rect 4939 37825 4951 37828
rect 4893 37819 4951 37825
rect 4430 37748 4436 37800
rect 4488 37788 4494 37800
rect 4632 37788 4660 37819
rect 5074 37816 5080 37828
rect 5132 37816 5138 37868
rect 5537 37859 5595 37865
rect 5537 37825 5549 37859
rect 5583 37825 5595 37859
rect 5537 37819 5595 37825
rect 9309 37859 9367 37865
rect 9309 37825 9321 37859
rect 9355 37825 9367 37859
rect 9309 37819 9367 37825
rect 4488 37760 4660 37788
rect 4488 37748 4494 37760
rect 4798 37748 4804 37800
rect 4856 37788 4862 37800
rect 5552 37788 5580 37819
rect 4856 37760 5580 37788
rect 9324 37788 9352 37819
rect 9398 37816 9404 37868
rect 9456 37856 9462 37868
rect 11517 37859 11575 37865
rect 11517 37856 11529 37859
rect 9456 37828 11529 37856
rect 9456 37816 9462 37828
rect 11517 37825 11529 37828
rect 11563 37825 11575 37859
rect 11517 37819 11575 37825
rect 11606 37816 11612 37868
rect 11664 37856 11670 37868
rect 11716 37865 11744 37964
rect 13170 37952 13176 37964
rect 13228 37992 13234 38004
rect 13725 37995 13783 38001
rect 13228 37964 13400 37992
rect 13228 37952 13234 37964
rect 11793 37927 11851 37933
rect 11793 37893 11805 37927
rect 11839 37924 11851 37927
rect 12158 37924 12164 37936
rect 11839 37896 12164 37924
rect 11839 37893 11851 37896
rect 11793 37887 11851 37893
rect 12158 37884 12164 37896
rect 12216 37884 12222 37936
rect 13372 37933 13400 37964
rect 13725 37961 13737 37995
rect 13771 37961 13783 37995
rect 13725 37955 13783 37961
rect 13357 37927 13415 37933
rect 13357 37893 13369 37927
rect 13403 37893 13415 37927
rect 13357 37887 13415 37893
rect 13449 37927 13507 37933
rect 13449 37893 13461 37927
rect 13495 37924 13507 37927
rect 13740 37924 13768 37955
rect 18322 37952 18328 38004
rect 18380 37992 18386 38004
rect 18380 37964 19196 37992
rect 18380 37952 18386 37964
rect 19168 37933 19196 37964
rect 19334 37952 19340 38004
rect 19392 37952 19398 38004
rect 27706 37952 27712 38004
rect 27764 37992 27770 38004
rect 28077 37995 28135 38001
rect 28077 37992 28089 37995
rect 27764 37964 28089 37992
rect 27764 37952 27770 37964
rect 28077 37961 28089 37964
rect 28123 37961 28135 37995
rect 28902 37992 28908 38004
rect 28863 37964 28908 37992
rect 28077 37955 28135 37961
rect 28902 37952 28908 37964
rect 28960 37952 28966 38004
rect 29822 37952 29828 38004
rect 29880 37992 29886 38004
rect 29917 37995 29975 38001
rect 29917 37992 29929 37995
rect 29880 37964 29929 37992
rect 29880 37952 29886 37964
rect 29917 37961 29929 37964
rect 29963 37992 29975 37995
rect 31018 37992 31024 38004
rect 29963 37964 30880 37992
rect 30979 37964 31024 37992
rect 29963 37961 29975 37964
rect 29917 37955 29975 37961
rect 19153 37927 19211 37933
rect 13495 37896 13676 37924
rect 13740 37896 18920 37924
rect 13495 37893 13507 37896
rect 13449 37887 13507 37893
rect 11701 37859 11759 37865
rect 11701 37856 11713 37859
rect 11664 37828 11713 37856
rect 11664 37816 11670 37828
rect 11701 37825 11713 37828
rect 11747 37825 11759 37859
rect 11882 37856 11888 37868
rect 11843 37828 11888 37856
rect 11701 37819 11759 37825
rect 11882 37816 11888 37828
rect 11940 37816 11946 37868
rect 11974 37816 11980 37868
rect 12032 37856 12038 37868
rect 13173 37859 13231 37865
rect 13173 37856 13185 37859
rect 12032 37828 13185 37856
rect 12032 37816 12038 37828
rect 13173 37825 13185 37828
rect 13219 37825 13231 37859
rect 13173 37819 13231 37825
rect 13262 37816 13268 37868
rect 13320 37856 13326 37868
rect 13541 37859 13599 37865
rect 13541 37856 13553 37859
rect 13320 37828 13553 37856
rect 13320 37816 13326 37828
rect 13541 37825 13553 37828
rect 13587 37825 13599 37859
rect 13648 37856 13676 37896
rect 16022 37856 16028 37868
rect 13648 37828 16028 37856
rect 13541 37819 13599 37825
rect 16022 37816 16028 37828
rect 16080 37816 16086 37868
rect 17126 37856 17132 37868
rect 17087 37828 17132 37856
rect 17126 37816 17132 37828
rect 17184 37816 17190 37868
rect 17222 37859 17280 37865
rect 17222 37825 17234 37859
rect 17268 37825 17280 37859
rect 17222 37819 17280 37825
rect 17405 37859 17463 37865
rect 17405 37825 17417 37859
rect 17451 37825 17463 37859
rect 17405 37819 17463 37825
rect 12618 37788 12624 37800
rect 9324 37760 12624 37788
rect 4856 37748 4862 37760
rect 12618 37748 12624 37760
rect 12676 37748 12682 37800
rect 17034 37748 17040 37800
rect 17092 37788 17098 37800
rect 17236 37788 17264 37819
rect 17092 37760 17264 37788
rect 17420 37788 17448 37819
rect 17494 37816 17500 37868
rect 17552 37856 17558 37868
rect 17635 37859 17693 37865
rect 17552 37828 17597 37856
rect 17552 37816 17558 37828
rect 17635 37825 17647 37859
rect 17681 37856 17693 37859
rect 18506 37856 18512 37868
rect 17681 37828 18512 37856
rect 17681 37825 17693 37828
rect 17635 37819 17693 37825
rect 18506 37816 18512 37828
rect 18564 37816 18570 37868
rect 18892 37865 18920 37896
rect 19153 37893 19165 37927
rect 19199 37893 19211 37927
rect 19153 37887 19211 37893
rect 19245 37927 19303 37933
rect 19245 37893 19257 37927
rect 19291 37924 19303 37927
rect 19352 37924 19380 37952
rect 20070 37924 20076 37936
rect 19291 37896 19380 37924
rect 19996 37896 20076 37924
rect 19291 37893 19303 37896
rect 19245 37887 19303 37893
rect 19058 37865 19064 37868
rect 18877 37859 18935 37865
rect 18877 37825 18889 37859
rect 18923 37825 18935 37859
rect 18877 37819 18935 37825
rect 19025 37859 19064 37865
rect 19025 37825 19037 37859
rect 19025 37819 19064 37825
rect 19058 37816 19064 37819
rect 19116 37816 19122 37868
rect 19996 37865 20024 37896
rect 20070 37884 20076 37896
rect 20128 37884 20134 37936
rect 20438 37924 20444 37936
rect 20272 37896 20444 37924
rect 19342 37859 19400 37865
rect 19342 37856 19354 37859
rect 19260 37828 19354 37856
rect 18322 37788 18328 37800
rect 17420 37760 18328 37788
rect 17092 37748 17098 37760
rect 18322 37748 18328 37760
rect 18380 37748 18386 37800
rect 18524 37788 18552 37816
rect 19260 37788 19288 37828
rect 19342 37825 19354 37828
rect 19388 37825 19400 37859
rect 19342 37819 19400 37825
rect 19981 37859 20039 37865
rect 19981 37825 19993 37859
rect 20027 37825 20039 37859
rect 20162 37856 20168 37868
rect 20123 37828 20168 37856
rect 19981 37819 20039 37825
rect 20162 37816 20168 37828
rect 20220 37816 20226 37868
rect 20272 37865 20300 37896
rect 20438 37884 20444 37896
rect 20496 37884 20502 37936
rect 26053 37927 26111 37933
rect 26053 37924 26065 37927
rect 22066 37896 26065 37924
rect 20257 37859 20315 37865
rect 20257 37825 20269 37859
rect 20303 37825 20315 37859
rect 20257 37819 20315 37825
rect 20349 37859 20407 37865
rect 20349 37825 20361 37859
rect 20395 37856 20407 37859
rect 21085 37859 21143 37865
rect 21085 37856 21097 37859
rect 20395 37828 21097 37856
rect 20395 37825 20407 37828
rect 20349 37819 20407 37825
rect 21085 37825 21097 37828
rect 21131 37856 21143 37859
rect 22066 37856 22094 37896
rect 26053 37893 26065 37896
rect 26099 37924 26111 37927
rect 26510 37924 26516 37936
rect 26099 37896 26516 37924
rect 26099 37893 26111 37896
rect 26053 37887 26111 37893
rect 26510 37884 26516 37896
rect 26568 37884 26574 37936
rect 28261 37927 28319 37933
rect 28261 37893 28273 37927
rect 28307 37924 28319 37927
rect 28810 37924 28816 37936
rect 28307 37896 28816 37924
rect 28307 37893 28319 37896
rect 28261 37887 28319 37893
rect 28810 37884 28816 37896
rect 28868 37884 28874 37936
rect 29270 37924 29276 37936
rect 29012 37896 29276 37924
rect 21131 37828 22094 37856
rect 24213 37859 24271 37865
rect 21131 37825 21143 37828
rect 21085 37819 21143 37825
rect 24213 37825 24225 37859
rect 24259 37856 24271 37859
rect 24302 37856 24308 37868
rect 24259 37828 24308 37856
rect 24259 37825 24271 37828
rect 24213 37819 24271 37825
rect 20364 37788 20392 37819
rect 24302 37816 24308 37828
rect 24360 37816 24366 37868
rect 24480 37859 24538 37865
rect 24480 37825 24492 37859
rect 24526 37856 24538 37859
rect 26234 37856 26240 37868
rect 24526 37828 26240 37856
rect 24526 37825 24538 37828
rect 24480 37819 24538 37825
rect 26234 37816 26240 37828
rect 26292 37816 26298 37868
rect 28445 37859 28503 37865
rect 28445 37825 28457 37859
rect 28491 37856 28503 37859
rect 29012 37856 29040 37896
rect 29270 37884 29276 37896
rect 29328 37884 29334 37936
rect 30466 37924 30472 37936
rect 30463 37884 30472 37924
rect 30524 37884 30530 37936
rect 28491 37828 29040 37856
rect 29089 37859 29147 37865
rect 28491 37825 28503 37828
rect 28445 37819 28503 37825
rect 29089 37825 29101 37859
rect 29135 37856 29147 37859
rect 29178 37856 29184 37868
rect 29135 37828 29184 37856
rect 29135 37825 29147 37828
rect 29089 37819 29147 37825
rect 29178 37816 29184 37828
rect 29236 37816 29242 37868
rect 30098 37816 30104 37868
rect 30156 37856 30162 37868
rect 30377 37859 30435 37865
rect 30377 37856 30389 37859
rect 30156 37828 30389 37856
rect 30156 37816 30162 37828
rect 30377 37825 30389 37828
rect 30423 37825 30435 37859
rect 30463 37856 30491 37884
rect 30556 37859 30614 37865
rect 30556 37856 30568 37859
rect 30463 37828 30568 37856
rect 30377 37819 30435 37825
rect 30556 37825 30568 37828
rect 30602 37825 30614 37859
rect 30556 37819 30614 37825
rect 30653 37862 30711 37868
rect 30765 37862 30823 37865
rect 30852 37862 30880 37964
rect 31018 37952 31024 37964
rect 31076 37952 31082 38004
rect 33042 37992 33048 38004
rect 33003 37964 33048 37992
rect 33042 37952 33048 37964
rect 33100 37952 33106 38004
rect 34606 37992 34612 38004
rect 33152 37964 34612 37992
rect 33152 37924 33180 37964
rect 32692 37896 33180 37924
rect 34532 37924 34560 37964
rect 34606 37952 34612 37964
rect 34664 37952 34670 38004
rect 34532 37896 34652 37924
rect 30653 37828 30665 37862
rect 30699 37828 30711 37862
rect 30760 37859 30880 37862
rect 30760 37828 30777 37859
rect 30653 37822 30711 37828
rect 30765 37825 30777 37828
rect 30811 37834 30880 37859
rect 30811 37825 30823 37834
rect 18524 37760 19288 37788
rect 19444 37760 20392 37788
rect 30668 37788 30696 37822
rect 30765 37819 30823 37825
rect 31294 37816 31300 37868
rect 31352 37856 31358 37868
rect 31570 37856 31576 37868
rect 31352 37828 31576 37856
rect 31352 37816 31358 37828
rect 31570 37816 31576 37828
rect 31628 37856 31634 37868
rect 32401 37859 32459 37865
rect 32401 37856 32413 37859
rect 31628 37828 32413 37856
rect 31628 37816 31634 37828
rect 32401 37825 32413 37828
rect 32447 37825 32459 37859
rect 32582 37856 32588 37868
rect 32543 37828 32588 37856
rect 32401 37819 32459 37825
rect 32582 37816 32588 37828
rect 32640 37816 32646 37868
rect 32692 37865 32720 37896
rect 32677 37859 32735 37865
rect 32677 37825 32689 37859
rect 32723 37825 32735 37859
rect 32677 37819 32735 37825
rect 32769 37859 32827 37865
rect 32769 37825 32781 37859
rect 32815 37825 32827 37859
rect 32769 37819 32827 37825
rect 31018 37788 31024 37800
rect 30668 37760 31024 37788
rect 5718 37720 5724 37732
rect 4356 37692 5724 37720
rect 5718 37680 5724 37692
rect 5776 37680 5782 37732
rect 5902 37680 5908 37732
rect 5960 37720 5966 37732
rect 6457 37723 6515 37729
rect 6457 37720 6469 37723
rect 5960 37692 6469 37720
rect 5960 37680 5966 37692
rect 6457 37689 6469 37692
rect 6503 37720 6515 37723
rect 11790 37720 11796 37732
rect 6503 37692 11796 37720
rect 6503 37689 6515 37692
rect 6457 37683 6515 37689
rect 11790 37680 11796 37692
rect 11848 37680 11854 37732
rect 11900 37692 13860 37720
rect 3789 37655 3847 37661
rect 3789 37621 3801 37655
rect 3835 37652 3847 37655
rect 4706 37652 4712 37664
rect 3835 37624 4712 37652
rect 3835 37621 3847 37624
rect 3789 37615 3847 37621
rect 4706 37612 4712 37624
rect 4764 37612 4770 37664
rect 10778 37612 10784 37664
rect 10836 37652 10842 37664
rect 11900 37652 11928 37692
rect 10836 37624 11928 37652
rect 12069 37655 12127 37661
rect 10836 37612 10842 37624
rect 12069 37621 12081 37655
rect 12115 37652 12127 37655
rect 13630 37652 13636 37664
rect 12115 37624 13636 37652
rect 12115 37621 12127 37624
rect 12069 37615 12127 37621
rect 13630 37612 13636 37624
rect 13688 37612 13694 37664
rect 13832 37652 13860 37692
rect 13906 37680 13912 37732
rect 13964 37720 13970 37732
rect 19444 37720 19472 37760
rect 31018 37748 31024 37760
rect 31076 37748 31082 37800
rect 32784 37788 32812 37819
rect 34238 37816 34244 37868
rect 34296 37856 34302 37868
rect 34333 37859 34391 37865
rect 34333 37856 34345 37859
rect 34296 37828 34345 37856
rect 34296 37816 34302 37828
rect 34333 37825 34345 37828
rect 34379 37825 34391 37859
rect 34514 37856 34520 37868
rect 34475 37828 34520 37856
rect 34333 37819 34391 37825
rect 34514 37816 34520 37828
rect 34572 37816 34578 37868
rect 34624 37865 34652 37896
rect 34609 37859 34667 37865
rect 34609 37825 34621 37859
rect 34655 37825 34667 37859
rect 34609 37819 34667 37825
rect 34701 37859 34759 37865
rect 34701 37825 34713 37859
rect 34747 37825 34759 37859
rect 34701 37819 34759 37825
rect 34716 37788 34744 37819
rect 31726 37760 32812 37788
rect 34164 37760 34744 37788
rect 13964 37692 19472 37720
rect 19521 37723 19579 37729
rect 13964 37680 13970 37692
rect 19521 37689 19533 37723
rect 19567 37720 19579 37723
rect 21266 37720 21272 37732
rect 19567 37692 21272 37720
rect 19567 37689 19579 37692
rect 19521 37683 19579 37689
rect 21266 37680 21272 37692
rect 21324 37680 21330 37732
rect 26510 37680 26516 37732
rect 26568 37720 26574 37732
rect 27430 37720 27436 37732
rect 26568 37692 27436 37720
rect 26568 37680 26574 37692
rect 27430 37680 27436 37692
rect 27488 37720 27494 37732
rect 27488 37692 29960 37720
rect 27488 37680 27494 37692
rect 16942 37652 16948 37664
rect 13832 37624 16948 37652
rect 16942 37612 16948 37624
rect 17000 37612 17006 37664
rect 17494 37612 17500 37664
rect 17552 37652 17558 37664
rect 17773 37655 17831 37661
rect 17773 37652 17785 37655
rect 17552 37624 17785 37652
rect 17552 37612 17558 37624
rect 17773 37621 17785 37624
rect 17819 37621 17831 37655
rect 17773 37615 17831 37621
rect 20625 37655 20683 37661
rect 20625 37621 20637 37655
rect 20671 37652 20683 37655
rect 20990 37652 20996 37664
rect 20671 37624 20996 37652
rect 20671 37621 20683 37624
rect 20625 37615 20683 37621
rect 20990 37612 20996 37624
rect 21048 37612 21054 37664
rect 22278 37612 22284 37664
rect 22336 37652 22342 37664
rect 22557 37655 22615 37661
rect 22557 37652 22569 37655
rect 22336 37624 22569 37652
rect 22336 37612 22342 37624
rect 22557 37621 22569 37624
rect 22603 37621 22615 37655
rect 23106 37652 23112 37664
rect 23067 37624 23112 37652
rect 22557 37615 22615 37621
rect 23106 37612 23112 37624
rect 23164 37612 23170 37664
rect 25590 37652 25596 37664
rect 25551 37624 25596 37652
rect 25590 37612 25596 37624
rect 25648 37612 25654 37664
rect 29932 37652 29960 37692
rect 31481 37655 31539 37661
rect 31481 37652 31493 37655
rect 29932 37624 31493 37652
rect 31481 37621 31493 37624
rect 31527 37652 31539 37655
rect 31726 37652 31754 37760
rect 34164 37664 34192 37760
rect 31527 37624 31754 37652
rect 33873 37655 33931 37661
rect 31527 37621 31539 37624
rect 31481 37615 31539 37621
rect 33873 37621 33885 37655
rect 33919 37652 33931 37655
rect 34146 37652 34152 37664
rect 33919 37624 34152 37652
rect 33919 37621 33931 37624
rect 33873 37615 33931 37621
rect 34146 37612 34152 37624
rect 34204 37612 34210 37664
rect 34977 37655 35035 37661
rect 34977 37621 34989 37655
rect 35023 37652 35035 37655
rect 35342 37652 35348 37664
rect 35023 37624 35348 37652
rect 35023 37621 35035 37624
rect 34977 37615 35035 37621
rect 35342 37612 35348 37624
rect 35400 37612 35406 37664
rect 58158 37652 58164 37664
rect 58119 37624 58164 37652
rect 58158 37612 58164 37624
rect 58216 37612 58222 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 20162 37448 20168 37460
rect 20123 37420 20168 37448
rect 20162 37408 20168 37420
rect 20220 37408 20226 37460
rect 26234 37448 26240 37460
rect 26195 37420 26240 37448
rect 26234 37408 26240 37420
rect 26292 37408 26298 37460
rect 30098 37408 30104 37460
rect 30156 37448 30162 37460
rect 31294 37448 31300 37460
rect 30156 37420 31300 37448
rect 30156 37408 30162 37420
rect 31294 37408 31300 37420
rect 31352 37408 31358 37460
rect 32674 37408 32680 37460
rect 32732 37448 32738 37460
rect 33689 37451 33747 37457
rect 33689 37448 33701 37451
rect 32732 37420 33701 37448
rect 32732 37408 32738 37420
rect 33689 37417 33701 37420
rect 33735 37417 33747 37451
rect 33689 37411 33747 37417
rect 5077 37315 5135 37321
rect 5077 37281 5089 37315
rect 5123 37312 5135 37315
rect 5718 37312 5724 37324
rect 5123 37284 5724 37312
rect 5123 37281 5135 37284
rect 5077 37275 5135 37281
rect 5718 37272 5724 37284
rect 5776 37272 5782 37324
rect 13354 37312 13360 37324
rect 13315 37284 13360 37312
rect 13354 37272 13360 37284
rect 13412 37272 13418 37324
rect 4614 37204 4620 37256
rect 4672 37244 4678 37256
rect 5997 37247 6055 37253
rect 5997 37244 6009 37247
rect 4672 37216 6009 37244
rect 4672 37204 4678 37216
rect 5997 37213 6009 37216
rect 6043 37213 6055 37247
rect 7834 37244 7840 37256
rect 5997 37207 6055 37213
rect 7392 37216 7840 37244
rect 6264 37179 6322 37185
rect 6264 37145 6276 37179
rect 6310 37176 6322 37179
rect 7006 37176 7012 37188
rect 6310 37148 7012 37176
rect 6310 37145 6322 37148
rect 6264 37139 6322 37145
rect 7006 37136 7012 37148
rect 7064 37136 7070 37188
rect 7392 37117 7420 37216
rect 7834 37204 7840 37216
rect 7892 37204 7898 37256
rect 8110 37244 8116 37256
rect 8071 37216 8116 37244
rect 8110 37204 8116 37216
rect 8168 37204 8174 37256
rect 8202 37204 8208 37256
rect 8260 37244 8266 37256
rect 11882 37244 11888 37256
rect 8260 37216 11888 37244
rect 8260 37204 8266 37216
rect 11882 37204 11888 37216
rect 11940 37244 11946 37256
rect 13262 37244 13268 37256
rect 11940 37216 13268 37244
rect 11940 37204 11946 37216
rect 13262 37204 13268 37216
rect 13320 37204 13326 37256
rect 15654 37244 15660 37256
rect 15615 37216 15660 37244
rect 15654 37204 15660 37216
rect 15712 37204 15718 37256
rect 18049 37247 18107 37253
rect 18049 37244 18061 37247
rect 15764 37216 18061 37244
rect 7926 37136 7932 37188
rect 7984 37176 7990 37188
rect 8021 37179 8079 37185
rect 8021 37176 8033 37179
rect 7984 37148 8033 37176
rect 7984 37136 7990 37148
rect 8021 37145 8033 37148
rect 8067 37176 8079 37179
rect 11606 37176 11612 37188
rect 8067 37148 11612 37176
rect 8067 37145 8079 37148
rect 8021 37139 8079 37145
rect 11606 37136 11612 37148
rect 11664 37136 11670 37188
rect 13173 37179 13231 37185
rect 13173 37145 13185 37179
rect 13219 37145 13231 37179
rect 13173 37139 13231 37145
rect 7377 37111 7435 37117
rect 7377 37077 7389 37111
rect 7423 37077 7435 37111
rect 7377 37071 7435 37077
rect 8294 37068 8300 37120
rect 8352 37108 8358 37120
rect 8389 37111 8447 37117
rect 8389 37108 8401 37111
rect 8352 37080 8401 37108
rect 8352 37068 8358 37080
rect 8389 37077 8401 37080
rect 8435 37077 8447 37111
rect 8389 37071 8447 37077
rect 11701 37111 11759 37117
rect 11701 37077 11713 37111
rect 11747 37108 11759 37111
rect 11790 37108 11796 37120
rect 11747 37080 11796 37108
rect 11747 37077 11759 37080
rect 11701 37071 11759 37077
rect 11790 37068 11796 37080
rect 11848 37068 11854 37120
rect 12621 37111 12679 37117
rect 12621 37077 12633 37111
rect 12667 37108 12679 37111
rect 12710 37108 12716 37120
rect 12667 37080 12716 37108
rect 12667 37077 12679 37080
rect 12621 37071 12679 37077
rect 12710 37068 12716 37080
rect 12768 37108 12774 37120
rect 13188 37108 13216 37139
rect 13630 37136 13636 37188
rect 13688 37176 13694 37188
rect 15764 37176 15792 37216
rect 18049 37213 18061 37216
rect 18095 37213 18107 37247
rect 18049 37207 18107 37213
rect 18142 37247 18200 37253
rect 18142 37213 18154 37247
rect 18188 37213 18200 37247
rect 18142 37207 18200 37213
rect 13688 37148 15792 37176
rect 15924 37179 15982 37185
rect 13688 37136 13694 37148
rect 15924 37145 15936 37179
rect 15970 37176 15982 37179
rect 16666 37176 16672 37188
rect 15970 37148 16672 37176
rect 15970 37145 15982 37148
rect 15924 37139 15982 37145
rect 16666 37136 16672 37148
rect 16724 37136 16730 37188
rect 18156 37176 18184 37207
rect 18506 37204 18512 37256
rect 18564 37253 18570 37256
rect 18564 37244 18572 37253
rect 19981 37247 20039 37253
rect 19981 37244 19993 37247
rect 18564 37216 18609 37244
rect 19720 37216 19993 37244
rect 18564 37207 18572 37216
rect 18564 37204 18570 37207
rect 18322 37176 18328 37188
rect 16776 37148 18184 37176
rect 18283 37148 18328 37176
rect 12768 37080 13216 37108
rect 12768 37068 12774 37080
rect 15470 37068 15476 37120
rect 15528 37108 15534 37120
rect 16776 37108 16804 37148
rect 18322 37136 18328 37148
rect 18380 37136 18386 37188
rect 18417 37179 18475 37185
rect 18417 37145 18429 37179
rect 18463 37176 18475 37179
rect 19720 37176 19748 37216
rect 19981 37213 19993 37216
rect 20027 37213 20039 37247
rect 19981 37207 20039 37213
rect 18463 37148 19748 37176
rect 19797 37179 19855 37185
rect 18463 37145 18475 37148
rect 18417 37139 18475 37145
rect 19797 37145 19809 37179
rect 19843 37145 19855 37179
rect 19797 37139 19855 37145
rect 17034 37108 17040 37120
rect 15528 37080 16804 37108
rect 16995 37080 17040 37108
rect 15528 37068 15534 37080
rect 17034 37068 17040 37080
rect 17092 37068 17098 37120
rect 18690 37108 18696 37120
rect 18651 37080 18696 37108
rect 18690 37068 18696 37080
rect 18748 37068 18754 37120
rect 19334 37068 19340 37120
rect 19392 37108 19398 37120
rect 19812 37108 19840 37139
rect 19392 37080 19840 37108
rect 19996 37108 20024 37207
rect 20990 37204 20996 37256
rect 21048 37244 21054 37256
rect 21738 37247 21796 37253
rect 21738 37244 21750 37247
rect 21048 37216 21750 37244
rect 21048 37204 21054 37216
rect 21738 37213 21750 37216
rect 21784 37213 21796 37247
rect 21738 37207 21796 37213
rect 21910 37204 21916 37256
rect 21968 37244 21974 37256
rect 22005 37247 22063 37253
rect 22005 37244 22017 37247
rect 21968 37216 22017 37244
rect 21968 37204 21974 37216
rect 22005 37213 22017 37216
rect 22051 37213 22063 37247
rect 22005 37207 22063 37213
rect 22278 37204 22284 37256
rect 22336 37244 22342 37256
rect 22925 37247 22983 37253
rect 22925 37244 22937 37247
rect 22336 37216 22937 37244
rect 22336 37204 22342 37216
rect 22925 37213 22937 37216
rect 22971 37213 22983 37247
rect 22925 37207 22983 37213
rect 23198 37204 23204 37256
rect 23256 37244 23262 37256
rect 23293 37247 23351 37253
rect 23293 37244 23305 37247
rect 23256 37216 23305 37244
rect 23256 37204 23262 37216
rect 23293 37213 23305 37216
rect 23339 37213 23351 37247
rect 24394 37244 24400 37256
rect 24355 37216 24400 37244
rect 23293 37207 23351 37213
rect 24394 37204 24400 37216
rect 24452 37204 24458 37256
rect 26510 37244 26516 37256
rect 26471 37216 26516 37244
rect 26510 37204 26516 37216
rect 26568 37204 26574 37256
rect 26605 37247 26663 37253
rect 26605 37213 26617 37247
rect 26651 37213 26663 37247
rect 26605 37207 26663 37213
rect 23017 37179 23075 37185
rect 23017 37145 23029 37179
rect 23063 37145 23075 37179
rect 23017 37139 23075 37145
rect 20625 37111 20683 37117
rect 20625 37108 20637 37111
rect 19996 37080 20637 37108
rect 19392 37068 19398 37080
rect 20625 37077 20637 37080
rect 20671 37077 20683 37111
rect 22738 37108 22744 37120
rect 22699 37080 22744 37108
rect 20625 37071 20683 37077
rect 22738 37068 22744 37080
rect 22796 37068 22802 37120
rect 23032 37108 23060 37139
rect 23106 37136 23112 37188
rect 23164 37176 23170 37188
rect 24670 37185 24676 37188
rect 23164 37148 23209 37176
rect 23164 37136 23170 37148
rect 24664 37139 24676 37185
rect 24728 37176 24734 37188
rect 24728 37148 24764 37176
rect 24670 37136 24676 37139
rect 24728 37136 24734 37148
rect 24946 37136 24952 37188
rect 25004 37176 25010 37188
rect 26620 37176 26648 37207
rect 26694 37204 26700 37256
rect 26752 37244 26758 37256
rect 26752 37216 26797 37244
rect 26752 37204 26758 37216
rect 26878 37204 26884 37256
rect 26936 37244 26942 37256
rect 27341 37247 27399 37253
rect 27341 37244 27353 37247
rect 26936 37216 27353 37244
rect 26936 37204 26942 37216
rect 27341 37213 27353 37216
rect 27387 37213 27399 37247
rect 33704 37244 33732 37411
rect 34790 37244 34796 37256
rect 33704 37216 34796 37244
rect 27341 37207 27399 37213
rect 34790 37204 34796 37216
rect 34848 37244 34854 37256
rect 35342 37253 35348 37256
rect 35069 37247 35127 37253
rect 35069 37244 35081 37247
rect 34848 37216 35081 37244
rect 34848 37204 34854 37216
rect 35069 37213 35081 37216
rect 35115 37213 35127 37247
rect 35336 37244 35348 37253
rect 35303 37216 35348 37244
rect 35069 37207 35127 37213
rect 35336 37207 35348 37216
rect 35342 37204 35348 37207
rect 35400 37204 35406 37256
rect 25004 37148 26648 37176
rect 25004 37136 25010 37148
rect 30282 37136 30288 37188
rect 30340 37176 30346 37188
rect 31941 37179 31999 37185
rect 31941 37176 31953 37179
rect 30340 37148 31953 37176
rect 30340 37136 30346 37148
rect 31941 37145 31953 37148
rect 31987 37176 31999 37179
rect 32401 37179 32459 37185
rect 32401 37176 32413 37179
rect 31987 37148 32413 37176
rect 31987 37145 31999 37148
rect 31941 37139 31999 37145
rect 32401 37145 32413 37148
rect 32447 37145 32459 37179
rect 32401 37139 32459 37145
rect 25777 37111 25835 37117
rect 25777 37108 25789 37111
rect 23032 37080 25789 37108
rect 25777 37077 25789 37080
rect 25823 37108 25835 37111
rect 26234 37108 26240 37120
rect 25823 37080 26240 37108
rect 25823 37077 25835 37080
rect 25777 37071 25835 37077
rect 26234 37068 26240 37080
rect 26292 37068 26298 37120
rect 27982 37068 27988 37120
rect 28040 37108 28046 37120
rect 28169 37111 28227 37117
rect 28169 37108 28181 37111
rect 28040 37080 28181 37108
rect 28040 37068 28046 37080
rect 28169 37077 28181 37080
rect 28215 37077 28227 37111
rect 28169 37071 28227 37077
rect 29641 37111 29699 37117
rect 29641 37077 29653 37111
rect 29687 37108 29699 37111
rect 30098 37108 30104 37120
rect 29687 37080 30104 37108
rect 29687 37077 29699 37080
rect 29641 37071 29699 37077
rect 30098 37068 30104 37080
rect 30156 37068 30162 37120
rect 35526 37068 35532 37120
rect 35584 37108 35590 37120
rect 36449 37111 36507 37117
rect 36449 37108 36461 37111
rect 35584 37080 36461 37108
rect 35584 37068 35590 37080
rect 36449 37077 36461 37080
rect 36495 37077 36507 37111
rect 36449 37071 36507 37077
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 12161 36907 12219 36913
rect 12161 36873 12173 36907
rect 12207 36904 12219 36907
rect 15470 36904 15476 36916
rect 12207 36876 15332 36904
rect 15431 36876 15476 36904
rect 12207 36873 12219 36876
rect 12161 36867 12219 36873
rect 6546 36796 6552 36848
rect 6604 36836 6610 36848
rect 6917 36839 6975 36845
rect 6917 36836 6929 36839
rect 6604 36808 6929 36836
rect 6604 36796 6610 36808
rect 6917 36805 6929 36808
rect 6963 36805 6975 36839
rect 7834 36836 7840 36848
rect 7795 36808 7840 36836
rect 6917 36799 6975 36805
rect 7834 36796 7840 36808
rect 7892 36796 7898 36848
rect 8202 36836 8208 36848
rect 7944 36808 8208 36836
rect 5166 36728 5172 36780
rect 5224 36768 5230 36780
rect 6641 36771 6699 36777
rect 6641 36768 6653 36771
rect 5224 36740 6653 36768
rect 5224 36728 5230 36740
rect 6641 36737 6653 36740
rect 6687 36737 6699 36771
rect 6641 36731 6699 36737
rect 6825 36771 6883 36777
rect 6825 36737 6837 36771
rect 6871 36737 6883 36771
rect 6825 36731 6883 36737
rect 7009 36771 7067 36777
rect 7009 36737 7021 36771
rect 7055 36768 7067 36771
rect 7944 36768 7972 36808
rect 8202 36796 8208 36808
rect 8260 36796 8266 36848
rect 7055 36740 7972 36768
rect 7055 36737 7067 36740
rect 7009 36731 7067 36737
rect 6840 36700 6868 36731
rect 8018 36728 8024 36780
rect 8076 36768 8082 36780
rect 8076 36740 8121 36768
rect 8076 36728 8082 36740
rect 9950 36728 9956 36780
rect 10008 36768 10014 36780
rect 12069 36771 12127 36777
rect 12069 36768 12081 36771
rect 10008 36740 12081 36768
rect 10008 36728 10014 36740
rect 12069 36737 12081 36740
rect 12115 36737 12127 36771
rect 12069 36731 12127 36737
rect 12342 36728 12348 36780
rect 12400 36768 12406 36780
rect 14093 36771 14151 36777
rect 14093 36768 14105 36771
rect 12400 36740 14105 36768
rect 12400 36728 12406 36740
rect 14093 36737 14105 36740
rect 14139 36737 14151 36771
rect 14093 36731 14151 36737
rect 14360 36771 14418 36777
rect 14360 36737 14372 36771
rect 14406 36768 14418 36771
rect 14734 36768 14740 36780
rect 14406 36740 14740 36768
rect 14406 36737 14418 36740
rect 14360 36731 14418 36737
rect 14734 36728 14740 36740
rect 14792 36728 14798 36780
rect 7926 36700 7932 36712
rect 6840 36672 7932 36700
rect 7926 36660 7932 36672
rect 7984 36660 7990 36712
rect 13262 36700 13268 36712
rect 13223 36672 13268 36700
rect 13262 36660 13268 36672
rect 13320 36660 13326 36712
rect 13541 36703 13599 36709
rect 13541 36669 13553 36703
rect 13587 36669 13599 36703
rect 13541 36663 13599 36669
rect 12986 36592 12992 36644
rect 13044 36632 13050 36644
rect 13556 36632 13584 36663
rect 13044 36604 13584 36632
rect 15304 36632 15332 36876
rect 15470 36864 15476 36876
rect 15528 36864 15534 36916
rect 16666 36904 16672 36916
rect 16627 36876 16672 36904
rect 16666 36864 16672 36876
rect 16724 36864 16730 36916
rect 18417 36907 18475 36913
rect 18417 36873 18429 36907
rect 18463 36904 18475 36907
rect 19426 36904 19432 36916
rect 18463 36876 19432 36904
rect 18463 36873 18475 36876
rect 18417 36867 18475 36873
rect 19426 36864 19432 36876
rect 19484 36864 19490 36916
rect 30101 36907 30159 36913
rect 30101 36873 30113 36907
rect 30147 36904 30159 36907
rect 30190 36904 30196 36916
rect 30147 36876 30196 36904
rect 30147 36873 30159 36876
rect 30101 36867 30159 36873
rect 30190 36864 30196 36876
rect 30248 36864 30254 36916
rect 32582 36864 32588 36916
rect 32640 36904 32646 36916
rect 32861 36907 32919 36913
rect 32861 36904 32873 36907
rect 32640 36876 32873 36904
rect 32640 36864 32646 36876
rect 32861 36873 32873 36876
rect 32907 36873 32919 36907
rect 32861 36867 32919 36873
rect 34514 36864 34520 36916
rect 34572 36904 34578 36916
rect 35713 36907 35771 36913
rect 35713 36904 35725 36907
rect 34572 36876 35725 36904
rect 34572 36864 34578 36876
rect 35713 36873 35725 36876
rect 35759 36873 35771 36907
rect 35713 36867 35771 36873
rect 17052 36808 18092 36836
rect 16942 36768 16948 36780
rect 16903 36740 16948 36768
rect 16942 36728 16948 36740
rect 17000 36728 17006 36780
rect 17052 36777 17080 36808
rect 17037 36771 17095 36777
rect 17037 36737 17049 36771
rect 17083 36737 17095 36771
rect 17037 36731 17095 36737
rect 16850 36660 16856 36712
rect 16908 36700 16914 36712
rect 17052 36700 17080 36731
rect 17126 36728 17132 36780
rect 17184 36768 17190 36780
rect 18064 36777 18092 36808
rect 18230 36796 18236 36848
rect 18288 36836 18294 36848
rect 19058 36836 19064 36848
rect 18288 36808 18920 36836
rect 19019 36808 19064 36836
rect 18288 36796 18294 36808
rect 17313 36771 17371 36777
rect 17184 36740 17229 36768
rect 17184 36728 17190 36740
rect 17313 36737 17325 36771
rect 17359 36768 17371 36771
rect 17773 36771 17831 36777
rect 17773 36768 17785 36771
rect 17359 36740 17785 36768
rect 17359 36737 17371 36740
rect 17313 36731 17371 36737
rect 17773 36737 17785 36740
rect 17819 36737 17831 36771
rect 17773 36731 17831 36737
rect 17957 36771 18015 36777
rect 17957 36737 17969 36771
rect 18003 36737 18015 36771
rect 17957 36731 18015 36737
rect 18049 36771 18107 36777
rect 18049 36737 18061 36771
rect 18095 36737 18107 36771
rect 18049 36731 18107 36737
rect 16908 36672 17080 36700
rect 16908 36660 16914 36672
rect 17328 36632 17356 36731
rect 15304 36604 17356 36632
rect 17788 36632 17816 36731
rect 17972 36700 18000 36731
rect 18138 36728 18144 36780
rect 18196 36768 18202 36780
rect 18892 36777 18920 36808
rect 19058 36796 19064 36808
rect 19116 36796 19122 36848
rect 21910 36796 21916 36848
rect 21968 36836 21974 36848
rect 23845 36839 23903 36845
rect 23845 36836 23857 36839
rect 21968 36808 23857 36836
rect 21968 36796 21974 36808
rect 23845 36805 23857 36808
rect 23891 36836 23903 36839
rect 24394 36836 24400 36848
rect 23891 36808 24400 36836
rect 23891 36805 23903 36808
rect 23845 36799 23903 36805
rect 24394 36796 24400 36808
rect 24452 36796 24458 36848
rect 25593 36839 25651 36845
rect 25593 36805 25605 36839
rect 25639 36836 25651 36839
rect 27065 36839 27123 36845
rect 27065 36836 27077 36839
rect 25639 36808 27077 36836
rect 25639 36805 25651 36808
rect 25593 36799 25651 36805
rect 27065 36805 27077 36808
rect 27111 36836 27123 36839
rect 28994 36836 29000 36848
rect 27111 36808 29000 36836
rect 27111 36805 27123 36808
rect 27065 36799 27123 36805
rect 28994 36796 29000 36808
rect 29052 36836 29058 36848
rect 30282 36836 30288 36848
rect 29052 36808 30288 36836
rect 29052 36796 29058 36808
rect 30282 36796 30288 36808
rect 30340 36796 30346 36848
rect 33045 36839 33103 36845
rect 33045 36805 33057 36839
rect 33091 36836 33103 36839
rect 33870 36836 33876 36848
rect 33091 36808 33876 36836
rect 33091 36805 33103 36808
rect 33045 36799 33103 36805
rect 33870 36796 33876 36808
rect 33928 36796 33934 36848
rect 34054 36796 34060 36848
rect 34112 36836 34118 36848
rect 34112 36808 34376 36836
rect 34112 36796 34118 36808
rect 18877 36771 18935 36777
rect 18196 36740 18241 36768
rect 18196 36728 18202 36740
rect 18877 36737 18889 36771
rect 18923 36737 18935 36771
rect 22278 36768 22284 36780
rect 22239 36740 22284 36768
rect 18877 36731 18935 36737
rect 22278 36728 22284 36740
rect 22336 36728 22342 36780
rect 22373 36771 22431 36777
rect 22373 36737 22385 36771
rect 22419 36737 22431 36771
rect 22373 36731 22431 36737
rect 19245 36703 19303 36709
rect 19245 36700 19257 36703
rect 17972 36672 19257 36700
rect 19245 36669 19257 36672
rect 19291 36669 19303 36703
rect 22388 36700 22416 36731
rect 22462 36728 22468 36780
rect 22520 36768 22526 36780
rect 22646 36768 22652 36780
rect 22520 36740 22565 36768
rect 22607 36740 22652 36768
rect 22520 36728 22526 36740
rect 22646 36728 22652 36740
rect 22704 36728 22710 36780
rect 25682 36728 25688 36780
rect 25740 36768 25746 36780
rect 26053 36771 26111 36777
rect 26053 36768 26065 36771
rect 25740 36740 26065 36768
rect 25740 36728 25746 36740
rect 26053 36737 26065 36740
rect 26099 36737 26111 36771
rect 26234 36768 26240 36780
rect 26195 36740 26240 36768
rect 26053 36731 26111 36737
rect 26234 36728 26240 36740
rect 26292 36728 26298 36780
rect 27614 36768 27620 36780
rect 27575 36740 27620 36768
rect 27614 36728 27620 36740
rect 27672 36728 27678 36780
rect 27706 36728 27712 36780
rect 27764 36768 27770 36780
rect 27873 36771 27931 36777
rect 27873 36768 27885 36771
rect 27764 36740 27885 36768
rect 27764 36728 27770 36740
rect 27873 36737 27885 36740
rect 27919 36737 27931 36771
rect 27873 36731 27931 36737
rect 28902 36728 28908 36780
rect 28960 36768 28966 36780
rect 29457 36771 29515 36777
rect 29457 36768 29469 36771
rect 28960 36740 29469 36768
rect 28960 36728 28966 36740
rect 29457 36737 29469 36740
rect 29503 36737 29515 36771
rect 29457 36731 29515 36737
rect 29546 36728 29552 36780
rect 29604 36768 29610 36780
rect 29641 36771 29699 36777
rect 29641 36768 29653 36771
rect 29604 36740 29653 36768
rect 29604 36728 29610 36740
rect 29641 36737 29653 36740
rect 29687 36737 29699 36771
rect 29641 36731 29699 36737
rect 29733 36771 29791 36777
rect 29733 36737 29745 36771
rect 29779 36737 29791 36771
rect 29733 36731 29791 36737
rect 29825 36771 29883 36777
rect 29825 36737 29837 36771
rect 29871 36768 29883 36771
rect 30098 36768 30104 36780
rect 29871 36740 30104 36768
rect 29871 36737 29883 36740
rect 29825 36731 29883 36737
rect 25590 36700 25596 36712
rect 22388 36672 25596 36700
rect 19245 36663 19303 36669
rect 25590 36660 25596 36672
rect 25648 36660 25654 36712
rect 29748 36700 29776 36731
rect 30098 36728 30104 36740
rect 30156 36728 30162 36780
rect 31294 36768 31300 36780
rect 31255 36740 31300 36768
rect 31294 36728 31300 36740
rect 31352 36728 31358 36780
rect 33226 36768 33232 36780
rect 33187 36740 33232 36768
rect 33226 36728 33232 36740
rect 33284 36728 33290 36780
rect 34238 36768 34244 36780
rect 34151 36740 34244 36768
rect 34238 36728 34244 36740
rect 34296 36728 34302 36780
rect 34348 36768 34376 36808
rect 34404 36771 34462 36777
rect 34404 36768 34416 36771
rect 34348 36740 34416 36768
rect 34404 36737 34416 36740
rect 34450 36737 34462 36771
rect 34404 36731 34462 36737
rect 34517 36771 34575 36777
rect 34517 36737 34529 36771
rect 34563 36737 34575 36771
rect 34517 36731 34575 36737
rect 34629 36771 34687 36777
rect 34629 36737 34641 36771
rect 34675 36768 34687 36771
rect 35342 36768 35348 36780
rect 34675 36737 34698 36768
rect 35303 36740 35348 36768
rect 34629 36731 34698 36737
rect 30558 36700 30564 36712
rect 29748 36672 30564 36700
rect 30558 36660 30564 36672
rect 30616 36660 30622 36712
rect 31570 36700 31576 36712
rect 31531 36672 31576 36700
rect 31570 36660 31576 36672
rect 31628 36660 31634 36712
rect 33594 36660 33600 36712
rect 33652 36700 33658 36712
rect 34256 36700 34284 36728
rect 34532 36700 34560 36731
rect 33652 36672 34284 36700
rect 34348 36672 34560 36700
rect 33652 36660 33658 36672
rect 18138 36632 18144 36644
rect 17788 36604 18144 36632
rect 13044 36592 13050 36604
rect 18138 36592 18144 36604
rect 18196 36592 18202 36644
rect 34348 36632 34376 36672
rect 34422 36632 34428 36644
rect 34348 36604 34428 36632
rect 34422 36592 34428 36604
rect 34480 36592 34486 36644
rect 34670 36632 34698 36731
rect 35342 36728 35348 36740
rect 35400 36728 35406 36780
rect 35526 36768 35532 36780
rect 35487 36740 35532 36768
rect 35526 36728 35532 36740
rect 35584 36728 35590 36780
rect 34624 36604 34698 36632
rect 7190 36564 7196 36576
rect 7151 36536 7196 36564
rect 7190 36524 7196 36536
rect 7248 36524 7254 36576
rect 7466 36524 7472 36576
rect 7524 36564 7530 36576
rect 7653 36567 7711 36573
rect 7653 36564 7665 36567
rect 7524 36536 7665 36564
rect 7524 36524 7530 36536
rect 7653 36533 7665 36536
rect 7699 36533 7711 36567
rect 7653 36527 7711 36533
rect 19426 36524 19432 36576
rect 19484 36564 19490 36576
rect 19797 36567 19855 36573
rect 19797 36564 19809 36567
rect 19484 36536 19809 36564
rect 19484 36524 19490 36536
rect 19797 36533 19809 36536
rect 19843 36564 19855 36567
rect 20070 36564 20076 36576
rect 19843 36536 20076 36564
rect 19843 36533 19855 36536
rect 19797 36527 19855 36533
rect 20070 36524 20076 36536
rect 20128 36524 20134 36576
rect 21358 36524 21364 36576
rect 21416 36564 21422 36576
rect 22097 36567 22155 36573
rect 22097 36564 22109 36567
rect 21416 36536 22109 36564
rect 21416 36524 21422 36536
rect 22097 36533 22109 36536
rect 22143 36533 22155 36567
rect 22097 36527 22155 36533
rect 22462 36524 22468 36576
rect 22520 36564 22526 36576
rect 22646 36564 22652 36576
rect 22520 36536 22652 36564
rect 22520 36524 22526 36536
rect 22646 36524 22652 36536
rect 22704 36564 22710 36576
rect 23106 36564 23112 36576
rect 22704 36536 23112 36564
rect 22704 36524 22710 36536
rect 23106 36524 23112 36536
rect 23164 36524 23170 36576
rect 25038 36524 25044 36576
rect 25096 36564 25102 36576
rect 26421 36567 26479 36573
rect 26421 36564 26433 36567
rect 25096 36536 26433 36564
rect 25096 36524 25102 36536
rect 26421 36533 26433 36536
rect 26467 36533 26479 36567
rect 26421 36527 26479 36533
rect 28997 36567 29055 36573
rect 28997 36533 29009 36567
rect 29043 36564 29055 36567
rect 29270 36564 29276 36576
rect 29043 36536 29276 36564
rect 29043 36533 29055 36536
rect 28997 36527 29055 36533
rect 29270 36524 29276 36536
rect 29328 36524 29334 36576
rect 33686 36564 33692 36576
rect 33647 36536 33692 36564
rect 33686 36524 33692 36536
rect 33744 36564 33750 36576
rect 34624 36564 34652 36604
rect 33744 36536 34652 36564
rect 33744 36524 33750 36536
rect 34698 36524 34704 36576
rect 34756 36564 34762 36576
rect 34885 36567 34943 36573
rect 34885 36564 34897 36567
rect 34756 36536 34897 36564
rect 34756 36524 34762 36536
rect 34885 36533 34897 36536
rect 34931 36533 34943 36567
rect 34885 36527 34943 36533
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 5166 36360 5172 36372
rect 5127 36332 5172 36360
rect 5166 36320 5172 36332
rect 5224 36320 5230 36372
rect 7006 36360 7012 36372
rect 6967 36332 7012 36360
rect 7006 36320 7012 36332
rect 7064 36320 7070 36372
rect 9490 36360 9496 36372
rect 9451 36332 9496 36360
rect 9490 36320 9496 36332
rect 9548 36320 9554 36372
rect 11422 36320 11428 36372
rect 11480 36360 11486 36372
rect 12342 36360 12348 36372
rect 11480 36332 12348 36360
rect 11480 36320 11486 36332
rect 12342 36320 12348 36332
rect 12400 36360 12406 36372
rect 13081 36363 13139 36369
rect 13081 36360 13093 36363
rect 12400 36332 13093 36360
rect 12400 36320 12406 36332
rect 13081 36329 13093 36332
rect 13127 36329 13139 36363
rect 14734 36360 14740 36372
rect 14695 36332 14740 36360
rect 13081 36323 13139 36329
rect 14734 36320 14740 36332
rect 14792 36320 14798 36372
rect 16669 36363 16727 36369
rect 16669 36329 16681 36363
rect 16715 36360 16727 36363
rect 17126 36360 17132 36372
rect 16715 36332 17132 36360
rect 16715 36329 16727 36332
rect 16669 36323 16727 36329
rect 17126 36320 17132 36332
rect 17184 36320 17190 36372
rect 18046 36320 18052 36372
rect 18104 36360 18110 36372
rect 18509 36363 18567 36369
rect 18509 36360 18521 36363
rect 18104 36332 18521 36360
rect 18104 36320 18110 36332
rect 18509 36329 18521 36332
rect 18555 36329 18567 36363
rect 18509 36323 18567 36329
rect 24581 36363 24639 36369
rect 24581 36329 24593 36363
rect 24627 36360 24639 36363
rect 24670 36360 24676 36372
rect 24627 36332 24676 36360
rect 24627 36329 24639 36332
rect 24581 36323 24639 36329
rect 24670 36320 24676 36332
rect 24728 36320 24734 36372
rect 26053 36363 26111 36369
rect 26053 36329 26065 36363
rect 26099 36360 26111 36363
rect 26694 36360 26700 36372
rect 26099 36332 26700 36360
rect 26099 36329 26111 36332
rect 26053 36323 26111 36329
rect 26694 36320 26700 36332
rect 26752 36320 26758 36372
rect 27706 36360 27712 36372
rect 27667 36332 27712 36360
rect 27706 36320 27712 36332
rect 27764 36320 27770 36372
rect 29546 36360 29552 36372
rect 29507 36332 29552 36360
rect 29546 36320 29552 36332
rect 29604 36320 29610 36372
rect 34054 36320 34060 36372
rect 34112 36360 34118 36372
rect 34149 36363 34207 36369
rect 34149 36360 34161 36363
rect 34112 36332 34161 36360
rect 34112 36320 34118 36332
rect 34149 36329 34161 36332
rect 34195 36329 34207 36363
rect 34149 36323 34207 36329
rect 24762 36252 24768 36304
rect 24820 36292 24826 36304
rect 25682 36292 25688 36304
rect 24820 36264 25688 36292
rect 24820 36252 24826 36264
rect 25682 36252 25688 36264
rect 25740 36252 25746 36304
rect 16850 36224 16856 36236
rect 14384 36196 16856 36224
rect 14384 36168 14412 36196
rect 16850 36184 16856 36196
rect 16908 36184 16914 36236
rect 24302 36184 24308 36236
rect 24360 36224 24366 36236
rect 26878 36224 26884 36236
rect 24360 36196 26884 36224
rect 24360 36184 24366 36196
rect 2498 36116 2504 36168
rect 2556 36156 2562 36168
rect 3789 36159 3847 36165
rect 3789 36156 3801 36159
rect 2556 36128 3801 36156
rect 2556 36116 2562 36128
rect 3789 36125 3801 36128
rect 3835 36156 3847 36159
rect 4614 36156 4620 36168
rect 3835 36128 4620 36156
rect 3835 36125 3847 36128
rect 3789 36119 3847 36125
rect 4614 36116 4620 36128
rect 4672 36116 4678 36168
rect 7239 36159 7297 36165
rect 7239 36156 7251 36159
rect 6564 36128 7251 36156
rect 4056 36091 4114 36097
rect 4056 36057 4068 36091
rect 4102 36088 4114 36091
rect 4102 36060 4660 36088
rect 4102 36057 4114 36060
rect 4056 36051 4114 36057
rect 4632 36032 4660 36060
rect 6564 36032 6592 36128
rect 7239 36125 7251 36128
rect 7285 36125 7297 36159
rect 7374 36156 7380 36168
rect 7335 36128 7380 36156
rect 7239 36119 7297 36125
rect 7374 36116 7380 36128
rect 7432 36116 7438 36168
rect 7466 36116 7472 36168
rect 7524 36165 7530 36168
rect 7524 36156 7532 36165
rect 7653 36159 7711 36165
rect 7524 36128 7569 36156
rect 7524 36119 7532 36128
rect 7653 36125 7665 36159
rect 7699 36125 7711 36159
rect 7653 36119 7711 36125
rect 7524 36116 7530 36119
rect 7668 36088 7696 36119
rect 8938 36116 8944 36168
rect 8996 36156 9002 36168
rect 9309 36159 9367 36165
rect 9309 36156 9321 36159
rect 8996 36128 9321 36156
rect 8996 36116 9002 36128
rect 9309 36125 9321 36128
rect 9355 36125 9367 36159
rect 9309 36119 9367 36125
rect 9858 36116 9864 36168
rect 9916 36156 9922 36168
rect 9953 36159 10011 36165
rect 9953 36156 9965 36159
rect 9916 36128 9965 36156
rect 9916 36116 9922 36128
rect 9953 36125 9965 36128
rect 9999 36125 10011 36159
rect 14090 36156 14096 36168
rect 14051 36128 14096 36156
rect 9953 36119 10011 36125
rect 14090 36116 14096 36128
rect 14148 36116 14154 36168
rect 14277 36159 14335 36165
rect 14277 36125 14289 36159
rect 14323 36125 14335 36159
rect 14277 36119 14335 36125
rect 10220 36091 10278 36097
rect 7668 36060 9674 36088
rect 4614 35980 4620 36032
rect 4672 35980 4678 36032
rect 6546 36020 6552 36032
rect 6507 35992 6552 36020
rect 6546 35980 6552 35992
rect 6604 35980 6610 36032
rect 9646 36020 9674 36060
rect 10220 36057 10232 36091
rect 10266 36088 10278 36091
rect 10318 36088 10324 36100
rect 10266 36060 10324 36088
rect 10266 36057 10278 36060
rect 10220 36051 10278 36057
rect 10318 36048 10324 36060
rect 10376 36048 10382 36100
rect 11790 36088 11796 36100
rect 11751 36060 11796 36088
rect 11790 36048 11796 36060
rect 11848 36048 11854 36100
rect 14292 36088 14320 36119
rect 14366 36116 14372 36168
rect 14424 36156 14430 36168
rect 14507 36159 14565 36165
rect 14424 36128 14469 36156
rect 14424 36116 14430 36128
rect 14507 36125 14519 36159
rect 14553 36156 14565 36159
rect 15010 36156 15016 36168
rect 14553 36128 15016 36156
rect 14553 36125 14565 36128
rect 14507 36119 14565 36125
rect 15010 36116 15016 36128
rect 15068 36116 15074 36168
rect 15381 36159 15439 36165
rect 15381 36125 15393 36159
rect 15427 36156 15439 36159
rect 15470 36156 15476 36168
rect 15427 36128 15476 36156
rect 15427 36125 15439 36128
rect 15381 36119 15439 36125
rect 15470 36116 15476 36128
rect 15528 36116 15534 36168
rect 16485 36159 16543 36165
rect 16485 36125 16497 36159
rect 16531 36156 16543 36159
rect 17034 36156 17040 36168
rect 16531 36128 17040 36156
rect 16531 36125 16543 36128
rect 16485 36119 16543 36125
rect 17034 36116 17040 36128
rect 17092 36116 17098 36168
rect 24670 36116 24676 36168
rect 24728 36156 24734 36168
rect 24811 36159 24869 36165
rect 24811 36156 24823 36159
rect 24728 36128 24823 36156
rect 24728 36116 24734 36128
rect 24811 36125 24823 36128
rect 24857 36125 24869 36159
rect 24946 36156 24952 36168
rect 24907 36128 24952 36156
rect 24811 36119 24869 36125
rect 24946 36116 24952 36128
rect 25004 36116 25010 36168
rect 25038 36116 25044 36168
rect 25096 36156 25102 36168
rect 25240 36165 25268 36196
rect 26878 36184 26884 36196
rect 26936 36184 26942 36236
rect 30558 36224 30564 36236
rect 28092 36196 30564 36224
rect 25225 36159 25283 36165
rect 25096 36128 25141 36156
rect 25096 36116 25102 36128
rect 25225 36125 25237 36159
rect 25271 36125 25283 36159
rect 25225 36119 25283 36125
rect 25590 36116 25596 36168
rect 25648 36156 25654 36168
rect 25869 36159 25927 36165
rect 25869 36156 25881 36159
rect 25648 36128 25881 36156
rect 25648 36116 25654 36128
rect 25869 36125 25881 36128
rect 25915 36125 25927 36159
rect 27982 36156 27988 36168
rect 25869 36119 25927 36125
rect 27172 36128 27988 36156
rect 15197 36091 15255 36097
rect 15197 36088 15209 36091
rect 14292 36060 15209 36088
rect 15197 36057 15209 36060
rect 15243 36057 15255 36091
rect 15197 36051 15255 36057
rect 15565 36091 15623 36097
rect 15565 36057 15577 36091
rect 15611 36088 15623 36091
rect 15654 36088 15660 36100
rect 15611 36060 15660 36088
rect 15611 36057 15623 36060
rect 15565 36051 15623 36057
rect 15654 36048 15660 36060
rect 15712 36088 15718 36100
rect 16301 36091 16359 36097
rect 16301 36088 16313 36091
rect 15712 36060 16313 36088
rect 15712 36048 15718 36060
rect 16301 36057 16313 36060
rect 16347 36088 16359 36091
rect 18230 36088 18236 36100
rect 16347 36060 18236 36088
rect 16347 36057 16359 36060
rect 16301 36051 16359 36057
rect 18230 36048 18236 36060
rect 18288 36048 18294 36100
rect 25682 36088 25688 36100
rect 25643 36060 25688 36088
rect 25682 36048 25688 36060
rect 25740 36048 25746 36100
rect 27172 36032 27200 36128
rect 27982 36116 27988 36128
rect 28040 36116 28046 36168
rect 28092 36165 28120 36196
rect 30558 36184 30564 36196
rect 30616 36184 30622 36236
rect 34790 36224 34796 36236
rect 34751 36196 34796 36224
rect 34790 36184 34796 36196
rect 34848 36184 34854 36236
rect 28077 36159 28135 36165
rect 28077 36125 28089 36159
rect 28123 36125 28135 36159
rect 28077 36119 28135 36125
rect 28166 36116 28172 36168
rect 28224 36156 28230 36168
rect 28353 36159 28411 36165
rect 28224 36128 28269 36156
rect 28224 36116 28230 36128
rect 28353 36125 28365 36159
rect 28399 36125 28411 36159
rect 29730 36156 29736 36168
rect 29691 36128 29736 36156
rect 28353 36119 28411 36125
rect 27890 36048 27896 36100
rect 27948 36088 27954 36100
rect 28368 36088 28396 36119
rect 29730 36116 29736 36128
rect 29788 36116 29794 36168
rect 31849 36159 31907 36165
rect 31849 36156 31861 36159
rect 31726 36128 31861 36156
rect 28902 36088 28908 36100
rect 27948 36060 28908 36088
rect 27948 36048 27954 36060
rect 28902 36048 28908 36060
rect 28960 36048 28966 36100
rect 29914 36088 29920 36100
rect 29875 36060 29920 36088
rect 29914 36048 29920 36060
rect 29972 36048 29978 36100
rect 10134 36020 10140 36032
rect 9646 35992 10140 36020
rect 10134 35980 10140 35992
rect 10192 35980 10198 36032
rect 11330 36020 11336 36032
rect 11291 35992 11336 36020
rect 11330 35980 11336 35992
rect 11388 35980 11394 36032
rect 16942 35980 16948 36032
rect 17000 36020 17006 36032
rect 17497 36023 17555 36029
rect 17497 36020 17509 36023
rect 17000 35992 17509 36020
rect 17000 35980 17006 35992
rect 17497 35989 17509 35992
rect 17543 36020 17555 36023
rect 18598 36020 18604 36032
rect 17543 35992 18604 36020
rect 17543 35989 17555 35992
rect 17497 35983 17555 35989
rect 18598 35980 18604 35992
rect 18656 35980 18662 36032
rect 22557 36023 22615 36029
rect 22557 35989 22569 36023
rect 22603 36020 22615 36023
rect 22646 36020 22652 36032
rect 22603 35992 22652 36020
rect 22603 35989 22615 35992
rect 22557 35983 22615 35989
rect 22646 35980 22652 35992
rect 22704 35980 22710 36032
rect 23014 36020 23020 36032
rect 22975 35992 23020 36020
rect 23014 35980 23020 35992
rect 23072 35980 23078 36032
rect 27154 36020 27160 36032
rect 27115 35992 27160 36020
rect 27154 35980 27160 35992
rect 27212 35980 27218 36032
rect 30650 36020 30656 36032
rect 30611 35992 30656 36020
rect 30650 35980 30656 35992
rect 30708 36020 30714 36032
rect 31297 36023 31355 36029
rect 31297 36020 31309 36023
rect 30708 35992 31309 36020
rect 30708 35980 30714 35992
rect 31297 35989 31309 35992
rect 31343 36020 31355 36023
rect 31570 36020 31576 36032
rect 31343 35992 31576 36020
rect 31343 35989 31355 35992
rect 31297 35983 31355 35989
rect 31570 35980 31576 35992
rect 31628 36020 31634 36032
rect 31726 36020 31754 36128
rect 31849 36125 31861 36128
rect 31895 36125 31907 36159
rect 31849 36119 31907 36125
rect 32125 36159 32183 36165
rect 32125 36125 32137 36159
rect 32171 36156 32183 36159
rect 33594 36156 33600 36168
rect 32171 36128 33600 36156
rect 32171 36125 32183 36128
rect 32125 36119 32183 36125
rect 33594 36116 33600 36128
rect 33652 36116 33658 36168
rect 33778 36156 33784 36168
rect 33739 36128 33784 36156
rect 33778 36116 33784 36128
rect 33836 36116 33842 36168
rect 34698 36116 34704 36168
rect 34756 36156 34762 36168
rect 35049 36159 35107 36165
rect 35049 36156 35061 36159
rect 34756 36128 35061 36156
rect 34756 36116 34762 36128
rect 35049 36125 35061 36128
rect 35095 36125 35107 36159
rect 58158 36156 58164 36168
rect 58119 36128 58164 36156
rect 35049 36119 35107 36125
rect 58158 36116 58164 36128
rect 58216 36116 58222 36168
rect 33965 36091 34023 36097
rect 33965 36057 33977 36091
rect 34011 36057 34023 36091
rect 33965 36051 34023 36057
rect 31628 35992 31754 36020
rect 33980 36020 34008 36051
rect 34698 36020 34704 36032
rect 33980 35992 34704 36020
rect 31628 35980 31634 35992
rect 34698 35980 34704 35992
rect 34756 36020 34762 36032
rect 36173 36023 36231 36029
rect 36173 36020 36185 36023
rect 34756 35992 36185 36020
rect 34756 35980 34762 35992
rect 36173 35989 36185 35992
rect 36219 35989 36231 36023
rect 36173 35983 36231 35989
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 9766 35776 9772 35828
rect 9824 35816 9830 35828
rect 13909 35819 13967 35825
rect 13909 35816 13921 35819
rect 9824 35788 13921 35816
rect 9824 35776 9830 35788
rect 13909 35785 13921 35788
rect 13955 35816 13967 35819
rect 14090 35816 14096 35828
rect 13955 35788 14096 35816
rect 13955 35785 13967 35788
rect 13909 35779 13967 35785
rect 14090 35776 14096 35788
rect 14148 35776 14154 35828
rect 27341 35819 27399 35825
rect 27341 35816 27353 35819
rect 14200 35788 27353 35816
rect 4617 35751 4675 35757
rect 4617 35717 4629 35751
rect 4663 35748 4675 35751
rect 5166 35748 5172 35760
rect 4663 35720 5172 35748
rect 4663 35717 4675 35720
rect 4617 35711 4675 35717
rect 5166 35708 5172 35720
rect 5224 35708 5230 35760
rect 6564 35720 7604 35748
rect 4433 35683 4491 35689
rect 4433 35649 4445 35683
rect 4479 35680 4491 35683
rect 4890 35680 4896 35692
rect 4479 35652 4896 35680
rect 4479 35649 4491 35652
rect 4433 35643 4491 35649
rect 4890 35640 4896 35652
rect 4948 35680 4954 35692
rect 6564 35680 6592 35720
rect 7466 35680 7472 35692
rect 7524 35689 7530 35692
rect 4948 35652 6592 35680
rect 7436 35652 7472 35680
rect 4948 35640 4954 35652
rect 7466 35640 7472 35652
rect 7524 35643 7536 35689
rect 7576 35680 7604 35720
rect 11054 35708 11060 35760
rect 11112 35748 11118 35760
rect 11514 35748 11520 35760
rect 11112 35720 11520 35748
rect 11112 35708 11118 35720
rect 11514 35708 11520 35720
rect 11572 35708 11578 35760
rect 11606 35708 11612 35760
rect 11664 35748 11670 35760
rect 11664 35720 12434 35748
rect 11664 35708 11670 35720
rect 7745 35683 7803 35689
rect 7576 35652 7696 35680
rect 7524 35640 7530 35643
rect 7668 35612 7696 35652
rect 7745 35649 7757 35683
rect 7791 35680 7803 35683
rect 9858 35680 9864 35692
rect 7791 35652 9864 35680
rect 7791 35649 7803 35652
rect 7745 35643 7803 35649
rect 9858 35640 9864 35652
rect 9916 35640 9922 35692
rect 9950 35640 9956 35692
rect 10008 35680 10014 35692
rect 10008 35652 10053 35680
rect 10008 35640 10014 35652
rect 10134 35640 10140 35692
rect 10192 35680 10198 35692
rect 10229 35683 10287 35689
rect 10229 35680 10241 35683
rect 10192 35652 10241 35680
rect 10192 35640 10198 35652
rect 10229 35649 10241 35652
rect 10275 35680 10287 35683
rect 10778 35680 10784 35692
rect 10275 35652 10784 35680
rect 10275 35649 10287 35652
rect 10229 35643 10287 35649
rect 10778 35640 10784 35652
rect 10836 35680 10842 35692
rect 10962 35680 10968 35692
rect 10836 35652 10968 35680
rect 10836 35640 10842 35652
rect 10962 35640 10968 35652
rect 11020 35640 11026 35692
rect 11698 35680 11704 35692
rect 11659 35652 11704 35680
rect 11698 35640 11704 35652
rect 11756 35640 11762 35692
rect 12406 35680 12434 35720
rect 13354 35708 13360 35760
rect 13412 35748 13418 35760
rect 13630 35748 13636 35760
rect 13412 35720 13636 35748
rect 13412 35708 13418 35720
rect 13630 35708 13636 35720
rect 13688 35748 13694 35760
rect 14200 35748 14228 35788
rect 27341 35785 27353 35788
rect 27387 35816 27399 35819
rect 27890 35816 27896 35828
rect 27387 35788 27896 35816
rect 27387 35785 27399 35788
rect 27341 35779 27399 35785
rect 27890 35776 27896 35788
rect 27948 35776 27954 35828
rect 28166 35776 28172 35828
rect 28224 35816 28230 35828
rect 28353 35819 28411 35825
rect 28353 35816 28365 35819
rect 28224 35788 28365 35816
rect 28224 35776 28230 35788
rect 28353 35785 28365 35788
rect 28399 35785 28411 35819
rect 28353 35779 28411 35785
rect 28626 35776 28632 35828
rect 28684 35816 28690 35828
rect 30098 35816 30104 35828
rect 28684 35788 30104 35816
rect 28684 35776 28690 35788
rect 30098 35776 30104 35788
rect 30156 35776 30162 35828
rect 30558 35776 30564 35828
rect 30616 35816 30622 35828
rect 30616 35788 30696 35816
rect 30616 35776 30622 35788
rect 13688 35720 14228 35748
rect 14921 35751 14979 35757
rect 13688 35708 13694 35720
rect 14921 35717 14933 35751
rect 14967 35748 14979 35751
rect 15010 35748 15016 35760
rect 14967 35720 15016 35748
rect 14967 35717 14979 35720
rect 14921 35711 14979 35717
rect 15010 35708 15016 35720
rect 15068 35708 15074 35760
rect 18230 35748 18236 35760
rect 18191 35720 18236 35748
rect 18230 35708 18236 35720
rect 18288 35708 18294 35760
rect 22646 35708 22652 35760
rect 22704 35748 22710 35760
rect 23201 35751 23259 35757
rect 23201 35748 23213 35751
rect 22704 35720 23213 35748
rect 22704 35708 22710 35720
rect 23201 35717 23213 35720
rect 23247 35717 23259 35751
rect 23201 35711 23259 35717
rect 28537 35751 28595 35757
rect 28537 35717 28549 35751
rect 28583 35748 28595 35751
rect 29270 35748 29276 35760
rect 28583 35720 29276 35748
rect 28583 35717 28595 35720
rect 28537 35711 28595 35717
rect 29270 35708 29276 35720
rect 29328 35708 29334 35760
rect 30668 35748 30696 35788
rect 30576 35720 30696 35748
rect 13081 35683 13139 35689
rect 13081 35680 13093 35683
rect 12406 35652 13093 35680
rect 13081 35649 13093 35652
rect 13127 35649 13139 35683
rect 18046 35680 18052 35692
rect 18007 35652 18052 35680
rect 13081 35643 13139 35649
rect 18046 35640 18052 35652
rect 18104 35640 18110 35692
rect 22370 35640 22376 35692
rect 22428 35680 22434 35692
rect 23014 35680 23020 35692
rect 22428 35652 23020 35680
rect 22428 35640 22434 35652
rect 23014 35640 23020 35652
rect 23072 35640 23078 35692
rect 23106 35640 23112 35692
rect 23164 35680 23170 35692
rect 23385 35683 23443 35689
rect 23164 35652 23209 35680
rect 23164 35640 23170 35652
rect 23385 35649 23397 35683
rect 23431 35680 23443 35683
rect 24854 35680 24860 35692
rect 23431 35652 24860 35680
rect 23431 35649 23443 35652
rect 23385 35643 23443 35649
rect 24854 35640 24860 35652
rect 24912 35640 24918 35692
rect 28721 35683 28779 35689
rect 28721 35649 28733 35683
rect 28767 35680 28779 35683
rect 29914 35680 29920 35692
rect 28767 35652 29920 35680
rect 28767 35649 28779 35652
rect 28721 35643 28779 35649
rect 29914 35640 29920 35652
rect 29972 35640 29978 35692
rect 30190 35640 30196 35692
rect 30248 35680 30254 35692
rect 30576 35689 30604 35720
rect 30285 35683 30343 35689
rect 30285 35680 30297 35683
rect 30248 35652 30297 35680
rect 30248 35640 30254 35652
rect 30285 35649 30297 35652
rect 30331 35649 30343 35683
rect 30448 35683 30506 35689
rect 30448 35680 30460 35683
rect 30285 35643 30343 35649
rect 30392 35652 30460 35680
rect 8018 35612 8024 35624
rect 7668 35584 8024 35612
rect 8018 35572 8024 35584
rect 8076 35612 8082 35624
rect 8757 35615 8815 35621
rect 8757 35612 8769 35615
rect 8076 35584 8769 35612
rect 8076 35572 8082 35584
rect 8757 35581 8769 35584
rect 8803 35581 8815 35615
rect 8757 35575 8815 35581
rect 8938 35572 8944 35624
rect 8996 35612 9002 35624
rect 9033 35615 9091 35621
rect 9033 35612 9045 35615
rect 8996 35584 9045 35612
rect 8996 35572 9002 35584
rect 9033 35581 9045 35584
rect 9079 35581 9091 35615
rect 9033 35575 9091 35581
rect 13357 35615 13415 35621
rect 13357 35581 13369 35615
rect 13403 35612 13415 35615
rect 13538 35612 13544 35624
rect 13403 35584 13544 35612
rect 13403 35581 13415 35584
rect 13357 35575 13415 35581
rect 13538 35572 13544 35584
rect 13596 35572 13602 35624
rect 17034 35504 17040 35556
rect 17092 35544 17098 35556
rect 29733 35547 29791 35553
rect 29733 35544 29745 35547
rect 17092 35516 29745 35544
rect 17092 35504 17098 35516
rect 29733 35513 29745 35516
rect 29779 35544 29791 35547
rect 29822 35544 29828 35556
rect 29779 35516 29828 35544
rect 29779 35513 29791 35516
rect 29733 35507 29791 35513
rect 29822 35504 29828 35516
rect 29880 35504 29886 35556
rect 30392 35544 30420 35652
rect 30448 35649 30460 35652
rect 30494 35649 30506 35683
rect 30448 35643 30506 35649
rect 30561 35683 30619 35689
rect 30561 35649 30573 35683
rect 30607 35649 30619 35683
rect 30561 35643 30619 35649
rect 30653 35683 30711 35689
rect 30653 35649 30665 35683
rect 30699 35655 30880 35683
rect 30699 35649 30711 35655
rect 30653 35643 30711 35649
rect 30466 35544 30472 35556
rect 30392 35516 30472 35544
rect 30466 35504 30472 35516
rect 30524 35504 30530 35556
rect 30852 35544 30880 35655
rect 30760 35516 30880 35544
rect 4798 35476 4804 35488
rect 4759 35448 4804 35476
rect 4798 35436 4804 35448
rect 4856 35436 4862 35488
rect 6365 35479 6423 35485
rect 6365 35445 6377 35479
rect 6411 35476 6423 35479
rect 6638 35476 6644 35488
rect 6411 35448 6644 35476
rect 6411 35445 6423 35448
rect 6365 35439 6423 35445
rect 6638 35436 6644 35448
rect 6696 35436 6702 35488
rect 10962 35436 10968 35488
rect 11020 35476 11026 35488
rect 11885 35479 11943 35485
rect 11885 35476 11897 35479
rect 11020 35448 11897 35476
rect 11020 35436 11026 35448
rect 11885 35445 11897 35448
rect 11931 35445 11943 35479
rect 11885 35439 11943 35445
rect 17865 35479 17923 35485
rect 17865 35445 17877 35479
rect 17911 35476 17923 35479
rect 17954 35476 17960 35488
rect 17911 35448 17960 35476
rect 17911 35445 17923 35448
rect 17865 35439 17923 35445
rect 17954 35436 17960 35448
rect 18012 35436 18018 35488
rect 22370 35476 22376 35488
rect 22331 35448 22376 35476
rect 22370 35436 22376 35448
rect 22428 35436 22434 35488
rect 22833 35479 22891 35485
rect 22833 35445 22845 35479
rect 22879 35476 22891 35479
rect 23014 35476 23020 35488
rect 22879 35448 23020 35476
rect 22879 35445 22891 35448
rect 22833 35439 22891 35445
rect 23014 35436 23020 35448
rect 23072 35436 23078 35488
rect 24302 35436 24308 35488
rect 24360 35476 24366 35488
rect 24397 35479 24455 35485
rect 24397 35476 24409 35479
rect 24360 35448 24409 35476
rect 24360 35436 24366 35448
rect 24397 35445 24409 35448
rect 24443 35445 24455 35479
rect 24397 35439 24455 35445
rect 24670 35436 24676 35488
rect 24728 35476 24734 35488
rect 25314 35476 25320 35488
rect 24728 35448 25320 35476
rect 24728 35436 24734 35448
rect 25314 35436 25320 35448
rect 25372 35476 25378 35488
rect 25409 35479 25467 35485
rect 25409 35476 25421 35479
rect 25372 35448 25421 35476
rect 25372 35436 25378 35448
rect 25409 35445 25421 35448
rect 25455 35476 25467 35479
rect 25958 35476 25964 35488
rect 25455 35448 25964 35476
rect 25455 35445 25467 35448
rect 25409 35439 25467 35445
rect 25958 35436 25964 35448
rect 26016 35436 26022 35488
rect 29840 35476 29868 35504
rect 30760 35476 30788 35516
rect 30926 35476 30932 35488
rect 29840 35448 30788 35476
rect 30887 35448 30932 35476
rect 30926 35436 30932 35448
rect 30984 35436 30990 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 4341 35275 4399 35281
rect 4341 35241 4353 35275
rect 4387 35272 4399 35275
rect 4614 35272 4620 35284
rect 4387 35244 4620 35272
rect 4387 35241 4399 35244
rect 4341 35235 4399 35241
rect 4614 35232 4620 35244
rect 4672 35232 4678 35284
rect 7285 35275 7343 35281
rect 7285 35241 7297 35275
rect 7331 35272 7343 35275
rect 7466 35272 7472 35284
rect 7331 35244 7472 35272
rect 7331 35241 7343 35244
rect 7285 35235 7343 35241
rect 7466 35232 7472 35244
rect 7524 35232 7530 35284
rect 18046 35232 18052 35284
rect 18104 35272 18110 35284
rect 18693 35275 18751 35281
rect 18693 35272 18705 35275
rect 18104 35244 18705 35272
rect 18104 35232 18110 35244
rect 18693 35241 18705 35244
rect 18739 35241 18751 35275
rect 18693 35235 18751 35241
rect 25958 35232 25964 35284
rect 26016 35272 26022 35284
rect 30098 35272 30104 35284
rect 26016 35244 30104 35272
rect 26016 35232 26022 35244
rect 30098 35232 30104 35244
rect 30156 35232 30162 35284
rect 30285 35275 30343 35281
rect 30285 35241 30297 35275
rect 30331 35272 30343 35275
rect 30466 35272 30472 35284
rect 30331 35244 30472 35272
rect 30331 35241 30343 35244
rect 30285 35235 30343 35241
rect 30466 35232 30472 35244
rect 30524 35232 30530 35284
rect 7374 35204 7380 35216
rect 4724 35176 7380 35204
rect 3234 35096 3240 35148
rect 3292 35136 3298 35148
rect 4724 35136 4752 35176
rect 7374 35164 7380 35176
rect 7432 35164 7438 35216
rect 9033 35207 9091 35213
rect 9033 35173 9045 35207
rect 9079 35204 9091 35207
rect 9079 35176 17172 35204
rect 9079 35173 9091 35176
rect 9033 35167 9091 35173
rect 3292 35108 4752 35136
rect 3292 35096 3298 35108
rect 4724 35077 4752 35108
rect 6825 35139 6883 35145
rect 6825 35105 6837 35139
rect 6871 35136 6883 35139
rect 6871 35108 7788 35136
rect 6871 35105 6883 35108
rect 6825 35099 6883 35105
rect 4617 35071 4675 35077
rect 4617 35037 4629 35071
rect 4663 35037 4675 35071
rect 4617 35031 4675 35037
rect 4709 35071 4767 35077
rect 4709 35037 4721 35071
rect 4755 35037 4767 35071
rect 4709 35031 4767 35037
rect 4632 35000 4660 35031
rect 4798 35028 4804 35080
rect 4856 35068 4862 35080
rect 4856 35040 4901 35068
rect 4856 35028 4862 35040
rect 4982 35028 4988 35080
rect 5040 35068 5046 35080
rect 7558 35068 7564 35080
rect 5040 35040 5085 35068
rect 7519 35040 7564 35068
rect 5040 35028 5046 35040
rect 7558 35028 7564 35040
rect 7616 35028 7622 35080
rect 7760 35077 7788 35108
rect 7653 35071 7711 35077
rect 7653 35037 7665 35071
rect 7699 35037 7711 35071
rect 7653 35031 7711 35037
rect 7745 35071 7803 35077
rect 7745 35037 7757 35071
rect 7791 35037 7803 35071
rect 7745 35031 7803 35037
rect 7929 35071 7987 35077
rect 7929 35037 7941 35071
rect 7975 35068 7987 35071
rect 9048 35068 9076 35167
rect 9769 35139 9827 35145
rect 9769 35105 9781 35139
rect 9815 35136 9827 35139
rect 10410 35136 10416 35148
rect 9815 35108 10416 35136
rect 9815 35105 9827 35108
rect 9769 35099 9827 35105
rect 10410 35096 10416 35108
rect 10468 35136 10474 35148
rect 10686 35136 10692 35148
rect 10468 35108 10692 35136
rect 10468 35096 10474 35108
rect 10686 35096 10692 35108
rect 10744 35136 10750 35148
rect 11974 35136 11980 35148
rect 10744 35108 11100 35136
rect 10744 35096 10750 35108
rect 7975 35040 9076 35068
rect 9493 35071 9551 35077
rect 7975 35037 7987 35040
rect 7929 35031 7987 35037
rect 9493 35037 9505 35071
rect 9539 35068 9551 35071
rect 9582 35068 9588 35080
rect 9539 35040 9588 35068
rect 9539 35037 9551 35040
rect 9493 35031 9551 35037
rect 4632 34972 5580 35000
rect 5552 34941 5580 34972
rect 5626 34960 5632 35012
rect 5684 35000 5690 35012
rect 6457 35003 6515 35009
rect 6457 35000 6469 35003
rect 5684 34972 6469 35000
rect 5684 34960 5690 34972
rect 6457 34969 6469 34972
rect 6503 34969 6515 35003
rect 6638 35000 6644 35012
rect 6599 34972 6644 35000
rect 6457 34963 6515 34969
rect 6638 34960 6644 34972
rect 6696 34960 6702 35012
rect 5537 34935 5595 34941
rect 5537 34901 5549 34935
rect 5583 34932 5595 34935
rect 6086 34932 6092 34944
rect 5583 34904 6092 34932
rect 5583 34901 5595 34904
rect 5537 34895 5595 34901
rect 6086 34892 6092 34904
rect 6144 34892 6150 34944
rect 6822 34892 6828 34944
rect 6880 34932 6886 34944
rect 7668 34932 7696 35031
rect 9582 35028 9588 35040
rect 9640 35028 9646 35080
rect 10778 35068 10784 35080
rect 10739 35040 10784 35068
rect 10778 35028 10784 35040
rect 10836 35028 10842 35080
rect 10962 35068 10968 35080
rect 10923 35040 10968 35068
rect 10962 35028 10968 35040
rect 11020 35028 11026 35080
rect 11072 35077 11100 35108
rect 11164 35108 11980 35136
rect 11164 35077 11192 35108
rect 11974 35096 11980 35108
rect 12032 35136 12038 35148
rect 16942 35136 16948 35148
rect 12032 35108 16948 35136
rect 12032 35096 12038 35108
rect 16942 35096 16948 35108
rect 17000 35096 17006 35148
rect 11057 35071 11115 35077
rect 11057 35037 11069 35071
rect 11103 35037 11115 35071
rect 11057 35031 11115 35037
rect 11149 35071 11207 35077
rect 11149 35037 11161 35071
rect 11195 35037 11207 35071
rect 11149 35031 11207 35037
rect 11330 35028 11336 35080
rect 11388 35068 11394 35080
rect 12529 35071 12587 35077
rect 12529 35068 12541 35071
rect 11388 35040 12541 35068
rect 11388 35028 11394 35040
rect 12529 35037 12541 35040
rect 12575 35037 12587 35071
rect 12802 35068 12808 35080
rect 12763 35040 12808 35068
rect 12529 35031 12587 35037
rect 12802 35028 12808 35040
rect 12860 35028 12866 35080
rect 12897 35071 12955 35077
rect 12897 35037 12909 35071
rect 12943 35068 12955 35071
rect 12986 35068 12992 35080
rect 12943 35040 12992 35068
rect 12943 35037 12955 35040
rect 12897 35031 12955 35037
rect 12986 35028 12992 35040
rect 13044 35028 13050 35080
rect 11885 35003 11943 35009
rect 11885 35000 11897 35003
rect 10980 34972 11897 35000
rect 10980 34944 11008 34972
rect 11885 34969 11897 34972
rect 11931 34969 11943 35003
rect 11885 34963 11943 34969
rect 12713 35003 12771 35009
rect 12713 34969 12725 35003
rect 12759 35000 12771 35003
rect 13538 35000 13544 35012
rect 12759 34972 13544 35000
rect 12759 34969 12771 34972
rect 12713 34963 12771 34969
rect 6880 34904 7696 34932
rect 6880 34892 6886 34904
rect 10962 34892 10968 34944
rect 11020 34892 11026 34944
rect 11425 34935 11483 34941
rect 11425 34901 11437 34935
rect 11471 34932 11483 34935
rect 11606 34932 11612 34944
rect 11471 34904 11612 34932
rect 11471 34901 11483 34904
rect 11425 34895 11483 34901
rect 11606 34892 11612 34904
rect 11664 34892 11670 34944
rect 12526 34892 12532 34944
rect 12584 34932 12590 34944
rect 12728 34932 12756 34963
rect 13538 34960 13544 34972
rect 13596 34960 13602 35012
rect 12584 34904 12756 34932
rect 13081 34935 13139 34941
rect 12584 34892 12590 34904
rect 13081 34901 13093 34935
rect 13127 34932 13139 34935
rect 14918 34932 14924 34944
rect 13127 34904 14924 34932
rect 13127 34901 13139 34904
rect 13081 34895 13139 34901
rect 14918 34892 14924 34904
rect 14976 34892 14982 34944
rect 17144 34932 17172 35176
rect 22094 35164 22100 35216
rect 22152 35164 22158 35216
rect 25685 35207 25743 35213
rect 25685 35204 25697 35207
rect 24964 35176 25697 35204
rect 20806 35096 20812 35148
rect 20864 35136 20870 35148
rect 22112 35136 22140 35164
rect 20864 35108 22140 35136
rect 20864 35096 20870 35108
rect 17310 35068 17316 35080
rect 17271 35040 17316 35068
rect 17310 35028 17316 35040
rect 17368 35028 17374 35080
rect 21928 35077 21956 35108
rect 20993 35071 21051 35077
rect 20993 35068 21005 35071
rect 18248 35040 21005 35068
rect 18248 35012 18276 35040
rect 20993 35037 21005 35040
rect 21039 35068 21051 35071
rect 21821 35071 21879 35077
rect 21821 35068 21833 35071
rect 21039 35040 21833 35068
rect 21039 35037 21051 35040
rect 20993 35031 21051 35037
rect 21821 35037 21833 35040
rect 21867 35037 21879 35071
rect 21821 35031 21879 35037
rect 21913 35071 21971 35077
rect 21913 35037 21925 35071
rect 21959 35037 21971 35071
rect 21913 35031 21971 35037
rect 22005 35071 22063 35077
rect 22005 35037 22017 35071
rect 22051 35068 22063 35071
rect 22094 35068 22100 35080
rect 22051 35040 22100 35068
rect 22051 35037 22063 35040
rect 22005 35031 22063 35037
rect 22094 35028 22100 35040
rect 22152 35028 22158 35080
rect 22186 35028 22192 35080
rect 22244 35068 22250 35080
rect 22244 35040 22289 35068
rect 22244 35028 22250 35040
rect 23106 35028 23112 35080
rect 23164 35068 23170 35080
rect 24964 35077 24992 35176
rect 25685 35173 25697 35176
rect 25731 35173 25743 35207
rect 25685 35167 25743 35173
rect 32125 35139 32183 35145
rect 32125 35105 32137 35139
rect 32171 35136 32183 35139
rect 32674 35136 32680 35148
rect 32171 35108 32680 35136
rect 32171 35105 32183 35108
rect 32125 35099 32183 35105
rect 24949 35071 25007 35077
rect 24949 35068 24961 35071
rect 23164 35040 24961 35068
rect 23164 35028 23170 35040
rect 24949 35037 24961 35040
rect 24995 35037 25007 35071
rect 24949 35031 25007 35037
rect 27065 35071 27123 35077
rect 27065 35037 27077 35071
rect 27111 35068 27123 35071
rect 27522 35068 27528 35080
rect 27111 35040 27528 35068
rect 27111 35037 27123 35040
rect 27065 35031 27123 35037
rect 27522 35028 27528 35040
rect 27580 35028 27586 35080
rect 30926 35028 30932 35080
rect 30984 35068 30990 35080
rect 31858 35071 31916 35077
rect 31858 35068 31870 35071
rect 30984 35040 31870 35068
rect 30984 35028 30990 35040
rect 31858 35037 31870 35040
rect 31904 35037 31916 35071
rect 31858 35031 31916 35037
rect 32030 35028 32036 35080
rect 32088 35068 32094 35080
rect 32140 35068 32168 35099
rect 32674 35096 32680 35108
rect 32732 35096 32738 35148
rect 58158 35068 58164 35080
rect 32088 35040 32168 35068
rect 58119 35040 58164 35068
rect 32088 35028 32094 35040
rect 58158 35028 58164 35040
rect 58216 35028 58222 35080
rect 17586 35009 17592 35012
rect 17580 34963 17592 35009
rect 17644 35000 17650 35012
rect 17644 34972 17680 35000
rect 17586 34960 17592 34963
rect 17644 34960 17650 34972
rect 18230 34960 18236 35012
rect 18288 34960 18294 35012
rect 18690 34960 18696 35012
rect 18748 35000 18754 35012
rect 21082 35000 21088 35012
rect 18748 34972 21088 35000
rect 18748 34960 18754 34972
rect 21082 34960 21088 34972
rect 21140 34960 21146 35012
rect 24762 35000 24768 35012
rect 24723 34972 24768 35000
rect 24762 34960 24768 34972
rect 24820 34960 24826 35012
rect 25498 34960 25504 35012
rect 25556 35000 25562 35012
rect 26798 35003 26856 35009
rect 26798 35000 26810 35003
rect 25556 34972 26810 35000
rect 25556 34960 25562 34972
rect 26798 34969 26810 34972
rect 26844 34969 26856 35003
rect 29914 35000 29920 35012
rect 29875 34972 29920 35000
rect 26798 34963 26856 34969
rect 29914 34960 29920 34972
rect 29972 34960 29978 35012
rect 30101 35003 30159 35009
rect 30101 34969 30113 35003
rect 30147 35000 30159 35003
rect 30147 34972 30788 35000
rect 30147 34969 30159 34972
rect 30101 34963 30159 34969
rect 19426 34932 19432 34944
rect 17144 34904 19432 34932
rect 19426 34892 19432 34904
rect 19484 34932 19490 34944
rect 19705 34935 19763 34941
rect 19705 34932 19717 34935
rect 19484 34904 19717 34932
rect 19484 34892 19490 34904
rect 19705 34901 19717 34904
rect 19751 34901 19763 34935
rect 21542 34932 21548 34944
rect 21503 34904 21548 34932
rect 19705 34895 19763 34901
rect 21542 34892 21548 34904
rect 21600 34892 21606 34944
rect 25038 34892 25044 34944
rect 25096 34932 25102 34944
rect 30760 34941 30788 34972
rect 25133 34935 25191 34941
rect 25133 34932 25145 34935
rect 25096 34904 25145 34932
rect 25096 34892 25102 34904
rect 25133 34901 25145 34904
rect 25179 34901 25191 34935
rect 25133 34895 25191 34901
rect 30745 34935 30803 34941
rect 30745 34901 30757 34935
rect 30791 34932 30803 34935
rect 31110 34932 31116 34944
rect 30791 34904 31116 34932
rect 30791 34901 30803 34904
rect 30745 34895 30803 34901
rect 31110 34892 31116 34904
rect 31168 34892 31174 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 3881 34731 3939 34737
rect 3881 34697 3893 34731
rect 3927 34697 3939 34731
rect 3881 34691 3939 34697
rect 3896 34660 3924 34691
rect 6638 34688 6644 34740
rect 6696 34728 6702 34740
rect 8478 34728 8484 34740
rect 6696 34700 8484 34728
rect 6696 34688 6702 34700
rect 8478 34688 8484 34700
rect 8536 34688 8542 34740
rect 8757 34731 8815 34737
rect 8757 34697 8769 34731
rect 8803 34728 8815 34731
rect 8846 34728 8852 34740
rect 8803 34700 8852 34728
rect 8803 34697 8815 34700
rect 8757 34691 8815 34697
rect 8846 34688 8852 34700
rect 8904 34688 8910 34740
rect 10318 34728 10324 34740
rect 10279 34700 10324 34728
rect 10318 34688 10324 34700
rect 10376 34688 10382 34740
rect 10686 34688 10692 34740
rect 10744 34688 10750 34740
rect 11698 34688 11704 34740
rect 11756 34728 11762 34740
rect 12897 34731 12955 34737
rect 12897 34728 12909 34731
rect 11756 34700 12909 34728
rect 11756 34688 11762 34700
rect 12897 34697 12909 34700
rect 12943 34697 12955 34731
rect 13722 34728 13728 34740
rect 12897 34691 12955 34697
rect 13648 34700 13728 34728
rect 4525 34663 4583 34669
rect 4525 34660 4537 34663
rect 3896 34632 4537 34660
rect 4525 34629 4537 34632
rect 4571 34660 4583 34663
rect 5074 34660 5080 34672
rect 4571 34632 5080 34660
rect 4571 34629 4583 34632
rect 4525 34623 4583 34629
rect 5074 34620 5080 34632
rect 5132 34620 5138 34672
rect 8294 34660 8300 34672
rect 8128 34632 8300 34660
rect 2498 34592 2504 34604
rect 2459 34564 2504 34592
rect 2498 34552 2504 34564
rect 2556 34552 2562 34604
rect 2774 34601 2780 34604
rect 2768 34555 2780 34601
rect 2832 34592 2838 34604
rect 4709 34595 4767 34601
rect 2832 34564 2868 34592
rect 2774 34552 2780 34555
rect 2832 34552 2838 34564
rect 4709 34561 4721 34595
rect 4755 34592 4767 34595
rect 5626 34592 5632 34604
rect 4755 34564 5632 34592
rect 4755 34561 4767 34564
rect 4709 34555 4767 34561
rect 5626 34552 5632 34564
rect 5684 34552 5690 34604
rect 8128 34601 8156 34632
rect 8294 34620 8300 34632
rect 8352 34620 8358 34672
rect 8389 34663 8447 34669
rect 8389 34629 8401 34663
rect 8435 34660 8447 34663
rect 10410 34660 10416 34672
rect 8435 34632 10416 34660
rect 8435 34629 8447 34632
rect 8389 34623 8447 34629
rect 10410 34620 10416 34632
rect 10468 34620 10474 34672
rect 10704 34607 10732 34688
rect 8113 34595 8171 34601
rect 8113 34561 8125 34595
rect 8159 34561 8171 34595
rect 8113 34555 8171 34561
rect 8202 34552 8208 34604
rect 8260 34592 8266 34604
rect 8260 34564 8305 34592
rect 8260 34552 8266 34564
rect 8478 34552 8484 34604
rect 8536 34592 8542 34604
rect 8619 34595 8677 34601
rect 8536 34564 8578 34592
rect 8536 34552 8542 34564
rect 8619 34561 8631 34595
rect 8665 34592 8677 34595
rect 9674 34592 9680 34604
rect 8665 34564 9680 34592
rect 8665 34561 8677 34564
rect 8619 34555 8677 34561
rect 9674 34552 9680 34564
rect 9732 34552 9738 34604
rect 9769 34595 9827 34601
rect 9769 34561 9781 34595
rect 9815 34592 9827 34595
rect 9950 34592 9956 34604
rect 9815 34564 9956 34592
rect 9815 34561 9827 34564
rect 9769 34555 9827 34561
rect 9950 34552 9956 34564
rect 10008 34592 10014 34604
rect 10226 34592 10232 34604
rect 10008 34564 10232 34592
rect 10008 34552 10014 34564
rect 10226 34552 10232 34564
rect 10284 34552 10290 34604
rect 10686 34601 10744 34607
rect 10551 34595 10609 34601
rect 10551 34592 10563 34595
rect 10541 34561 10563 34592
rect 10597 34561 10609 34595
rect 10686 34567 10698 34601
rect 10732 34567 10744 34601
rect 10686 34561 10744 34567
rect 10541 34555 10609 34561
rect 7558 34484 7564 34536
rect 7616 34524 7622 34536
rect 7653 34527 7711 34533
rect 7653 34524 7665 34527
rect 7616 34496 7665 34524
rect 7616 34484 7622 34496
rect 7653 34493 7665 34496
rect 7699 34524 7711 34527
rect 7742 34524 7748 34536
rect 7699 34496 7748 34524
rect 7699 34493 7711 34496
rect 7653 34487 7711 34493
rect 7742 34484 7748 34496
rect 7800 34484 7806 34536
rect 4982 34416 4988 34468
rect 5040 34456 5046 34468
rect 10541 34456 10569 34555
rect 10778 34552 10784 34604
rect 10836 34601 10842 34604
rect 10836 34592 10844 34601
rect 10836 34564 10881 34592
rect 10836 34555 10844 34564
rect 10836 34552 10842 34555
rect 10962 34552 10968 34604
rect 11020 34592 11026 34604
rect 11020 34564 11065 34592
rect 11020 34552 11026 34564
rect 11606 34552 11612 34604
rect 11664 34592 11670 34604
rect 11773 34595 11831 34601
rect 11773 34592 11785 34595
rect 11664 34564 11785 34592
rect 11664 34552 11670 34564
rect 11773 34561 11785 34564
rect 11819 34561 11831 34595
rect 12912 34592 12940 34691
rect 13538 34660 13544 34672
rect 13499 34632 13544 34660
rect 13538 34620 13544 34632
rect 13596 34620 13602 34672
rect 13648 34669 13676 34700
rect 13722 34688 13728 34700
rect 13780 34688 13786 34740
rect 16942 34728 16948 34740
rect 16903 34700 16948 34728
rect 16942 34688 16948 34700
rect 17000 34688 17006 34740
rect 17497 34731 17555 34737
rect 17497 34697 17509 34731
rect 17543 34728 17555 34731
rect 17586 34728 17592 34740
rect 17543 34700 17592 34728
rect 17543 34697 17555 34700
rect 17497 34691 17555 34697
rect 17586 34688 17592 34700
rect 17644 34688 17650 34740
rect 18322 34728 18328 34740
rect 17972 34700 18328 34728
rect 13633 34663 13691 34669
rect 13633 34629 13645 34663
rect 13679 34629 13691 34663
rect 13633 34623 13691 34629
rect 15470 34620 15476 34672
rect 15528 34660 15534 34672
rect 17972 34660 18000 34700
rect 18322 34688 18328 34700
rect 18380 34728 18386 34740
rect 19429 34731 19487 34737
rect 18380 34700 19104 34728
rect 18380 34688 18386 34700
rect 15528 34632 18000 34660
rect 15528 34620 15534 34632
rect 18046 34620 18052 34672
rect 18104 34660 18110 34672
rect 19076 34669 19104 34700
rect 19429 34697 19441 34731
rect 19475 34728 19487 34731
rect 20162 34728 20168 34740
rect 19475 34700 20168 34728
rect 19475 34697 19487 34700
rect 19429 34691 19487 34697
rect 20162 34688 20168 34700
rect 20220 34688 20226 34740
rect 24670 34728 24676 34740
rect 21008 34700 24676 34728
rect 19061 34663 19119 34669
rect 18104 34632 18920 34660
rect 18104 34620 18110 34632
rect 13357 34595 13415 34601
rect 13357 34592 13369 34595
rect 12912 34564 13369 34592
rect 11773 34555 11831 34561
rect 13357 34561 13369 34564
rect 13403 34561 13415 34595
rect 13357 34555 13415 34561
rect 13725 34595 13783 34601
rect 13725 34561 13737 34595
rect 13771 34561 13783 34595
rect 13725 34555 13783 34561
rect 11422 34484 11428 34536
rect 11480 34524 11486 34536
rect 11517 34527 11575 34533
rect 11517 34524 11529 34527
rect 11480 34496 11529 34524
rect 11480 34484 11486 34496
rect 11517 34493 11529 34496
rect 11563 34493 11575 34527
rect 11517 34487 11575 34493
rect 12986 34484 12992 34536
rect 13044 34524 13050 34536
rect 13740 34524 13768 34555
rect 16942 34552 16948 34604
rect 17000 34592 17006 34604
rect 17727 34595 17785 34601
rect 17727 34592 17739 34595
rect 17000 34564 17739 34592
rect 17000 34552 17006 34564
rect 17727 34561 17739 34564
rect 17773 34561 17785 34595
rect 17862 34592 17868 34604
rect 17823 34564 17868 34592
rect 17727 34555 17785 34561
rect 17862 34552 17868 34564
rect 17920 34552 17926 34604
rect 17954 34552 17960 34604
rect 18012 34592 18018 34604
rect 18012 34564 18057 34592
rect 18012 34552 18018 34564
rect 18138 34552 18144 34604
rect 18196 34592 18202 34604
rect 18892 34601 18920 34632
rect 19061 34629 19073 34663
rect 19107 34629 19119 34663
rect 19061 34623 19119 34629
rect 19153 34663 19211 34669
rect 19153 34629 19165 34663
rect 19199 34660 19211 34663
rect 19794 34660 19800 34672
rect 19199 34632 19800 34660
rect 19199 34629 19211 34632
rect 19153 34623 19211 34629
rect 19794 34620 19800 34632
rect 19852 34620 19858 34672
rect 18785 34595 18843 34601
rect 18196 34564 18241 34592
rect 18196 34552 18202 34564
rect 18785 34561 18797 34595
rect 18831 34561 18843 34595
rect 18785 34555 18843 34561
rect 18878 34595 18936 34601
rect 18878 34561 18890 34595
rect 18924 34561 18936 34595
rect 18878 34555 18936 34561
rect 18800 34524 18828 34555
rect 19242 34552 19248 34604
rect 19300 34601 19306 34604
rect 19300 34592 19308 34601
rect 19300 34564 19345 34592
rect 19300 34555 19308 34564
rect 19300 34552 19306 34555
rect 19518 34552 19524 34604
rect 19576 34592 19582 34604
rect 19889 34595 19947 34601
rect 19889 34592 19901 34595
rect 19576 34564 19901 34592
rect 19576 34552 19582 34564
rect 19889 34561 19901 34564
rect 19935 34561 19947 34595
rect 20070 34592 20076 34604
rect 20031 34564 20076 34592
rect 19889 34555 19947 34561
rect 20070 34552 20076 34564
rect 20128 34552 20134 34604
rect 20165 34595 20223 34601
rect 20165 34561 20177 34595
rect 20211 34561 20223 34595
rect 20165 34555 20223 34561
rect 13044 34496 13768 34524
rect 13924 34496 18828 34524
rect 13044 34484 13050 34496
rect 11238 34456 11244 34468
rect 5040 34428 5534 34456
rect 10541 34428 11244 34456
rect 5040 34416 5046 34428
rect 3142 34348 3148 34400
rect 3200 34388 3206 34400
rect 4341 34391 4399 34397
rect 4341 34388 4353 34391
rect 3200 34360 4353 34388
rect 3200 34348 3206 34360
rect 4341 34357 4353 34360
rect 4387 34357 4399 34391
rect 5506 34388 5534 34428
rect 11238 34416 11244 34428
rect 11296 34416 11302 34468
rect 13924 34465 13952 34496
rect 19426 34484 19432 34536
rect 19484 34524 19490 34536
rect 20180 34524 20208 34555
rect 20254 34552 20260 34604
rect 20312 34592 20318 34604
rect 21008 34601 21036 34700
rect 24670 34688 24676 34700
rect 24728 34688 24734 34740
rect 25498 34728 25504 34740
rect 25459 34700 25504 34728
rect 25498 34688 25504 34700
rect 25556 34688 25562 34740
rect 32309 34731 32367 34737
rect 32309 34697 32321 34731
rect 32355 34728 32367 34731
rect 33778 34728 33784 34740
rect 32355 34700 33784 34728
rect 32355 34697 32367 34700
rect 32309 34691 32367 34697
rect 33778 34688 33784 34700
rect 33836 34688 33842 34740
rect 21542 34620 21548 34672
rect 21600 34660 21606 34672
rect 22066 34663 22124 34669
rect 22066 34660 22078 34663
rect 21600 34632 22078 34660
rect 21600 34620 21606 34632
rect 22066 34629 22078 34632
rect 22112 34629 22124 34663
rect 22066 34623 22124 34629
rect 24946 34620 24952 34672
rect 25004 34660 25010 34672
rect 25004 34632 25176 34660
rect 25004 34620 25010 34632
rect 20993 34595 21051 34601
rect 20993 34592 21005 34595
rect 20312 34564 21005 34592
rect 20312 34552 20318 34564
rect 20993 34561 21005 34564
rect 21039 34561 21051 34595
rect 20993 34555 21051 34561
rect 21821 34595 21879 34601
rect 21821 34561 21833 34595
rect 21867 34592 21879 34595
rect 21910 34592 21916 34604
rect 21867 34564 21916 34592
rect 21867 34561 21879 34564
rect 21821 34555 21879 34561
rect 21910 34552 21916 34564
rect 21968 34552 21974 34604
rect 24394 34552 24400 34604
rect 24452 34592 24458 34604
rect 24857 34595 24915 34601
rect 24857 34592 24869 34595
rect 24452 34564 24869 34592
rect 24452 34552 24458 34564
rect 24857 34561 24869 34564
rect 24903 34561 24915 34595
rect 25038 34592 25044 34604
rect 24999 34564 25044 34592
rect 24857 34555 24915 34561
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 25148 34601 25176 34632
rect 30098 34620 30104 34672
rect 30156 34660 30162 34672
rect 34517 34663 34575 34669
rect 34517 34660 34529 34663
rect 30156 34632 34529 34660
rect 30156 34620 30162 34632
rect 34517 34629 34529 34632
rect 34563 34660 34575 34663
rect 35710 34660 35716 34672
rect 34563 34632 35716 34660
rect 34563 34629 34575 34632
rect 34517 34623 34575 34629
rect 35710 34620 35716 34632
rect 35768 34620 35774 34672
rect 25133 34595 25191 34601
rect 25133 34561 25145 34595
rect 25179 34561 25191 34595
rect 25133 34555 25191 34561
rect 25222 34552 25228 34604
rect 25280 34592 25286 34604
rect 25961 34595 26019 34601
rect 25961 34592 25973 34595
rect 25280 34564 25973 34592
rect 25280 34552 25286 34564
rect 25961 34561 25973 34564
rect 26007 34592 26019 34595
rect 26050 34592 26056 34604
rect 26007 34564 26056 34592
rect 26007 34561 26019 34564
rect 25961 34555 26019 34561
rect 26050 34552 26056 34564
rect 26108 34552 26114 34604
rect 30650 34592 30656 34604
rect 29748 34564 30656 34592
rect 20438 34524 20444 34536
rect 19484 34496 20444 34524
rect 19484 34484 19490 34496
rect 20438 34484 20444 34496
rect 20496 34484 20502 34536
rect 20533 34527 20591 34533
rect 20533 34493 20545 34527
rect 20579 34524 20591 34527
rect 21542 34524 21548 34536
rect 20579 34496 21548 34524
rect 20579 34493 20591 34496
rect 20533 34487 20591 34493
rect 21542 34484 21548 34496
rect 21600 34484 21606 34536
rect 29638 34484 29644 34536
rect 29696 34524 29702 34536
rect 29748 34533 29776 34564
rect 30650 34552 30656 34564
rect 30708 34592 30714 34604
rect 31113 34595 31171 34601
rect 31113 34592 31125 34595
rect 30708 34564 31125 34592
rect 30708 34552 30714 34564
rect 31113 34561 31125 34564
rect 31159 34561 31171 34595
rect 31113 34555 31171 34561
rect 31754 34552 31760 34604
rect 31812 34592 31818 34604
rect 32125 34595 32183 34601
rect 32125 34592 32137 34595
rect 31812 34564 32137 34592
rect 31812 34552 31818 34564
rect 32125 34561 32137 34564
rect 32171 34561 32183 34595
rect 32125 34555 32183 34561
rect 29733 34527 29791 34533
rect 29733 34524 29745 34527
rect 29696 34496 29745 34524
rect 29696 34484 29702 34496
rect 29733 34493 29745 34496
rect 29779 34493 29791 34527
rect 29733 34487 29791 34493
rect 30190 34484 30196 34536
rect 30248 34524 30254 34536
rect 30837 34527 30895 34533
rect 30837 34524 30849 34527
rect 30248 34496 30849 34524
rect 30248 34484 30254 34496
rect 30837 34493 30849 34496
rect 30883 34493 30895 34527
rect 30837 34487 30895 34493
rect 13909 34459 13967 34465
rect 13909 34425 13921 34459
rect 13955 34425 13967 34459
rect 27154 34456 27160 34468
rect 13909 34419 13967 34425
rect 16868 34428 21128 34456
rect 9677 34391 9735 34397
rect 9677 34388 9689 34391
rect 5506 34360 9689 34388
rect 4341 34351 4399 34357
rect 9677 34357 9689 34360
rect 9723 34388 9735 34391
rect 9858 34388 9864 34400
rect 9723 34360 9864 34388
rect 9723 34357 9735 34360
rect 9677 34351 9735 34357
rect 9858 34348 9864 34360
rect 9916 34348 9922 34400
rect 11698 34348 11704 34400
rect 11756 34388 11762 34400
rect 16868 34388 16896 34428
rect 11756 34360 16896 34388
rect 21100 34388 21128 34428
rect 22756 34428 27160 34456
rect 22756 34388 22784 34428
rect 27154 34416 27160 34428
rect 27212 34416 27218 34468
rect 21100 34360 22784 34388
rect 11756 34348 11762 34360
rect 22830 34348 22836 34400
rect 22888 34388 22894 34400
rect 23201 34391 23259 34397
rect 23201 34388 23213 34391
rect 22888 34360 23213 34388
rect 22888 34348 22894 34360
rect 23201 34357 23213 34360
rect 23247 34357 23259 34391
rect 23201 34351 23259 34357
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 2593 34187 2651 34193
rect 2593 34153 2605 34187
rect 2639 34184 2651 34187
rect 2774 34184 2780 34196
rect 2639 34156 2780 34184
rect 2639 34153 2651 34156
rect 2593 34147 2651 34153
rect 2774 34144 2780 34156
rect 2832 34144 2838 34196
rect 7374 34144 7380 34196
rect 7432 34184 7438 34196
rect 9401 34187 9459 34193
rect 9401 34184 9413 34187
rect 7432 34156 9413 34184
rect 7432 34144 7438 34156
rect 9401 34153 9413 34156
rect 9447 34153 9459 34187
rect 9401 34147 9459 34153
rect 10778 34144 10784 34196
rect 10836 34184 10842 34196
rect 10965 34187 11023 34193
rect 10965 34184 10977 34187
rect 10836 34156 10977 34184
rect 10836 34144 10842 34156
rect 10965 34153 10977 34156
rect 11011 34153 11023 34187
rect 10965 34147 11023 34153
rect 11238 34144 11244 34196
rect 11296 34184 11302 34196
rect 11425 34187 11483 34193
rect 11425 34184 11437 34187
rect 11296 34156 11437 34184
rect 11296 34144 11302 34156
rect 11425 34153 11437 34156
rect 11471 34153 11483 34187
rect 11974 34184 11980 34196
rect 11935 34156 11980 34184
rect 11425 34147 11483 34153
rect 11974 34144 11980 34156
rect 12032 34144 12038 34196
rect 14366 34144 14372 34196
rect 14424 34184 14430 34196
rect 15013 34187 15071 34193
rect 15013 34184 15025 34187
rect 14424 34156 15025 34184
rect 14424 34144 14430 34156
rect 15013 34153 15025 34156
rect 15059 34184 15071 34187
rect 17862 34184 17868 34196
rect 15059 34156 17868 34184
rect 15059 34153 15071 34156
rect 15013 34147 15071 34153
rect 6822 34116 6828 34128
rect 2976 34088 6828 34116
rect 2866 33980 2872 33992
rect 2827 33952 2872 33980
rect 2866 33940 2872 33952
rect 2924 33940 2930 33992
rect 2976 33989 3004 34088
rect 2961 33983 3019 33989
rect 2961 33949 2973 33983
rect 3007 33949 3019 33983
rect 2961 33943 3019 33949
rect 3053 33983 3111 33989
rect 3053 33949 3065 33983
rect 3099 33980 3111 33983
rect 3142 33980 3148 33992
rect 3099 33952 3148 33980
rect 3099 33949 3111 33952
rect 3053 33943 3111 33949
rect 3142 33940 3148 33952
rect 3200 33940 3206 33992
rect 3237 33983 3295 33989
rect 3237 33949 3249 33983
rect 3283 33949 3295 33983
rect 4062 33980 4068 33992
rect 4023 33952 4068 33980
rect 3237 33943 3295 33949
rect 2133 33915 2191 33921
rect 2133 33881 2145 33915
rect 2179 33912 2191 33915
rect 2884 33912 2912 33940
rect 2179 33884 2912 33912
rect 3252 33912 3280 33943
rect 4062 33940 4068 33952
rect 4120 33940 4126 33992
rect 4172 33989 4200 34088
rect 6822 34076 6828 34088
rect 6880 34076 6886 34128
rect 9674 34076 9680 34128
rect 9732 34116 9738 34128
rect 14093 34119 14151 34125
rect 14093 34116 14105 34119
rect 9732 34088 14105 34116
rect 9732 34076 9738 34088
rect 14093 34085 14105 34088
rect 14139 34085 14151 34119
rect 14093 34079 14151 34085
rect 5537 34051 5595 34057
rect 5537 34017 5549 34051
rect 5583 34048 5595 34051
rect 11698 34048 11704 34060
rect 5583 34020 11704 34048
rect 5583 34017 5595 34020
rect 5537 34011 5595 34017
rect 4157 33983 4215 33989
rect 4157 33949 4169 33983
rect 4203 33949 4215 33983
rect 4157 33943 4215 33949
rect 4249 33983 4307 33989
rect 4249 33949 4261 33983
rect 4295 33980 4307 33983
rect 4338 33980 4344 33992
rect 4295 33952 4344 33980
rect 4295 33949 4307 33952
rect 4249 33943 4307 33949
rect 4338 33940 4344 33952
rect 4396 33940 4402 33992
rect 4433 33983 4491 33989
rect 4433 33949 4445 33983
rect 4479 33949 4491 33983
rect 4433 33943 4491 33949
rect 4448 33912 4476 33943
rect 4893 33915 4951 33921
rect 4893 33912 4905 33915
rect 3252 33884 4905 33912
rect 2179 33881 2191 33884
rect 2133 33875 2191 33881
rect 4080 33856 4108 33884
rect 4893 33881 4905 33884
rect 4939 33881 4951 33915
rect 4893 33875 4951 33881
rect 3786 33844 3792 33856
rect 3747 33816 3792 33844
rect 3786 33804 3792 33816
rect 3844 33804 3850 33856
rect 4062 33804 4068 33856
rect 4120 33804 4126 33856
rect 4154 33804 4160 33856
rect 4212 33844 4218 33856
rect 5552 33844 5580 34011
rect 11698 34008 11704 34020
rect 11756 34008 11762 34060
rect 10781 33983 10839 33989
rect 10781 33949 10793 33983
rect 10827 33980 10839 33983
rect 11330 33980 11336 33992
rect 10827 33952 11336 33980
rect 10827 33949 10839 33952
rect 10781 33943 10839 33949
rect 11330 33940 11336 33952
rect 11388 33940 11394 33992
rect 9493 33915 9551 33921
rect 9493 33881 9505 33915
rect 9539 33912 9551 33915
rect 9582 33912 9588 33924
rect 9539 33884 9588 33912
rect 9539 33881 9551 33884
rect 9493 33875 9551 33881
rect 9582 33872 9588 33884
rect 9640 33872 9646 33924
rect 10597 33915 10655 33921
rect 10597 33881 10609 33915
rect 10643 33912 10655 33915
rect 11054 33912 11060 33924
rect 10643 33884 11060 33912
rect 10643 33881 10655 33884
rect 10597 33875 10655 33881
rect 11054 33872 11060 33884
rect 11112 33872 11118 33924
rect 5718 33844 5724 33856
rect 4212 33816 5724 33844
rect 4212 33804 4218 33816
rect 5718 33804 5724 33816
rect 5776 33804 5782 33856
rect 14108 33844 14136 34079
rect 16945 34051 17003 34057
rect 16945 34017 16957 34051
rect 16991 34048 17003 34051
rect 17310 34048 17316 34060
rect 16991 34020 17316 34048
rect 16991 34017 17003 34020
rect 16945 34011 17003 34017
rect 17310 34008 17316 34020
rect 17368 34008 17374 34060
rect 14277 33983 14335 33989
rect 14277 33949 14289 33983
rect 14323 33980 14335 33983
rect 16390 33980 16396 33992
rect 14323 33952 16396 33980
rect 14323 33949 14335 33952
rect 14277 33943 14335 33949
rect 16390 33940 16396 33952
rect 16448 33940 16454 33992
rect 17586 33940 17592 33992
rect 17644 33980 17650 33992
rect 17788 33989 17816 34156
rect 17862 34144 17868 34156
rect 17920 34144 17926 34196
rect 20070 34184 20076 34196
rect 20031 34156 20076 34184
rect 20070 34144 20076 34156
rect 20128 34144 20134 34196
rect 22094 34144 22100 34196
rect 22152 34184 22158 34196
rect 22557 34187 22615 34193
rect 22557 34184 22569 34187
rect 22152 34156 22569 34184
rect 22152 34144 22158 34156
rect 22557 34153 22569 34156
rect 22603 34153 22615 34187
rect 22557 34147 22615 34153
rect 27157 34187 27215 34193
rect 27157 34153 27169 34187
rect 27203 34184 27215 34187
rect 27890 34184 27896 34196
rect 27203 34156 27896 34184
rect 27203 34153 27215 34156
rect 27157 34147 27215 34153
rect 27890 34144 27896 34156
rect 27948 34184 27954 34196
rect 28350 34184 28356 34196
rect 27948 34156 28356 34184
rect 27948 34144 27954 34156
rect 28350 34144 28356 34156
rect 28408 34144 28414 34196
rect 20717 34119 20775 34125
rect 20717 34116 20729 34119
rect 19904 34088 20729 34116
rect 17681 33983 17739 33989
rect 17681 33980 17693 33983
rect 17644 33952 17693 33980
rect 17644 33940 17650 33952
rect 17681 33949 17693 33952
rect 17727 33949 17739 33983
rect 17681 33943 17739 33949
rect 17773 33983 17831 33989
rect 17773 33949 17785 33983
rect 17819 33949 17831 33983
rect 17773 33943 17831 33949
rect 17862 33940 17868 33992
rect 17920 33980 17926 33992
rect 18049 33983 18107 33989
rect 17920 33952 17965 33980
rect 17920 33940 17926 33952
rect 18049 33949 18061 33983
rect 18095 33980 18107 33983
rect 18138 33980 18144 33992
rect 18095 33952 18144 33980
rect 18095 33949 18107 33952
rect 18049 33943 18107 33949
rect 18138 33940 18144 33952
rect 18196 33940 18202 33992
rect 19334 33940 19340 33992
rect 19392 33980 19398 33992
rect 19705 33983 19763 33989
rect 19705 33980 19717 33983
rect 19392 33952 19717 33980
rect 19392 33940 19398 33952
rect 19705 33949 19717 33952
rect 19751 33949 19763 33983
rect 19705 33943 19763 33949
rect 19794 33940 19800 33992
rect 19852 33980 19858 33992
rect 19904 33989 19932 34088
rect 20717 34085 20729 34088
rect 20763 34085 20775 34119
rect 20717 34079 20775 34085
rect 24946 34048 24952 34060
rect 24688 34020 24952 34048
rect 19889 33983 19947 33989
rect 19889 33980 19901 33983
rect 19852 33952 19901 33980
rect 19852 33940 19858 33952
rect 19889 33949 19901 33952
rect 19935 33949 19947 33983
rect 19889 33943 19947 33949
rect 21542 33940 21548 33992
rect 21600 33980 21606 33992
rect 21830 33983 21888 33989
rect 21830 33980 21842 33983
rect 21600 33952 21842 33980
rect 21600 33940 21606 33952
rect 21830 33949 21842 33952
rect 21876 33949 21888 33983
rect 21830 33943 21888 33949
rect 22002 33940 22008 33992
rect 22060 33980 22066 33992
rect 22097 33983 22155 33989
rect 22097 33980 22109 33983
rect 22060 33952 22109 33980
rect 22060 33940 22066 33952
rect 22097 33949 22109 33952
rect 22143 33949 22155 33983
rect 24394 33980 24400 33992
rect 24355 33952 24400 33980
rect 22097 33943 22155 33949
rect 24394 33940 24400 33952
rect 24452 33940 24458 33992
rect 24578 33980 24584 33992
rect 24539 33952 24584 33980
rect 24578 33940 24584 33952
rect 24636 33940 24642 33992
rect 24688 33989 24716 34020
rect 24946 34008 24952 34020
rect 25004 34008 25010 34060
rect 30653 34051 30711 34057
rect 30653 34017 30665 34051
rect 30699 34048 30711 34051
rect 30699 34020 31754 34048
rect 30699 34017 30711 34020
rect 30653 34011 30711 34017
rect 31726 33992 31754 34020
rect 33594 34008 33600 34060
rect 33652 34048 33658 34060
rect 33652 34020 34744 34048
rect 33652 34008 33658 34020
rect 24673 33983 24731 33989
rect 24673 33949 24685 33983
rect 24719 33949 24731 33983
rect 24673 33943 24731 33949
rect 24765 33983 24823 33989
rect 24765 33949 24777 33983
rect 24811 33949 24823 33983
rect 24765 33943 24823 33949
rect 14366 33872 14372 33924
rect 14424 33912 14430 33924
rect 14921 33915 14979 33921
rect 14921 33912 14933 33915
rect 14424 33884 14933 33912
rect 14424 33872 14430 33884
rect 14921 33881 14933 33884
rect 14967 33881 14979 33915
rect 16700 33915 16758 33921
rect 14921 33875 14979 33881
rect 15396 33884 16620 33912
rect 15396 33844 15424 33884
rect 15562 33844 15568 33856
rect 14108 33816 15424 33844
rect 15523 33816 15568 33844
rect 15562 33804 15568 33816
rect 15620 33804 15626 33856
rect 16592 33844 16620 33884
rect 16700 33881 16712 33915
rect 16746 33912 16758 33915
rect 17405 33915 17463 33921
rect 17405 33912 17417 33915
rect 16746 33884 17417 33912
rect 16746 33881 16758 33884
rect 16700 33875 16758 33881
rect 17405 33881 17417 33884
rect 17451 33881 17463 33915
rect 17405 33875 17463 33881
rect 19058 33872 19064 33924
rect 19116 33912 19122 33924
rect 19518 33912 19524 33924
rect 19116 33884 19524 33912
rect 19116 33872 19122 33884
rect 19518 33872 19524 33884
rect 19576 33872 19582 33924
rect 22738 33912 22744 33924
rect 22699 33884 22744 33912
rect 22738 33872 22744 33884
rect 22796 33872 22802 33924
rect 22925 33915 22983 33921
rect 22925 33881 22937 33915
rect 22971 33912 22983 33915
rect 23290 33912 23296 33924
rect 22971 33884 23296 33912
rect 22971 33881 22983 33884
rect 22925 33875 22983 33881
rect 18506 33844 18512 33856
rect 16592 33816 18512 33844
rect 18506 33804 18512 33816
rect 18564 33844 18570 33856
rect 19242 33844 19248 33856
rect 18564 33816 19248 33844
rect 18564 33804 18570 33816
rect 19242 33804 19248 33816
rect 19300 33804 19306 33856
rect 22094 33804 22100 33856
rect 22152 33844 22158 33856
rect 22940 33844 22968 33875
rect 23290 33872 23296 33884
rect 23348 33872 23354 33924
rect 23750 33872 23756 33924
rect 23808 33912 23814 33924
rect 23845 33915 23903 33921
rect 23845 33912 23857 33915
rect 23808 33884 23857 33912
rect 23808 33872 23814 33884
rect 23845 33881 23857 33884
rect 23891 33912 23903 33915
rect 24780 33912 24808 33943
rect 27522 33940 27528 33992
rect 27580 33980 27586 33992
rect 27617 33983 27675 33989
rect 27617 33980 27629 33983
rect 27580 33952 27629 33980
rect 27580 33940 27586 33952
rect 27617 33949 27629 33952
rect 27663 33949 27675 33983
rect 27617 33943 27675 33949
rect 29825 33983 29883 33989
rect 29825 33949 29837 33983
rect 29871 33980 29883 33983
rect 29914 33980 29920 33992
rect 29871 33952 29920 33980
rect 29871 33949 29883 33952
rect 29825 33943 29883 33949
rect 29914 33940 29920 33952
rect 29972 33980 29978 33992
rect 30098 33980 30104 33992
rect 29972 33952 30104 33980
rect 29972 33940 29978 33952
rect 30098 33940 30104 33952
rect 30156 33940 30162 33992
rect 30742 33940 30748 33992
rect 30800 33980 30806 33992
rect 30929 33983 30987 33989
rect 30929 33980 30941 33983
rect 30800 33952 30941 33980
rect 30800 33940 30806 33952
rect 30929 33949 30941 33952
rect 30975 33949 30987 33983
rect 31726 33952 31760 33992
rect 30929 33943 30987 33949
rect 31754 33940 31760 33952
rect 31812 33940 31818 33992
rect 31941 33983 31999 33989
rect 31941 33949 31953 33983
rect 31987 33980 31999 33983
rect 32030 33980 32036 33992
rect 31987 33952 32036 33980
rect 31987 33949 31999 33952
rect 31941 33943 31999 33949
rect 32030 33940 32036 33952
rect 32088 33940 32094 33992
rect 33778 33980 33784 33992
rect 33739 33952 33784 33980
rect 33778 33940 33784 33952
rect 33836 33940 33842 33992
rect 33965 33983 34023 33989
rect 33965 33949 33977 33983
rect 34011 33980 34023 33983
rect 34606 33980 34612 33992
rect 34011 33952 34612 33980
rect 34011 33949 34023 33952
rect 33965 33943 34023 33949
rect 34606 33940 34612 33952
rect 34664 33940 34670 33992
rect 34716 33989 34744 34020
rect 34701 33983 34759 33989
rect 34701 33949 34713 33983
rect 34747 33949 34759 33983
rect 34864 33983 34922 33989
rect 34864 33980 34876 33983
rect 34701 33943 34759 33949
rect 34808 33952 34876 33980
rect 23891 33884 24808 33912
rect 23891 33881 23903 33884
rect 23845 33875 23903 33881
rect 27706 33872 27712 33924
rect 27764 33912 27770 33924
rect 27862 33915 27920 33921
rect 27862 33912 27874 33915
rect 27764 33884 27874 33912
rect 27764 33872 27770 33884
rect 27862 33881 27874 33884
rect 27908 33881 27920 33915
rect 30006 33912 30012 33924
rect 29967 33884 30012 33912
rect 27862 33875 27920 33881
rect 30006 33872 30012 33884
rect 30064 33872 30070 33924
rect 32214 33921 32220 33924
rect 32208 33875 32220 33921
rect 32272 33912 32278 33924
rect 34149 33915 34207 33921
rect 32272 33884 32308 33912
rect 32214 33872 32220 33875
rect 32272 33872 32278 33884
rect 34149 33881 34161 33915
rect 34195 33912 34207 33915
rect 34808 33912 34836 33952
rect 34864 33949 34876 33952
rect 34910 33949 34922 33983
rect 34864 33943 34922 33949
rect 34964 33980 35022 33986
rect 34964 33946 34976 33980
rect 35010 33977 35022 33980
rect 35115 33983 35173 33989
rect 35010 33946 35023 33977
rect 34964 33940 35023 33946
rect 35115 33949 35127 33983
rect 35161 33980 35173 33983
rect 35710 33980 35716 33992
rect 35161 33952 35716 33980
rect 35161 33949 35173 33952
rect 35115 33943 35173 33949
rect 35710 33940 35716 33952
rect 35768 33940 35774 33992
rect 34195 33884 34836 33912
rect 34195 33881 34207 33884
rect 34149 33875 34207 33881
rect 34995 33856 35023 33940
rect 25038 33844 25044 33856
rect 22152 33816 22968 33844
rect 24999 33816 25044 33844
rect 22152 33804 22158 33816
rect 25038 33804 25044 33816
rect 25096 33804 25102 33856
rect 28997 33847 29055 33853
rect 28997 33813 29009 33847
rect 29043 33844 29055 33847
rect 29086 33844 29092 33856
rect 29043 33816 29092 33844
rect 29043 33813 29055 33816
rect 28997 33807 29055 33813
rect 29086 33804 29092 33816
rect 29144 33804 29150 33856
rect 30193 33847 30251 33853
rect 30193 33813 30205 33847
rect 30239 33844 30251 33847
rect 30466 33844 30472 33856
rect 30239 33816 30472 33844
rect 30239 33813 30251 33816
rect 30193 33807 30251 33813
rect 30466 33804 30472 33816
rect 30524 33804 30530 33856
rect 33318 33844 33324 33856
rect 33279 33816 33324 33844
rect 33318 33804 33324 33816
rect 33376 33804 33382 33856
rect 34974 33804 34980 33856
rect 35032 33804 35038 33856
rect 35345 33847 35403 33853
rect 35345 33813 35357 33847
rect 35391 33844 35403 33847
rect 35986 33844 35992 33856
rect 35391 33816 35992 33844
rect 35391 33813 35403 33816
rect 35345 33807 35403 33813
rect 35986 33804 35992 33816
rect 36044 33804 36050 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 4338 33640 4344 33652
rect 4299 33612 4344 33640
rect 4338 33600 4344 33612
rect 4396 33600 4402 33652
rect 8202 33640 8208 33652
rect 8163 33612 8208 33640
rect 8202 33600 8208 33612
rect 8260 33600 8266 33652
rect 11238 33600 11244 33652
rect 11296 33640 11302 33652
rect 17037 33643 17095 33649
rect 11296 33612 16988 33640
rect 11296 33600 11302 33612
rect 6362 33572 6368 33584
rect 2516 33544 6368 33572
rect 2222 33396 2228 33448
rect 2280 33436 2286 33448
rect 2516 33445 2544 33544
rect 6362 33532 6368 33544
rect 6420 33572 6426 33584
rect 6420 33544 6868 33572
rect 6420 33532 6426 33544
rect 2768 33507 2826 33513
rect 2768 33473 2780 33507
rect 2814 33504 2826 33507
rect 3786 33504 3792 33516
rect 2814 33476 3792 33504
rect 2814 33473 2826 33476
rect 2768 33467 2826 33473
rect 3786 33464 3792 33476
rect 3844 33464 3850 33516
rect 4525 33507 4583 33513
rect 4525 33473 4537 33507
rect 4571 33473 4583 33507
rect 4525 33467 4583 33473
rect 4709 33507 4767 33513
rect 4709 33473 4721 33507
rect 4755 33504 4767 33507
rect 5626 33504 5632 33516
rect 4755 33476 5632 33504
rect 4755 33473 4767 33476
rect 4709 33467 4767 33473
rect 2501 33439 2559 33445
rect 2501 33436 2513 33439
rect 2280 33408 2513 33436
rect 2280 33396 2286 33408
rect 2501 33405 2513 33408
rect 2547 33405 2559 33439
rect 4540 33436 4568 33467
rect 5626 33464 5632 33476
rect 5684 33464 5690 33516
rect 6840 33513 6868 33544
rect 10410 33532 10416 33584
rect 10468 33572 10474 33584
rect 12713 33575 12771 33581
rect 12713 33572 12725 33575
rect 10468 33544 12725 33572
rect 10468 33532 10474 33544
rect 12713 33541 12725 33544
rect 12759 33572 12771 33575
rect 15470 33572 15476 33584
rect 12759 33544 15476 33572
rect 12759 33541 12771 33544
rect 12713 33535 12771 33541
rect 15470 33532 15476 33544
rect 15528 33532 15534 33584
rect 15562 33532 15568 33584
rect 15620 33572 15626 33584
rect 16298 33572 16304 33584
rect 15620 33544 16304 33572
rect 15620 33532 15626 33544
rect 16298 33532 16304 33544
rect 16356 33572 16362 33584
rect 16853 33575 16911 33581
rect 16853 33572 16865 33575
rect 16356 33544 16865 33572
rect 16356 33532 16362 33544
rect 16853 33541 16865 33544
rect 16899 33541 16911 33575
rect 16960 33572 16988 33612
rect 17037 33609 17049 33643
rect 17083 33640 17095 33643
rect 17862 33640 17868 33652
rect 17083 33612 17868 33640
rect 17083 33609 17095 33612
rect 17037 33603 17095 33609
rect 17862 33600 17868 33612
rect 17920 33600 17926 33652
rect 19058 33640 19064 33652
rect 19019 33612 19064 33640
rect 19058 33600 19064 33612
rect 19116 33600 19122 33652
rect 24762 33640 24768 33652
rect 23584 33612 24768 33640
rect 17497 33575 17555 33581
rect 17497 33572 17509 33575
rect 16960 33544 17509 33572
rect 16853 33535 16911 33541
rect 17497 33541 17509 33544
rect 17543 33572 17555 33575
rect 17586 33572 17592 33584
rect 17543 33544 17592 33572
rect 17543 33541 17555 33544
rect 17497 33535 17555 33541
rect 17586 33532 17592 33544
rect 17644 33532 17650 33584
rect 18325 33575 18383 33581
rect 18325 33541 18337 33575
rect 18371 33572 18383 33575
rect 18598 33572 18604 33584
rect 18371 33544 18604 33572
rect 18371 33541 18383 33544
rect 18325 33535 18383 33541
rect 18598 33532 18604 33544
rect 18656 33532 18662 33584
rect 19334 33572 19340 33584
rect 18800 33544 19340 33572
rect 6825 33507 6883 33513
rect 6825 33473 6837 33507
rect 6871 33473 6883 33507
rect 6825 33467 6883 33473
rect 6914 33464 6920 33516
rect 6972 33504 6978 33516
rect 7081 33507 7139 33513
rect 7081 33504 7093 33507
rect 6972 33476 7093 33504
rect 6972 33464 6978 33476
rect 7081 33473 7093 33476
rect 7127 33473 7139 33507
rect 7081 33467 7139 33473
rect 12342 33464 12348 33516
rect 12400 33504 12406 33516
rect 12897 33507 12955 33513
rect 12897 33504 12909 33507
rect 12400 33476 12909 33504
rect 12400 33464 12406 33476
rect 12897 33473 12909 33476
rect 12943 33504 12955 33507
rect 16482 33504 16488 33516
rect 12943 33476 16488 33504
rect 12943 33473 12955 33476
rect 12897 33467 12955 33473
rect 16482 33464 16488 33476
rect 16540 33464 16546 33516
rect 16669 33507 16727 33513
rect 16669 33473 16681 33507
rect 16715 33473 16727 33507
rect 16669 33467 16727 33473
rect 5350 33436 5356 33448
rect 2501 33399 2559 33405
rect 3896 33408 5356 33436
rect 3896 33377 3924 33408
rect 5350 33396 5356 33408
rect 5408 33396 5414 33448
rect 14550 33436 14556 33448
rect 14511 33408 14556 33436
rect 14550 33396 14556 33408
rect 14608 33396 14614 33448
rect 14829 33439 14887 33445
rect 14829 33405 14841 33439
rect 14875 33436 14887 33439
rect 15654 33436 15660 33448
rect 14875 33408 15660 33436
rect 14875 33405 14887 33408
rect 14829 33399 14887 33405
rect 15654 33396 15660 33408
rect 15712 33436 15718 33448
rect 16684 33436 16712 33467
rect 17954 33464 17960 33516
rect 18012 33504 18018 33516
rect 18509 33507 18567 33513
rect 18509 33504 18521 33507
rect 18012 33476 18521 33504
rect 18012 33464 18018 33476
rect 18509 33473 18521 33476
rect 18555 33504 18567 33507
rect 18800 33504 18828 33544
rect 19334 33532 19340 33544
rect 19392 33532 19398 33584
rect 23474 33532 23480 33584
rect 23532 33572 23538 33584
rect 23584 33581 23612 33612
rect 24762 33600 24768 33612
rect 24820 33600 24826 33652
rect 27706 33640 27712 33652
rect 27667 33612 27712 33640
rect 27706 33600 27712 33612
rect 27764 33600 27770 33652
rect 30558 33640 30564 33652
rect 28092 33612 30564 33640
rect 23569 33575 23627 33581
rect 23569 33572 23581 33575
rect 23532 33544 23581 33572
rect 23532 33532 23538 33544
rect 23569 33541 23581 33544
rect 23615 33541 23627 33575
rect 23569 33535 23627 33541
rect 23937 33575 23995 33581
rect 23937 33541 23949 33575
rect 23983 33572 23995 33575
rect 24946 33572 24952 33584
rect 23983 33544 24624 33572
rect 23983 33541 23995 33544
rect 23937 33535 23995 33541
rect 18555 33476 18828 33504
rect 19153 33507 19211 33513
rect 18555 33473 18567 33476
rect 18509 33467 18567 33473
rect 19153 33473 19165 33507
rect 19199 33504 19211 33507
rect 19702 33504 19708 33516
rect 19199 33476 19708 33504
rect 19199 33473 19211 33476
rect 19153 33467 19211 33473
rect 19702 33464 19708 33476
rect 19760 33464 19766 33516
rect 23753 33507 23811 33513
rect 23753 33473 23765 33507
rect 23799 33473 23811 33507
rect 24394 33504 24400 33516
rect 24355 33476 24400 33504
rect 23753 33467 23811 33473
rect 15712 33408 16712 33436
rect 15712 33396 15718 33408
rect 17126 33396 17132 33448
rect 17184 33436 17190 33448
rect 18141 33439 18199 33445
rect 18141 33436 18153 33439
rect 17184 33408 18153 33436
rect 17184 33396 17190 33408
rect 18141 33405 18153 33408
rect 18187 33405 18199 33439
rect 23768 33436 23796 33467
rect 24394 33464 24400 33476
rect 24452 33464 24458 33516
rect 24596 33513 24624 33544
rect 24688 33544 24952 33572
rect 24688 33513 24716 33544
rect 24946 33532 24952 33544
rect 25004 33532 25010 33584
rect 24581 33507 24639 33513
rect 24581 33473 24593 33507
rect 24627 33473 24639 33507
rect 24581 33467 24639 33473
rect 24673 33507 24731 33513
rect 24673 33473 24685 33507
rect 24719 33473 24731 33507
rect 24673 33467 24731 33473
rect 24762 33464 24768 33516
rect 24820 33504 24826 33516
rect 24820 33476 25636 33504
rect 24820 33464 24826 33476
rect 25130 33436 25136 33448
rect 23768 33408 25136 33436
rect 18141 33399 18199 33405
rect 25130 33396 25136 33408
rect 25188 33396 25194 33448
rect 25608 33445 25636 33476
rect 27154 33464 27160 33516
rect 27212 33504 27218 33516
rect 28092 33513 28120 33612
rect 30558 33600 30564 33612
rect 30616 33600 30622 33652
rect 34146 33640 34152 33652
rect 31726 33612 34152 33640
rect 29181 33575 29239 33581
rect 29181 33541 29193 33575
rect 29227 33572 29239 33575
rect 30098 33572 30104 33584
rect 29227 33544 30104 33572
rect 29227 33541 29239 33544
rect 29181 33535 29239 33541
rect 30098 33532 30104 33544
rect 30156 33532 30162 33584
rect 30576 33519 30604 33600
rect 27985 33507 28043 33513
rect 27985 33504 27997 33507
rect 27212 33476 27997 33504
rect 27212 33464 27218 33476
rect 27985 33473 27997 33476
rect 28031 33473 28043 33507
rect 27985 33467 28043 33473
rect 28077 33507 28135 33513
rect 28077 33473 28089 33507
rect 28123 33473 28135 33507
rect 28077 33467 28135 33473
rect 28169 33507 28227 33513
rect 28169 33473 28181 33507
rect 28215 33473 28227 33507
rect 28350 33504 28356 33516
rect 28311 33476 28356 33504
rect 28169 33467 28227 33473
rect 25593 33439 25651 33445
rect 25593 33405 25605 33439
rect 25639 33436 25651 33439
rect 28184 33436 28212 33467
rect 28350 33464 28356 33476
rect 28408 33464 28414 33516
rect 28997 33507 29055 33513
rect 28997 33473 29009 33507
rect 29043 33504 29055 33507
rect 29086 33504 29092 33516
rect 29043 33476 29092 33504
rect 29043 33473 29055 33476
rect 28997 33467 29055 33473
rect 29086 33464 29092 33476
rect 29144 33464 29150 33516
rect 30190 33464 30196 33516
rect 30248 33504 30254 33516
rect 30466 33513 30472 33516
rect 30285 33507 30343 33513
rect 30285 33504 30297 33507
rect 30248 33476 30297 33504
rect 30248 33464 30254 33476
rect 30285 33473 30297 33476
rect 30331 33473 30343 33507
rect 30464 33504 30472 33513
rect 30427 33476 30472 33504
rect 30285 33467 30343 33473
rect 30464 33467 30472 33476
rect 30466 33464 30472 33467
rect 30524 33464 30530 33516
rect 30564 33513 30622 33519
rect 30564 33479 30576 33513
rect 30610 33479 30622 33513
rect 30564 33473 30622 33479
rect 30653 33507 30711 33513
rect 30653 33473 30665 33507
rect 30699 33473 30711 33507
rect 30653 33467 30711 33473
rect 28813 33439 28871 33445
rect 28813 33436 28825 33439
rect 25639 33408 26372 33436
rect 28184 33408 28825 33436
rect 25639 33405 25651 33408
rect 25593 33399 25651 33405
rect 3881 33371 3939 33377
rect 3881 33337 3893 33371
rect 3927 33337 3939 33371
rect 3881 33331 3939 33337
rect 25041 33371 25099 33377
rect 25041 33337 25053 33371
rect 25087 33368 25099 33371
rect 26234 33368 26240 33380
rect 25087 33340 26240 33368
rect 25087 33337 25099 33340
rect 25041 33331 25099 33337
rect 26234 33328 26240 33340
rect 26292 33328 26298 33380
rect 26344 33368 26372 33408
rect 28813 33405 28825 33408
rect 28859 33405 28871 33439
rect 28813 33399 28871 33405
rect 30374 33396 30380 33448
rect 30432 33436 30438 33448
rect 30668 33436 30696 33467
rect 30432 33408 30696 33436
rect 30432 33396 30438 33408
rect 31726 33368 31754 33612
rect 34146 33600 34152 33612
rect 34204 33600 34210 33652
rect 34517 33575 34575 33581
rect 34517 33541 34529 33575
rect 34563 33572 34575 33575
rect 36090 33575 36148 33581
rect 36090 33572 36102 33575
rect 34563 33544 36102 33572
rect 34563 33541 34575 33544
rect 34517 33535 34575 33541
rect 36090 33541 36102 33544
rect 36136 33541 36148 33575
rect 36090 33535 36148 33541
rect 33594 33464 33600 33516
rect 33652 33504 33658 33516
rect 33873 33507 33931 33513
rect 33873 33504 33885 33507
rect 33652 33476 33885 33504
rect 33652 33464 33658 33476
rect 33873 33473 33885 33476
rect 33919 33473 33931 33507
rect 34054 33504 34060 33516
rect 34015 33476 34060 33504
rect 33873 33467 33931 33473
rect 34054 33464 34060 33476
rect 34112 33464 34118 33516
rect 34149 33507 34207 33513
rect 34149 33473 34161 33507
rect 34195 33473 34207 33507
rect 34149 33467 34207 33473
rect 34241 33507 34299 33513
rect 34241 33473 34253 33507
rect 34287 33504 34299 33507
rect 34422 33504 34428 33516
rect 34287 33476 34428 33504
rect 34287 33473 34299 33476
rect 34241 33467 34299 33473
rect 31846 33396 31852 33448
rect 31904 33436 31910 33448
rect 32401 33439 32459 33445
rect 32401 33436 32413 33439
rect 31904 33408 32413 33436
rect 31904 33396 31910 33408
rect 32401 33405 32413 33408
rect 32447 33405 32459 33439
rect 32401 33399 32459 33405
rect 32677 33439 32735 33445
rect 32677 33405 32689 33439
rect 32723 33436 32735 33439
rect 34164 33436 34192 33467
rect 34422 33464 34428 33476
rect 34480 33464 34486 33516
rect 36262 33464 36268 33516
rect 36320 33504 36326 33516
rect 36357 33507 36415 33513
rect 36357 33504 36369 33507
rect 36320 33476 36369 33504
rect 36320 33464 36326 33476
rect 36357 33473 36369 33476
rect 36403 33473 36415 33507
rect 36357 33467 36415 33473
rect 34514 33436 34520 33448
rect 32723 33408 34520 33436
rect 32723 33405 32735 33408
rect 32677 33399 32735 33405
rect 34514 33396 34520 33408
rect 34572 33436 34578 33448
rect 34974 33436 34980 33448
rect 34572 33408 34980 33436
rect 34572 33396 34578 33408
rect 34974 33396 34980 33408
rect 35032 33396 35038 33448
rect 58158 33368 58164 33380
rect 26344 33340 31754 33368
rect 58119 33340 58164 33368
rect 58158 33328 58164 33340
rect 58216 33328 58222 33380
rect 17586 33260 17592 33312
rect 17644 33300 17650 33312
rect 18230 33300 18236 33312
rect 17644 33272 18236 33300
rect 17644 33260 17650 33272
rect 18230 33260 18236 33272
rect 18288 33260 18294 33312
rect 19702 33300 19708 33312
rect 19663 33272 19708 33300
rect 19702 33260 19708 33272
rect 19760 33260 19766 33312
rect 27154 33300 27160 33312
rect 27115 33272 27160 33300
rect 27154 33260 27160 33272
rect 27212 33260 27218 33312
rect 29362 33260 29368 33312
rect 29420 33300 29426 33312
rect 29733 33303 29791 33309
rect 29733 33300 29745 33303
rect 29420 33272 29745 33300
rect 29420 33260 29426 33272
rect 29733 33269 29745 33272
rect 29779 33300 29791 33303
rect 30374 33300 30380 33312
rect 29779 33272 30380 33300
rect 29779 33269 29791 33272
rect 29733 33263 29791 33269
rect 30374 33260 30380 33272
rect 30432 33260 30438 33312
rect 30834 33260 30840 33312
rect 30892 33300 30898 33312
rect 30929 33303 30987 33309
rect 30929 33300 30941 33303
rect 30892 33272 30941 33300
rect 30892 33260 30898 33272
rect 30929 33269 30941 33272
rect 30975 33269 30987 33303
rect 30929 33263 30987 33269
rect 34514 33260 34520 33312
rect 34572 33300 34578 33312
rect 34977 33303 35035 33309
rect 34977 33300 34989 33303
rect 34572 33272 34989 33300
rect 34572 33260 34578 33272
rect 34977 33269 34989 33272
rect 35023 33269 35035 33303
rect 34977 33263 35035 33269
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 6825 33099 6883 33105
rect 6825 33065 6837 33099
rect 6871 33096 6883 33099
rect 6914 33096 6920 33108
rect 6871 33068 6920 33096
rect 6871 33065 6883 33068
rect 6825 33059 6883 33065
rect 6914 33056 6920 33068
rect 6972 33056 6978 33108
rect 13814 33056 13820 33108
rect 13872 33096 13878 33108
rect 18046 33096 18052 33108
rect 13872 33068 18052 33096
rect 13872 33056 13878 33068
rect 18046 33056 18052 33068
rect 18104 33056 18110 33108
rect 23845 33099 23903 33105
rect 23845 33065 23857 33099
rect 23891 33096 23903 33099
rect 24578 33096 24584 33108
rect 23891 33068 24584 33096
rect 23891 33065 23903 33068
rect 23845 33059 23903 33065
rect 24578 33056 24584 33068
rect 24636 33056 24642 33108
rect 24854 33056 24860 33108
rect 24912 33096 24918 33108
rect 25130 33096 25136 33108
rect 24912 33068 25136 33096
rect 24912 33056 24918 33068
rect 25130 33056 25136 33068
rect 25188 33056 25194 33108
rect 29549 33099 29607 33105
rect 29549 33096 29561 33099
rect 25240 33068 29561 33096
rect 15838 32988 15844 33040
rect 15896 33028 15902 33040
rect 18417 33031 18475 33037
rect 18417 33028 18429 33031
rect 15896 33000 18429 33028
rect 15896 32988 15902 33000
rect 7926 32960 7932 32972
rect 7208 32932 7932 32960
rect 7208 32901 7236 32932
rect 7926 32920 7932 32932
rect 7984 32920 7990 32972
rect 16390 32920 16396 32972
rect 16448 32960 16454 32972
rect 16448 32932 16712 32960
rect 16448 32920 16454 32932
rect 7101 32895 7159 32901
rect 7101 32892 7113 32895
rect 6564 32864 7113 32892
rect 6564 32768 6592 32864
rect 7101 32861 7113 32864
rect 7147 32861 7159 32895
rect 7101 32855 7159 32861
rect 7193 32895 7251 32901
rect 7193 32861 7205 32895
rect 7239 32861 7251 32895
rect 7193 32855 7251 32861
rect 7285 32895 7343 32901
rect 7285 32861 7297 32895
rect 7331 32861 7343 32895
rect 7466 32892 7472 32904
rect 7427 32864 7472 32892
rect 7285 32855 7343 32861
rect 7300 32824 7328 32855
rect 7466 32852 7472 32864
rect 7524 32852 7530 32904
rect 8113 32895 8171 32901
rect 8113 32861 8125 32895
rect 8159 32892 8171 32895
rect 8202 32892 8208 32904
rect 8159 32864 8208 32892
rect 8159 32861 8171 32864
rect 8113 32855 8171 32861
rect 8202 32852 8208 32864
rect 8260 32852 8266 32904
rect 14090 32892 14096 32904
rect 14051 32864 14096 32892
rect 14090 32852 14096 32864
rect 14148 32852 14154 32904
rect 14918 32852 14924 32904
rect 14976 32892 14982 32904
rect 16209 32895 16267 32901
rect 16209 32892 16221 32895
rect 14976 32864 16221 32892
rect 14976 32852 14982 32864
rect 16209 32861 16221 32864
rect 16255 32861 16267 32895
rect 16209 32855 16267 32861
rect 16298 32852 16304 32904
rect 16356 32892 16362 32904
rect 16356 32864 16401 32892
rect 16356 32852 16362 32864
rect 16482 32852 16488 32904
rect 16540 32892 16546 32904
rect 16684 32901 16712 32932
rect 16674 32895 16732 32901
rect 16540 32864 16585 32892
rect 16540 32852 16546 32864
rect 16674 32861 16686 32895
rect 16720 32861 16732 32895
rect 17052 32892 17080 33000
rect 18417 32997 18429 33000
rect 18463 32997 18475 33031
rect 19797 33031 19855 33037
rect 19797 33028 19809 33031
rect 18417 32991 18475 32997
rect 18524 33000 19809 33028
rect 17126 32920 17132 32972
rect 17184 32960 17190 32972
rect 18524 32960 18552 33000
rect 19797 32997 19809 33000
rect 19843 33028 19855 33031
rect 23750 33028 23756 33040
rect 19843 33000 23756 33028
rect 19843 32997 19855 33000
rect 19797 32991 19855 32997
rect 23750 32988 23756 33000
rect 23808 32988 23814 33040
rect 24210 32988 24216 33040
rect 24268 33028 24274 33040
rect 25240 33028 25268 33068
rect 29549 33065 29561 33068
rect 29595 33065 29607 33099
rect 29549 33059 29607 33065
rect 31941 33099 31999 33105
rect 31941 33065 31953 33099
rect 31987 33096 31999 33099
rect 32214 33096 32220 33108
rect 31987 33068 32220 33096
rect 31987 33065 31999 33068
rect 31941 33059 31999 33065
rect 32214 33056 32220 33068
rect 32272 33056 32278 33108
rect 34054 33056 34060 33108
rect 34112 33096 34118 33108
rect 34149 33099 34207 33105
rect 34149 33096 34161 33099
rect 34112 33068 34161 33096
rect 34112 33056 34118 33068
rect 34149 33065 34161 33068
rect 34195 33065 34207 33099
rect 34149 33059 34207 33065
rect 34606 33056 34612 33108
rect 34664 33096 34670 33108
rect 34790 33096 34796 33108
rect 34664 33068 34796 33096
rect 34664 33056 34670 33068
rect 34790 33056 34796 33068
rect 34848 33096 34854 33108
rect 34885 33099 34943 33105
rect 34885 33096 34897 33099
rect 34848 33068 34897 33096
rect 34848 33056 34854 33068
rect 34885 33065 34897 33068
rect 34931 33065 34943 33099
rect 35894 33096 35900 33108
rect 34885 33059 34943 33065
rect 35360 33068 35900 33096
rect 24268 33000 25268 33028
rect 24268 32988 24274 33000
rect 30190 32988 30196 33040
rect 30248 33028 30254 33040
rect 35360 33028 35388 33068
rect 35894 33056 35900 33068
rect 35952 33056 35958 33108
rect 30248 33000 35388 33028
rect 30248 32988 30254 33000
rect 17184 32932 17448 32960
rect 17184 32920 17190 32932
rect 17313 32895 17371 32901
rect 17313 32892 17325 32895
rect 17052 32864 17325 32892
rect 16674 32855 16732 32861
rect 17313 32861 17325 32864
rect 17359 32861 17371 32895
rect 17420 32892 17448 32932
rect 18432 32932 18552 32960
rect 17586 32901 17592 32904
rect 17476 32895 17534 32901
rect 17476 32892 17488 32895
rect 17420 32864 17488 32892
rect 17313 32855 17371 32861
rect 17476 32861 17488 32864
rect 17522 32861 17534 32895
rect 17476 32855 17534 32861
rect 17576 32895 17592 32901
rect 17576 32861 17588 32895
rect 17576 32855 17592 32861
rect 17586 32852 17592 32855
rect 17644 32852 17650 32904
rect 17678 32852 17684 32904
rect 17736 32892 17742 32904
rect 18432 32892 18460 32932
rect 18598 32920 18604 32972
rect 18656 32920 18662 32972
rect 29178 32920 29184 32972
rect 29236 32960 29242 32972
rect 33321 32963 33379 32969
rect 29236 32932 30144 32960
rect 29236 32920 29242 32932
rect 18616 32892 18644 32920
rect 23474 32892 23480 32904
rect 17736 32864 18460 32892
rect 18524 32864 18644 32892
rect 23435 32864 23480 32892
rect 17736 32852 17742 32864
rect 7929 32827 7987 32833
rect 7929 32824 7941 32827
rect 7300 32796 7941 32824
rect 7929 32793 7941 32796
rect 7975 32793 7987 32827
rect 7929 32787 7987 32793
rect 8297 32827 8355 32833
rect 8297 32793 8309 32827
rect 8343 32793 8355 32827
rect 8297 32787 8355 32793
rect 14360 32827 14418 32833
rect 14360 32793 14372 32827
rect 14406 32824 14418 32827
rect 14458 32824 14464 32836
rect 14406 32796 14464 32824
rect 14406 32793 14418 32796
rect 14360 32787 14418 32793
rect 3881 32759 3939 32765
rect 3881 32725 3893 32759
rect 3927 32756 3939 32759
rect 4062 32756 4068 32768
rect 3927 32728 4068 32756
rect 3927 32725 3939 32728
rect 3881 32719 3939 32725
rect 4062 32716 4068 32728
rect 4120 32716 4126 32768
rect 6365 32759 6423 32765
rect 6365 32725 6377 32759
rect 6411 32756 6423 32759
rect 6546 32756 6552 32768
rect 6411 32728 6552 32756
rect 6411 32725 6423 32728
rect 6365 32719 6423 32725
rect 6546 32716 6552 32728
rect 6604 32716 6610 32768
rect 7374 32716 7380 32768
rect 7432 32756 7438 32768
rect 8202 32756 8208 32768
rect 7432 32728 8208 32756
rect 7432 32716 7438 32728
rect 8202 32716 8208 32728
rect 8260 32756 8266 32768
rect 8312 32756 8340 32787
rect 14458 32784 14464 32796
rect 14516 32784 14522 32836
rect 16577 32827 16635 32833
rect 16577 32793 16589 32827
rect 16623 32824 16635 32827
rect 18524 32824 18552 32864
rect 23474 32852 23480 32864
rect 23532 32852 23538 32904
rect 26234 32852 26240 32904
rect 26292 32901 26298 32904
rect 26292 32892 26304 32901
rect 26510 32892 26516 32904
rect 26292 32864 26337 32892
rect 26423 32864 26516 32892
rect 26292 32855 26304 32864
rect 26292 32852 26298 32855
rect 26510 32852 26516 32864
rect 26568 32892 26574 32904
rect 29730 32892 29736 32904
rect 26568 32864 27476 32892
rect 29691 32864 29736 32892
rect 26568 32852 26574 32864
rect 16623 32796 18552 32824
rect 18601 32827 18659 32833
rect 16623 32793 16635 32796
rect 16577 32787 16635 32793
rect 18601 32793 18613 32827
rect 18647 32824 18659 32827
rect 19337 32827 19395 32833
rect 19337 32824 19349 32827
rect 18647 32796 19349 32824
rect 18647 32793 18659 32796
rect 18601 32787 18659 32793
rect 19337 32793 19349 32796
rect 19383 32824 19395 32827
rect 19702 32824 19708 32836
rect 19383 32796 19708 32824
rect 19383 32793 19395 32796
rect 19337 32787 19395 32793
rect 19702 32784 19708 32796
rect 19760 32824 19766 32836
rect 23658 32824 23664 32836
rect 19760 32796 22094 32824
rect 23619 32796 23664 32824
rect 19760 32784 19766 32796
rect 8260 32728 8340 32756
rect 8260 32716 8266 32728
rect 15194 32716 15200 32768
rect 15252 32756 15258 32768
rect 15473 32759 15531 32765
rect 15473 32756 15485 32759
rect 15252 32728 15485 32756
rect 15252 32716 15258 32728
rect 15473 32725 15485 32728
rect 15519 32725 15531 32759
rect 15473 32719 15531 32725
rect 16853 32759 16911 32765
rect 16853 32725 16865 32759
rect 16899 32756 16911 32759
rect 17862 32756 17868 32768
rect 16899 32728 17868 32756
rect 16899 32725 16911 32728
rect 16853 32719 16911 32725
rect 17862 32716 17868 32728
rect 17920 32716 17926 32768
rect 17957 32759 18015 32765
rect 17957 32725 17969 32759
rect 18003 32756 18015 32759
rect 18414 32756 18420 32768
rect 18003 32728 18420 32756
rect 18003 32725 18015 32728
rect 17957 32719 18015 32725
rect 18414 32716 18420 32728
rect 18472 32716 18478 32768
rect 22066 32756 22094 32796
rect 23658 32784 23664 32796
rect 23716 32784 23722 32836
rect 23566 32756 23572 32768
rect 22066 32728 23572 32756
rect 23566 32716 23572 32728
rect 23624 32716 23630 32768
rect 27448 32765 27476 32864
rect 29730 32852 29736 32864
rect 29788 32852 29794 32904
rect 30116 32901 30144 32932
rect 33321 32929 33333 32963
rect 33367 32960 33379 32963
rect 34422 32960 34428 32972
rect 33367 32932 34428 32960
rect 33367 32929 33379 32932
rect 33321 32923 33379 32929
rect 34422 32920 34428 32932
rect 34480 32920 34486 32972
rect 29825 32895 29883 32901
rect 29825 32861 29837 32895
rect 29871 32861 29883 32895
rect 29825 32855 29883 32861
rect 30101 32895 30159 32901
rect 30101 32861 30113 32895
rect 30147 32861 30159 32895
rect 31018 32892 31024 32904
rect 30101 32855 30159 32861
rect 30668 32864 31024 32892
rect 28721 32827 28779 32833
rect 28721 32793 28733 32827
rect 28767 32824 28779 32827
rect 28994 32824 29000 32836
rect 28767 32796 29000 32824
rect 28767 32793 28779 32796
rect 28721 32787 28779 32793
rect 28994 32784 29000 32796
rect 29052 32784 29058 32836
rect 29270 32784 29276 32836
rect 29328 32824 29334 32836
rect 29840 32824 29868 32855
rect 29328 32796 29868 32824
rect 29917 32827 29975 32833
rect 29328 32784 29334 32796
rect 29917 32793 29929 32827
rect 29963 32824 29975 32827
rect 30190 32824 30196 32836
rect 29963 32796 30196 32824
rect 29963 32793 29975 32796
rect 29917 32787 29975 32793
rect 30190 32784 30196 32796
rect 30248 32784 30254 32836
rect 30668 32768 30696 32864
rect 31018 32852 31024 32864
rect 31076 32852 31082 32904
rect 31478 32852 31484 32904
rect 31536 32892 31542 32904
rect 32217 32895 32275 32901
rect 32217 32892 32229 32895
rect 31536 32864 32229 32892
rect 31536 32852 31542 32864
rect 32217 32861 32229 32864
rect 32263 32861 32275 32895
rect 32217 32855 32275 32861
rect 32309 32895 32367 32901
rect 32309 32861 32321 32895
rect 32355 32861 32367 32895
rect 32309 32855 32367 32861
rect 32401 32895 32459 32901
rect 32401 32861 32413 32895
rect 32447 32892 32459 32895
rect 32490 32892 32496 32904
rect 32447 32864 32496 32892
rect 32447 32861 32459 32864
rect 32401 32855 32459 32861
rect 30745 32827 30803 32833
rect 30745 32793 30757 32827
rect 30791 32824 30803 32827
rect 31294 32824 31300 32836
rect 30791 32796 31300 32824
rect 30791 32793 30803 32796
rect 30745 32787 30803 32793
rect 31294 32784 31300 32796
rect 31352 32824 31358 32836
rect 31846 32824 31852 32836
rect 31352 32796 31852 32824
rect 31352 32784 31358 32796
rect 31846 32784 31852 32796
rect 31904 32824 31910 32836
rect 32324 32824 32352 32855
rect 32490 32852 32496 32864
rect 32548 32852 32554 32904
rect 32585 32895 32643 32901
rect 32585 32861 32597 32895
rect 32631 32892 32643 32895
rect 33594 32892 33600 32904
rect 32631 32864 33600 32892
rect 32631 32861 32643 32864
rect 32585 32855 32643 32861
rect 33594 32852 33600 32864
rect 33652 32852 33658 32904
rect 33778 32892 33784 32904
rect 33739 32864 33784 32892
rect 33778 32852 33784 32864
rect 33836 32852 33842 32904
rect 33965 32895 34023 32901
rect 33965 32861 33977 32895
rect 34011 32892 34023 32895
rect 34514 32892 34520 32904
rect 34011 32864 34520 32892
rect 34011 32861 34023 32864
rect 33965 32855 34023 32861
rect 34514 32852 34520 32864
rect 34572 32852 34578 32904
rect 35986 32852 35992 32904
rect 36044 32901 36050 32904
rect 36044 32892 36056 32901
rect 36262 32892 36268 32904
rect 36044 32864 36089 32892
rect 36223 32864 36268 32892
rect 36044 32855 36056 32864
rect 36044 32852 36050 32855
rect 36262 32852 36268 32864
rect 36320 32852 36326 32904
rect 31904 32796 32352 32824
rect 31904 32784 31910 32796
rect 27433 32759 27491 32765
rect 27433 32725 27445 32759
rect 27479 32756 27491 32759
rect 27522 32756 27528 32768
rect 27479 32728 27528 32756
rect 27479 32725 27491 32728
rect 27433 32719 27491 32725
rect 27522 32716 27528 32728
rect 27580 32716 27586 32768
rect 30650 32756 30656 32768
rect 30611 32728 30656 32756
rect 30650 32716 30656 32728
rect 30708 32716 30714 32768
rect 30926 32716 30932 32768
rect 30984 32756 30990 32768
rect 31389 32759 31447 32765
rect 31389 32756 31401 32759
rect 30984 32728 31401 32756
rect 30984 32716 30990 32728
rect 31389 32725 31401 32728
rect 31435 32756 31447 32759
rect 31478 32756 31484 32768
rect 31435 32728 31484 32756
rect 31435 32725 31447 32728
rect 31389 32719 31447 32725
rect 31478 32716 31484 32728
rect 31536 32716 31542 32768
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 7466 32512 7472 32564
rect 7524 32552 7530 32564
rect 8297 32555 8355 32561
rect 8297 32552 8309 32555
rect 7524 32524 8309 32552
rect 7524 32512 7530 32524
rect 8297 32521 8309 32524
rect 8343 32552 8355 32555
rect 9766 32552 9772 32564
rect 8343 32524 9772 32552
rect 8343 32521 8355 32524
rect 8297 32515 8355 32521
rect 9766 32512 9772 32524
rect 9824 32512 9830 32564
rect 10870 32512 10876 32564
rect 10928 32552 10934 32564
rect 14182 32552 14188 32564
rect 10928 32524 14188 32552
rect 10928 32512 10934 32524
rect 14182 32512 14188 32524
rect 14240 32512 14246 32564
rect 14458 32552 14464 32564
rect 14419 32524 14464 32552
rect 14458 32512 14464 32524
rect 14516 32512 14522 32564
rect 17310 32512 17316 32564
rect 17368 32552 17374 32564
rect 18417 32555 18475 32561
rect 18417 32552 18429 32555
rect 17368 32524 18429 32552
rect 17368 32512 17374 32524
rect 18417 32521 18429 32524
rect 18463 32521 18475 32555
rect 18417 32515 18475 32521
rect 8938 32444 8944 32496
rect 8996 32484 9002 32496
rect 10229 32487 10287 32493
rect 10229 32484 10241 32487
rect 8996 32456 10241 32484
rect 8996 32444 9002 32456
rect 10229 32453 10241 32456
rect 10275 32453 10287 32487
rect 10229 32447 10287 32453
rect 12529 32487 12587 32493
rect 12529 32453 12541 32487
rect 12575 32484 12587 32487
rect 12618 32484 12624 32496
rect 12575 32456 12624 32484
rect 12575 32453 12587 32456
rect 12529 32447 12587 32453
rect 12618 32444 12624 32456
rect 12676 32484 12682 32496
rect 13078 32484 13084 32496
rect 12676 32456 13084 32484
rect 12676 32444 12682 32456
rect 13078 32444 13084 32456
rect 13136 32444 13142 32496
rect 13446 32444 13452 32496
rect 13504 32484 13510 32496
rect 14366 32484 14372 32496
rect 13504 32456 14372 32484
rect 13504 32444 13510 32456
rect 2222 32416 2228 32428
rect 2183 32388 2228 32416
rect 2222 32376 2228 32388
rect 2280 32376 2286 32428
rect 2314 32376 2320 32428
rect 2372 32416 2378 32428
rect 2481 32419 2539 32425
rect 2481 32416 2493 32419
rect 2372 32388 2493 32416
rect 2372 32376 2378 32388
rect 2481 32385 2493 32388
rect 2527 32385 2539 32419
rect 6362 32416 6368 32428
rect 6323 32388 6368 32416
rect 2481 32379 2539 32385
rect 6362 32376 6368 32388
rect 6420 32376 6426 32428
rect 6454 32376 6460 32428
rect 6512 32416 6518 32428
rect 6621 32419 6679 32425
rect 6621 32416 6633 32419
rect 6512 32388 6633 32416
rect 6512 32376 6518 32388
rect 6621 32385 6633 32388
rect 6667 32385 6679 32419
rect 6621 32379 6679 32385
rect 8202 32376 8208 32428
rect 8260 32416 8266 32428
rect 9493 32419 9551 32425
rect 9493 32416 9505 32419
rect 8260 32388 9505 32416
rect 8260 32376 8266 32388
rect 9493 32385 9505 32388
rect 9539 32385 9551 32419
rect 9493 32379 9551 32385
rect 10413 32419 10471 32425
rect 10413 32385 10425 32419
rect 10459 32416 10471 32419
rect 11054 32416 11060 32428
rect 10459 32388 11060 32416
rect 10459 32385 10471 32388
rect 10413 32379 10471 32385
rect 11054 32376 11060 32388
rect 11112 32376 11118 32428
rect 12713 32419 12771 32425
rect 12713 32385 12725 32419
rect 12759 32416 12771 32419
rect 12894 32416 12900 32428
rect 12759 32388 12900 32416
rect 12759 32385 12771 32388
rect 12713 32379 12771 32385
rect 12894 32376 12900 32388
rect 12952 32376 12958 32428
rect 13814 32416 13820 32428
rect 13775 32388 13820 32416
rect 13814 32376 13820 32388
rect 13872 32376 13878 32428
rect 14108 32425 14136 32456
rect 14366 32444 14372 32456
rect 14424 32444 14430 32496
rect 15105 32487 15163 32493
rect 15105 32453 15117 32487
rect 15151 32484 15163 32487
rect 15194 32484 15200 32496
rect 15151 32456 15200 32484
rect 15151 32453 15163 32456
rect 15105 32447 15163 32453
rect 15194 32444 15200 32456
rect 15252 32484 15258 32496
rect 15378 32484 15384 32496
rect 15252 32456 15384 32484
rect 15252 32444 15258 32456
rect 15378 32444 15384 32456
rect 15436 32444 15442 32496
rect 16117 32487 16175 32493
rect 16117 32453 16129 32487
rect 16163 32484 16175 32487
rect 17586 32484 17592 32496
rect 16163 32456 17592 32484
rect 16163 32453 16175 32456
rect 16117 32447 16175 32453
rect 17586 32444 17592 32456
rect 17644 32444 17650 32496
rect 14001 32419 14059 32425
rect 14001 32385 14013 32419
rect 14047 32385 14059 32419
rect 14001 32379 14059 32385
rect 14093 32419 14151 32425
rect 14093 32385 14105 32419
rect 14139 32385 14151 32419
rect 14093 32379 14151 32385
rect 9769 32351 9827 32357
rect 9769 32317 9781 32351
rect 9815 32348 9827 32351
rect 12066 32348 12072 32360
rect 9815 32320 12072 32348
rect 9815 32317 9827 32320
rect 9769 32311 9827 32317
rect 12066 32308 12072 32320
rect 12124 32308 12130 32360
rect 14016 32348 14044 32379
rect 14182 32376 14188 32428
rect 14240 32416 14246 32428
rect 14240 32388 14285 32416
rect 14240 32376 14246 32388
rect 14550 32376 14556 32428
rect 14608 32416 14614 32428
rect 14918 32416 14924 32428
rect 14608 32388 14924 32416
rect 14608 32376 14614 32388
rect 14918 32376 14924 32388
rect 14976 32376 14982 32428
rect 15562 32376 15568 32428
rect 15620 32416 15626 32428
rect 15933 32419 15991 32425
rect 15933 32416 15945 32419
rect 15620 32388 15945 32416
rect 15620 32376 15626 32388
rect 15933 32385 15945 32388
rect 15979 32385 15991 32419
rect 17126 32416 17132 32428
rect 17087 32388 17132 32416
rect 15933 32379 15991 32385
rect 17126 32376 17132 32388
rect 17184 32376 17190 32428
rect 18432 32416 18460 32515
rect 18598 32512 18604 32564
rect 18656 32552 18662 32564
rect 20717 32555 20775 32561
rect 20717 32552 20729 32555
rect 18656 32524 20729 32552
rect 18656 32512 18662 32524
rect 20717 32521 20729 32524
rect 20763 32521 20775 32555
rect 20717 32515 20775 32521
rect 23658 32512 23664 32564
rect 23716 32552 23722 32564
rect 24118 32552 24124 32564
rect 23716 32524 24124 32552
rect 23716 32512 23722 32524
rect 24118 32512 24124 32524
rect 24176 32512 24182 32564
rect 29730 32552 29736 32564
rect 28552 32524 29736 32552
rect 18506 32444 18512 32496
rect 18564 32484 18570 32496
rect 19582 32487 19640 32493
rect 19582 32484 19594 32487
rect 18564 32456 19594 32484
rect 18564 32444 18570 32456
rect 19582 32453 19594 32456
rect 19628 32453 19640 32487
rect 19582 32447 19640 32453
rect 25038 32444 25044 32496
rect 25096 32484 25102 32496
rect 25234 32487 25292 32493
rect 25234 32484 25246 32487
rect 25096 32456 25246 32484
rect 25096 32444 25102 32456
rect 25234 32453 25246 32456
rect 25280 32453 25292 32487
rect 25234 32447 25292 32453
rect 19242 32416 19248 32428
rect 18432 32388 19248 32416
rect 19242 32376 19248 32388
rect 19300 32416 19306 32428
rect 19337 32419 19395 32425
rect 19337 32416 19349 32419
rect 19300 32388 19349 32416
rect 19300 32376 19306 32388
rect 19337 32385 19349 32388
rect 19383 32385 19395 32419
rect 19337 32379 19395 32385
rect 19426 32376 19432 32428
rect 19484 32376 19490 32428
rect 22649 32419 22707 32425
rect 22649 32416 22661 32419
rect 22066 32388 22661 32416
rect 15289 32351 15347 32357
rect 15289 32348 15301 32351
rect 14016 32320 15301 32348
rect 15289 32317 15301 32320
rect 15335 32317 15347 32351
rect 15289 32311 15347 32317
rect 16942 32308 16948 32360
rect 17000 32348 17006 32360
rect 17310 32348 17316 32360
rect 17000 32320 17316 32348
rect 17000 32308 17006 32320
rect 17310 32308 17316 32320
rect 17368 32308 17374 32360
rect 17586 32308 17592 32360
rect 17644 32348 17650 32360
rect 19444 32348 19472 32376
rect 17644 32320 19472 32348
rect 17644 32308 17650 32320
rect 21174 32308 21180 32360
rect 21232 32348 21238 32360
rect 21269 32351 21327 32357
rect 21269 32348 21281 32351
rect 21232 32320 21281 32348
rect 21232 32308 21238 32320
rect 21269 32317 21281 32320
rect 21315 32348 21327 32351
rect 22066 32348 22094 32388
rect 22649 32385 22661 32388
rect 22695 32385 22707 32419
rect 22649 32379 22707 32385
rect 23477 32419 23535 32425
rect 23477 32385 23489 32419
rect 23523 32416 23535 32419
rect 24026 32416 24032 32428
rect 23523 32388 24032 32416
rect 23523 32385 23535 32388
rect 23477 32379 23535 32385
rect 24026 32376 24032 32388
rect 24084 32376 24090 32428
rect 25501 32419 25559 32425
rect 25501 32385 25513 32419
rect 25547 32416 25559 32419
rect 26510 32416 26516 32428
rect 25547 32388 26516 32416
rect 25547 32385 25559 32388
rect 25501 32379 25559 32385
rect 26510 32376 26516 32388
rect 26568 32376 26574 32428
rect 28552 32425 28580 32524
rect 29730 32512 29736 32524
rect 29788 32512 29794 32564
rect 29914 32552 29920 32564
rect 29875 32524 29920 32552
rect 29914 32512 29920 32524
rect 29972 32512 29978 32564
rect 32306 32512 32312 32564
rect 32364 32552 32370 32564
rect 36262 32552 36268 32564
rect 32364 32524 36268 32552
rect 32364 32512 32370 32524
rect 36262 32512 36268 32524
rect 36320 32512 36326 32564
rect 28629 32487 28687 32493
rect 28629 32453 28641 32487
rect 28675 32484 28687 32487
rect 29086 32484 29092 32496
rect 28675 32456 29092 32484
rect 28675 32453 28687 32456
rect 28629 32447 28687 32453
rect 29086 32444 29092 32456
rect 29144 32444 29150 32496
rect 32490 32484 32496 32496
rect 32451 32456 32496 32484
rect 32490 32444 32496 32456
rect 32548 32444 32554 32496
rect 28537 32419 28595 32425
rect 28537 32385 28549 32419
rect 28583 32385 28595 32419
rect 28537 32379 28595 32385
rect 28721 32419 28779 32425
rect 28721 32385 28733 32419
rect 28767 32385 28779 32419
rect 28721 32379 28779 32385
rect 21315 32320 22094 32348
rect 21315 32317 21327 32320
rect 21269 32311 21327 32317
rect 22186 32308 22192 32360
rect 22244 32348 22250 32360
rect 22373 32351 22431 32357
rect 22373 32348 22385 32351
rect 22244 32320 22385 32348
rect 22244 32308 22250 32320
rect 22373 32317 22385 32320
rect 22419 32317 22431 32351
rect 28736 32348 28764 32379
rect 28810 32376 28816 32428
rect 28868 32416 28874 32428
rect 28905 32419 28963 32425
rect 28905 32416 28917 32419
rect 28868 32388 28917 32416
rect 28868 32376 28874 32388
rect 28905 32385 28917 32388
rect 28951 32385 28963 32419
rect 28905 32379 28963 32385
rect 29638 32376 29644 32428
rect 29696 32416 29702 32428
rect 29733 32419 29791 32425
rect 29733 32416 29745 32419
rect 29696 32388 29745 32416
rect 29696 32376 29702 32388
rect 29733 32385 29745 32388
rect 29779 32416 29791 32419
rect 30469 32419 30527 32425
rect 30469 32416 30481 32419
rect 29779 32388 30481 32416
rect 29779 32385 29791 32388
rect 29733 32379 29791 32385
rect 30469 32385 30481 32388
rect 30515 32385 30527 32419
rect 30469 32379 30527 32385
rect 31754 32376 31760 32428
rect 31812 32416 31818 32428
rect 32125 32419 32183 32425
rect 32125 32416 32137 32419
rect 31812 32388 32137 32416
rect 31812 32376 31818 32388
rect 32125 32385 32137 32388
rect 32171 32416 32183 32419
rect 32214 32416 32220 32428
rect 32171 32388 32220 32416
rect 32171 32385 32183 32388
rect 32125 32379 32183 32385
rect 32214 32376 32220 32388
rect 32272 32376 32278 32428
rect 32309 32419 32367 32425
rect 32309 32385 32321 32419
rect 32355 32416 32367 32419
rect 33318 32416 33324 32428
rect 32355 32388 33324 32416
rect 32355 32385 32367 32388
rect 32309 32379 32367 32385
rect 33318 32376 33324 32388
rect 33376 32376 33382 32428
rect 34977 32419 35035 32425
rect 34977 32416 34989 32419
rect 34532 32388 34989 32416
rect 30190 32348 30196 32360
rect 28736 32320 30196 32348
rect 22373 32311 22431 32317
rect 30190 32308 30196 32320
rect 30248 32308 30254 32360
rect 17034 32280 17040 32292
rect 7300 32252 17040 32280
rect 3602 32212 3608 32224
rect 3563 32184 3608 32212
rect 3602 32172 3608 32184
rect 3660 32172 3666 32224
rect 6730 32172 6736 32224
rect 6788 32212 6794 32224
rect 7300 32212 7328 32252
rect 17034 32240 17040 32252
rect 17092 32240 17098 32292
rect 23474 32240 23480 32292
rect 23532 32280 23538 32292
rect 23661 32283 23719 32289
rect 23661 32280 23673 32283
rect 23532 32252 23673 32280
rect 23532 32240 23538 32252
rect 23661 32249 23673 32252
rect 23707 32249 23719 32283
rect 23661 32243 23719 32249
rect 27430 32240 27436 32292
rect 27488 32280 27494 32292
rect 27488 32252 28948 32280
rect 27488 32240 27494 32252
rect 6788 32184 7328 32212
rect 7745 32215 7803 32221
rect 6788 32172 6794 32184
rect 7745 32181 7757 32215
rect 7791 32212 7803 32215
rect 8110 32212 8116 32224
rect 7791 32184 8116 32212
rect 7791 32181 7803 32184
rect 7745 32175 7803 32181
rect 8110 32172 8116 32184
rect 8168 32172 8174 32224
rect 10134 32172 10140 32224
rect 10192 32212 10198 32224
rect 10597 32215 10655 32221
rect 10597 32212 10609 32215
rect 10192 32184 10609 32212
rect 10192 32172 10198 32184
rect 10597 32181 10609 32184
rect 10643 32181 10655 32215
rect 10597 32175 10655 32181
rect 12897 32215 12955 32221
rect 12897 32181 12909 32215
rect 12943 32212 12955 32215
rect 13354 32212 13360 32224
rect 12943 32184 13360 32212
rect 12943 32181 12955 32184
rect 12897 32175 12955 32181
rect 13354 32172 13360 32184
rect 13412 32172 13418 32224
rect 27706 32172 27712 32224
rect 27764 32212 27770 32224
rect 28353 32215 28411 32221
rect 28353 32212 28365 32215
rect 27764 32184 28365 32212
rect 27764 32172 27770 32184
rect 28353 32181 28365 32184
rect 28399 32181 28411 32215
rect 28920 32212 28948 32252
rect 28994 32240 29000 32292
rect 29052 32280 29058 32292
rect 30282 32280 30288 32292
rect 29052 32252 30288 32280
rect 29052 32240 29058 32252
rect 30282 32240 30288 32252
rect 30340 32280 30346 32292
rect 34532 32289 34560 32388
rect 34977 32385 34989 32388
rect 35023 32385 35035 32419
rect 34977 32379 35035 32385
rect 34517 32283 34575 32289
rect 34517 32280 34529 32283
rect 30340 32252 34529 32280
rect 30340 32240 30346 32252
rect 34517 32249 34529 32252
rect 34563 32249 34575 32283
rect 34517 32243 34575 32249
rect 31202 32212 31208 32224
rect 28920 32184 31208 32212
rect 28353 32175 28411 32181
rect 31202 32172 31208 32184
rect 31260 32172 31266 32224
rect 58158 32212 58164 32224
rect 58119 32184 58164 32212
rect 58158 32172 58164 32184
rect 58216 32172 58222 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 2041 32011 2099 32017
rect 2041 31977 2053 32011
rect 2087 32008 2099 32011
rect 2314 32008 2320 32020
rect 2087 31980 2320 32008
rect 2087 31977 2099 31980
rect 2041 31971 2099 31977
rect 2314 31968 2320 31980
rect 2372 31968 2378 32020
rect 6362 31968 6368 32020
rect 6420 32008 6426 32020
rect 7009 32011 7067 32017
rect 7009 32008 7021 32011
rect 6420 31980 7021 32008
rect 6420 31968 6426 31980
rect 7009 31977 7021 31980
rect 7055 31977 7067 32011
rect 7009 31971 7067 31977
rect 3234 31940 3240 31952
rect 2424 31912 3240 31940
rect 2424 31813 2452 31912
rect 3234 31900 3240 31912
rect 3292 31900 3298 31952
rect 7024 31872 7052 31971
rect 7282 31968 7288 32020
rect 7340 32008 7346 32020
rect 11790 32008 11796 32020
rect 7340 31980 11796 32008
rect 7340 31968 7346 31980
rect 11790 31968 11796 31980
rect 11848 31968 11854 32020
rect 12066 31968 12072 32020
rect 12124 32008 12130 32020
rect 14918 32008 14924 32020
rect 12124 31980 14924 32008
rect 12124 31968 12130 31980
rect 14918 31968 14924 31980
rect 14976 31968 14982 32020
rect 17037 32011 17095 32017
rect 17037 31977 17049 32011
rect 17083 32008 17095 32011
rect 17126 32008 17132 32020
rect 17083 31980 17132 32008
rect 17083 31977 17095 31980
rect 17037 31971 17095 31977
rect 17126 31968 17132 31980
rect 17184 31968 17190 32020
rect 20622 31968 20628 32020
rect 20680 32008 20686 32020
rect 27154 32008 27160 32020
rect 20680 31980 27160 32008
rect 20680 31968 20686 31980
rect 27154 31968 27160 31980
rect 27212 31968 27218 32020
rect 28905 32011 28963 32017
rect 28905 31977 28917 32011
rect 28951 32008 28963 32011
rect 28994 32008 29000 32020
rect 28951 31980 29000 32008
rect 28951 31977 28963 31980
rect 28905 31971 28963 31977
rect 28994 31968 29000 31980
rect 29052 31968 29058 32020
rect 29733 32011 29791 32017
rect 29733 31977 29745 32011
rect 29779 32008 29791 32011
rect 30006 32008 30012 32020
rect 29779 31980 30012 32008
rect 29779 31977 29791 31980
rect 29733 31971 29791 31977
rect 30006 31968 30012 31980
rect 30064 31968 30070 32020
rect 30742 32008 30748 32020
rect 30208 31980 30748 32008
rect 10689 31943 10747 31949
rect 10689 31909 10701 31943
rect 10735 31940 10747 31943
rect 11054 31940 11060 31952
rect 10735 31912 11060 31940
rect 10735 31909 10747 31912
rect 10689 31903 10747 31909
rect 11054 31900 11060 31912
rect 11112 31900 11118 31952
rect 14182 31940 14188 31952
rect 14143 31912 14188 31940
rect 14182 31900 14188 31912
rect 14240 31900 14246 31952
rect 17310 31900 17316 31952
rect 17368 31940 17374 31952
rect 21545 31943 21603 31949
rect 21545 31940 21557 31943
rect 17368 31912 21557 31940
rect 17368 31900 17374 31912
rect 21545 31909 21557 31912
rect 21591 31940 21603 31943
rect 22278 31940 22284 31952
rect 21591 31912 22284 31940
rect 21591 31909 21603 31912
rect 21545 31903 21603 31909
rect 22278 31900 22284 31912
rect 22336 31900 22342 31952
rect 28534 31900 28540 31952
rect 28592 31940 28598 31952
rect 30208 31940 30236 31980
rect 30742 31968 30748 31980
rect 30800 31968 30806 32020
rect 31202 31968 31208 32020
rect 31260 32008 31266 32020
rect 35529 32011 35587 32017
rect 35529 32008 35541 32011
rect 31260 31980 35541 32008
rect 31260 31968 31266 31980
rect 35529 31977 35541 31980
rect 35575 32008 35587 32011
rect 36446 32008 36452 32020
rect 35575 31980 36452 32008
rect 35575 31977 35587 31980
rect 35529 31971 35587 31977
rect 36446 31968 36452 31980
rect 36504 31968 36510 32020
rect 28592 31912 30236 31940
rect 28592 31900 28598 31912
rect 36262 31900 36268 31952
rect 36320 31940 36326 31952
rect 36320 31912 37596 31940
rect 36320 31900 36326 31912
rect 37568 31884 37596 31912
rect 9309 31875 9367 31881
rect 9309 31872 9321 31875
rect 7024 31844 9321 31872
rect 9309 31841 9321 31844
rect 9355 31841 9367 31875
rect 11422 31872 11428 31884
rect 11383 31844 11428 31872
rect 9309 31835 9367 31841
rect 11422 31832 11428 31844
rect 11480 31832 11486 31884
rect 17773 31875 17831 31881
rect 17773 31841 17785 31875
rect 17819 31872 17831 31875
rect 17954 31872 17960 31884
rect 17819 31844 17960 31872
rect 17819 31841 17831 31844
rect 17773 31835 17831 31841
rect 17954 31832 17960 31844
rect 18012 31832 18018 31884
rect 23569 31875 23627 31881
rect 23569 31841 23581 31875
rect 23615 31872 23627 31875
rect 24394 31872 24400 31884
rect 23615 31844 24400 31872
rect 23615 31841 23627 31844
rect 23569 31835 23627 31841
rect 24394 31832 24400 31844
rect 24452 31872 24458 31884
rect 24670 31872 24676 31884
rect 24452 31844 24676 31872
rect 24452 31832 24458 31844
rect 24670 31832 24676 31844
rect 24728 31832 24734 31884
rect 24946 31872 24952 31884
rect 24907 31844 24952 31872
rect 24946 31832 24952 31844
rect 25004 31832 25010 31884
rect 36725 31875 36783 31881
rect 36725 31841 36737 31875
rect 36771 31841 36783 31875
rect 37550 31872 37556 31884
rect 37463 31844 37556 31872
rect 36725 31835 36783 31841
rect 2271 31807 2329 31813
rect 2271 31773 2283 31807
rect 2317 31804 2329 31807
rect 2390 31807 2452 31813
rect 2317 31773 2340 31804
rect 2271 31767 2340 31773
rect 2390 31773 2402 31807
rect 2436 31776 2452 31807
rect 2522 31807 2580 31813
rect 2436 31773 2448 31776
rect 2390 31767 2448 31773
rect 2522 31773 2534 31807
rect 2568 31804 2580 31807
rect 2568 31776 2636 31804
rect 2568 31773 2580 31776
rect 2522 31767 2580 31773
rect 2312 31668 2340 31767
rect 2608 31736 2636 31776
rect 2682 31764 2688 31816
rect 2740 31804 2746 31816
rect 4982 31804 4988 31816
rect 2740 31776 4988 31804
rect 2740 31764 2746 31776
rect 4982 31764 4988 31776
rect 5040 31764 5046 31816
rect 5721 31807 5779 31813
rect 5721 31773 5733 31807
rect 5767 31804 5779 31807
rect 7282 31804 7288 31816
rect 5767 31776 7288 31804
rect 5767 31773 5779 31776
rect 5721 31767 5779 31773
rect 7282 31764 7288 31776
rect 7340 31764 7346 31816
rect 7558 31764 7564 31816
rect 7616 31804 7622 31816
rect 8297 31807 8355 31813
rect 8297 31804 8309 31807
rect 7616 31776 8309 31804
rect 7616 31764 7622 31776
rect 8297 31773 8309 31776
rect 8343 31773 8355 31807
rect 8297 31767 8355 31773
rect 9576 31807 9634 31813
rect 9576 31773 9588 31807
rect 9622 31804 9634 31807
rect 11692 31807 11750 31813
rect 9622 31776 9720 31804
rect 9622 31773 9634 31776
rect 9576 31767 9634 31773
rect 9692 31748 9720 31776
rect 11692 31773 11704 31807
rect 11738 31804 11750 31807
rect 12802 31804 12808 31816
rect 11738 31776 12808 31804
rect 11738 31773 11750 31776
rect 11692 31767 11750 31773
rect 12802 31764 12808 31776
rect 12860 31764 12866 31816
rect 16666 31764 16672 31816
rect 16724 31804 16730 31816
rect 17497 31807 17555 31813
rect 17497 31804 17509 31807
rect 16724 31776 17509 31804
rect 16724 31764 16730 31776
rect 17497 31773 17509 31776
rect 17543 31773 17555 31807
rect 17497 31767 17555 31773
rect 22094 31764 22100 31816
rect 22152 31804 22158 31816
rect 23845 31807 23903 31813
rect 23845 31804 23857 31807
rect 22152 31776 22197 31804
rect 23676 31776 23857 31804
rect 22152 31764 22158 31776
rect 23676 31748 23704 31776
rect 23845 31773 23857 31776
rect 23891 31773 23903 31807
rect 25222 31804 25228 31816
rect 25183 31776 25228 31804
rect 23845 31767 23903 31773
rect 25222 31764 25228 31776
rect 25280 31764 25286 31816
rect 30834 31764 30840 31816
rect 30892 31813 30898 31816
rect 30892 31804 30904 31813
rect 31113 31807 31171 31813
rect 30892 31776 30937 31804
rect 30892 31767 30904 31776
rect 31113 31773 31125 31807
rect 31159 31804 31171 31807
rect 32306 31804 32312 31816
rect 31159 31776 32312 31804
rect 31159 31773 31171 31776
rect 31113 31767 31171 31773
rect 30892 31764 30898 31767
rect 32306 31764 32312 31776
rect 32364 31764 32370 31816
rect 36087 31807 36145 31813
rect 36087 31773 36099 31807
rect 36133 31773 36145 31807
rect 36262 31804 36268 31816
rect 36223 31776 36268 31804
rect 36087 31767 36145 31773
rect 2774 31736 2780 31748
rect 2608 31708 2780 31736
rect 2774 31696 2780 31708
rect 2832 31696 2838 31748
rect 5626 31696 5632 31748
rect 5684 31736 5690 31748
rect 7929 31739 7987 31745
rect 7929 31736 7941 31739
rect 5684 31708 7941 31736
rect 5684 31696 5690 31708
rect 7929 31705 7941 31708
rect 7975 31705 7987 31739
rect 8110 31736 8116 31748
rect 8071 31708 8116 31736
rect 7929 31699 7987 31705
rect 8110 31696 8116 31708
rect 8168 31696 8174 31748
rect 9674 31696 9680 31748
rect 9732 31696 9738 31748
rect 22279 31739 22337 31745
rect 22279 31705 22291 31739
rect 22325 31736 22337 31739
rect 22325 31708 22600 31736
rect 22325 31705 22337 31708
rect 22279 31699 22337 31705
rect 3237 31671 3295 31677
rect 3237 31668 3249 31671
rect 2312 31640 3249 31668
rect 3237 31637 3249 31640
rect 3283 31668 3295 31671
rect 3326 31668 3332 31680
rect 3283 31640 3332 31668
rect 3283 31637 3295 31640
rect 3237 31631 3295 31637
rect 3326 31628 3332 31640
rect 3384 31628 3390 31680
rect 12805 31671 12863 31677
rect 12805 31637 12817 31671
rect 12851 31668 12863 31671
rect 12894 31668 12900 31680
rect 12851 31640 12900 31668
rect 12851 31637 12863 31640
rect 12805 31631 12863 31637
rect 12894 31628 12900 31640
rect 12952 31628 12958 31680
rect 22462 31668 22468 31680
rect 22423 31640 22468 31668
rect 22462 31628 22468 31640
rect 22520 31628 22526 31680
rect 22572 31668 22600 31708
rect 22646 31696 22652 31748
rect 22704 31736 22710 31748
rect 22830 31736 22836 31748
rect 22704 31708 22836 31736
rect 22704 31696 22710 31708
rect 22830 31696 22836 31708
rect 22888 31696 22894 31748
rect 23658 31696 23664 31748
rect 23716 31696 23722 31748
rect 35986 31696 35992 31748
rect 36044 31736 36050 31748
rect 36096 31736 36124 31767
rect 36262 31764 36268 31776
rect 36320 31764 36326 31816
rect 36357 31807 36415 31813
rect 36357 31773 36369 31807
rect 36403 31773 36415 31807
rect 36357 31767 36415 31773
rect 36044 31708 36124 31736
rect 36044 31696 36050 31708
rect 36170 31696 36176 31748
rect 36228 31736 36234 31748
rect 36372 31736 36400 31767
rect 36446 31764 36452 31816
rect 36504 31813 36510 31816
rect 36504 31807 36553 31813
rect 36504 31773 36507 31807
rect 36541 31773 36553 31807
rect 36740 31804 36768 31835
rect 37550 31832 37556 31844
rect 37608 31832 37614 31884
rect 37809 31807 37867 31813
rect 37809 31804 37821 31807
rect 36740 31776 37821 31804
rect 36504 31767 36553 31773
rect 37809 31773 37821 31776
rect 37855 31773 37867 31807
rect 37809 31767 37867 31773
rect 36504 31764 36510 31767
rect 36228 31708 36400 31736
rect 36228 31696 36234 31708
rect 22922 31668 22928 31680
rect 22572 31640 22928 31668
rect 22922 31628 22928 31640
rect 22980 31628 22986 31680
rect 38930 31668 38936 31680
rect 38891 31640 38936 31668
rect 38930 31628 38936 31640
rect 38988 31628 38994 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 2409 31467 2467 31473
rect 2409 31433 2421 31467
rect 2455 31464 2467 31467
rect 2774 31464 2780 31476
rect 2455 31436 2780 31464
rect 2455 31433 2467 31436
rect 2409 31427 2467 31433
rect 2774 31424 2780 31436
rect 2832 31424 2838 31476
rect 5169 31467 5227 31473
rect 5169 31433 5181 31467
rect 5215 31464 5227 31467
rect 5258 31464 5264 31476
rect 5215 31436 5264 31464
rect 5215 31433 5227 31436
rect 5169 31427 5227 31433
rect 5258 31424 5264 31436
rect 5316 31424 5322 31476
rect 5626 31464 5632 31476
rect 5587 31436 5632 31464
rect 5626 31424 5632 31436
rect 5684 31424 5690 31476
rect 7282 31424 7288 31476
rect 7340 31464 7346 31476
rect 9125 31467 9183 31473
rect 9125 31464 9137 31467
rect 7340 31436 9137 31464
rect 7340 31424 7346 31436
rect 9125 31433 9137 31436
rect 9171 31433 9183 31467
rect 9674 31464 9680 31476
rect 9635 31436 9680 31464
rect 9125 31427 9183 31433
rect 9674 31424 9680 31436
rect 9732 31424 9738 31476
rect 10226 31464 10232 31476
rect 9876 31436 10232 31464
rect 2593 31399 2651 31405
rect 2593 31365 2605 31399
rect 2639 31396 2651 31399
rect 3602 31396 3608 31408
rect 2639 31368 3608 31396
rect 2639 31365 2651 31368
rect 2593 31359 2651 31365
rect 3602 31356 3608 31368
rect 3660 31356 3666 31408
rect 4062 31356 4068 31408
rect 4120 31396 4126 31408
rect 4120 31368 6684 31396
rect 4120 31356 4126 31368
rect 2774 31288 2780 31340
rect 2832 31328 2838 31340
rect 6656 31337 6684 31368
rect 6822 31356 6828 31408
rect 6880 31396 6886 31408
rect 8389 31399 8447 31405
rect 8389 31396 8401 31399
rect 6880 31368 8401 31396
rect 6880 31356 6886 31368
rect 5813 31331 5871 31337
rect 2832 31300 2877 31328
rect 2832 31288 2838 31300
rect 5813 31297 5825 31331
rect 5859 31297 5871 31331
rect 5813 31291 5871 31297
rect 6641 31331 6699 31337
rect 6641 31297 6653 31331
rect 6687 31328 6699 31331
rect 7098 31328 7104 31340
rect 6687 31300 7104 31328
rect 6687 31297 6699 31300
rect 6641 31291 6699 31297
rect 5828 31192 5856 31291
rect 7098 31288 7104 31300
rect 7156 31288 7162 31340
rect 7392 31337 7420 31368
rect 8389 31365 8401 31368
rect 8435 31365 8447 31399
rect 8389 31359 8447 31365
rect 8573 31399 8631 31405
rect 8573 31365 8585 31399
rect 8619 31396 8631 31399
rect 9876 31396 9904 31436
rect 10226 31424 10232 31436
rect 10284 31424 10290 31476
rect 10870 31464 10876 31476
rect 10831 31436 10876 31464
rect 10870 31424 10876 31436
rect 10928 31424 10934 31476
rect 12802 31424 12808 31476
rect 12860 31464 12866 31476
rect 12897 31467 12955 31473
rect 12897 31464 12909 31467
rect 12860 31436 12909 31464
rect 12860 31424 12866 31436
rect 12897 31433 12909 31436
rect 12943 31433 12955 31467
rect 12897 31427 12955 31433
rect 13262 31424 13268 31476
rect 13320 31424 13326 31476
rect 16298 31424 16304 31476
rect 16356 31464 16362 31476
rect 24394 31464 24400 31476
rect 16356 31436 24400 31464
rect 16356 31424 16362 31436
rect 24394 31424 24400 31436
rect 24452 31464 24458 31476
rect 24452 31436 27614 31464
rect 24452 31424 24458 31436
rect 10888 31396 10916 31424
rect 8619 31368 9904 31396
rect 9968 31368 10916 31396
rect 8619 31365 8631 31368
rect 8573 31359 8631 31365
rect 7285 31331 7343 31337
rect 7285 31297 7297 31331
rect 7331 31297 7343 31331
rect 7285 31291 7343 31297
rect 7377 31331 7435 31337
rect 7377 31297 7389 31331
rect 7423 31297 7435 31331
rect 7377 31291 7435 31297
rect 5902 31220 5908 31272
rect 5960 31260 5966 31272
rect 7300 31260 7328 31291
rect 7466 31288 7472 31340
rect 7524 31328 7530 31340
rect 9968 31337 9996 31368
rect 9953 31331 10011 31337
rect 7524 31300 7569 31328
rect 7524 31288 7530 31300
rect 9953 31297 9965 31331
rect 9999 31297 10011 31331
rect 9953 31291 10011 31297
rect 10045 31331 10103 31337
rect 10045 31297 10057 31331
rect 10091 31297 10103 31331
rect 10045 31291 10103 31297
rect 5960 31232 7328 31260
rect 7484 31260 7512 31288
rect 8570 31260 8576 31272
rect 7484 31232 8576 31260
rect 5960 31220 5966 31232
rect 8570 31220 8576 31232
rect 8628 31220 8634 31272
rect 9582 31220 9588 31272
rect 9640 31260 9646 31272
rect 10060 31260 10088 31291
rect 10134 31288 10140 31340
rect 10192 31328 10198 31340
rect 10321 31331 10379 31337
rect 10192 31300 10237 31328
rect 10192 31288 10198 31300
rect 10321 31297 10333 31331
rect 10367 31328 10379 31331
rect 10778 31328 10784 31340
rect 10367 31300 10784 31328
rect 10367 31297 10379 31300
rect 10321 31291 10379 31297
rect 10778 31288 10784 31300
rect 10836 31288 10842 31340
rect 11698 31328 11704 31340
rect 11659 31300 11704 31328
rect 11698 31288 11704 31300
rect 11756 31288 11762 31340
rect 11882 31328 11888 31340
rect 11843 31300 11888 31328
rect 11882 31288 11888 31300
rect 11940 31288 11946 31340
rect 13280 31337 13308 31424
rect 23385 31399 23443 31405
rect 23385 31396 23397 31399
rect 15120 31368 15792 31396
rect 13173 31331 13231 31337
rect 13173 31297 13185 31331
rect 13219 31297 13231 31331
rect 13173 31291 13231 31297
rect 13262 31331 13320 31337
rect 13262 31297 13274 31331
rect 13308 31297 13320 31331
rect 13262 31291 13320 31297
rect 9640 31232 10088 31260
rect 13188 31260 13216 31291
rect 13354 31288 13360 31340
rect 13412 31328 13418 31340
rect 13541 31331 13599 31337
rect 13412 31300 13457 31328
rect 13412 31288 13418 31300
rect 13541 31297 13553 31331
rect 13587 31328 13599 31331
rect 13722 31328 13728 31340
rect 13587 31300 13728 31328
rect 13587 31297 13599 31300
rect 13541 31291 13599 31297
rect 13722 31288 13728 31300
rect 13780 31288 13786 31340
rect 14274 31288 14280 31340
rect 14332 31328 14338 31340
rect 15120 31337 15148 31368
rect 15105 31331 15163 31337
rect 15105 31328 15117 31331
rect 14332 31300 15117 31328
rect 14332 31288 14338 31300
rect 15105 31297 15117 31300
rect 15151 31297 15163 31331
rect 15105 31291 15163 31297
rect 15197 31331 15255 31337
rect 15197 31297 15209 31331
rect 15243 31297 15255 31331
rect 15197 31291 15255 31297
rect 15289 31331 15347 31337
rect 15289 31297 15301 31331
rect 15335 31297 15347 31331
rect 15289 31291 15347 31297
rect 15473 31331 15531 31337
rect 15473 31297 15485 31331
rect 15519 31328 15531 31331
rect 15654 31328 15660 31340
rect 15519 31300 15660 31328
rect 15519 31297 15531 31300
rect 15473 31291 15531 31297
rect 14292 31260 14320 31288
rect 13188 31232 14320 31260
rect 9640 31220 9646 31232
rect 15010 31220 15016 31272
rect 15068 31260 15074 31272
rect 15212 31260 15240 31291
rect 15068 31232 15240 31260
rect 15068 31220 15074 31232
rect 13170 31192 13176 31204
rect 5828 31164 13176 31192
rect 13170 31152 13176 31164
rect 13228 31152 13234 31204
rect 7650 31084 7656 31136
rect 7708 31124 7714 31136
rect 7745 31127 7803 31133
rect 7745 31124 7757 31127
rect 7708 31096 7757 31124
rect 7708 31084 7714 31096
rect 7745 31093 7757 31096
rect 7791 31093 7803 31127
rect 7745 31087 7803 31093
rect 10410 31084 10416 31136
rect 10468 31124 10474 31136
rect 11517 31127 11575 31133
rect 11517 31124 11529 31127
rect 10468 31096 11529 31124
rect 10468 31084 10474 31096
rect 11517 31093 11529 31096
rect 11563 31093 11575 31127
rect 11517 31087 11575 31093
rect 12434 31084 12440 31136
rect 12492 31124 12498 31136
rect 12492 31096 12537 31124
rect 12492 31084 12498 31096
rect 13722 31084 13728 31136
rect 13780 31124 13786 31136
rect 14001 31127 14059 31133
rect 14001 31124 14013 31127
rect 13780 31096 14013 31124
rect 13780 31084 13786 31096
rect 14001 31093 14013 31096
rect 14047 31093 14059 31127
rect 14001 31087 14059 31093
rect 14829 31127 14887 31133
rect 14829 31093 14841 31127
rect 14875 31124 14887 31127
rect 14918 31124 14924 31136
rect 14875 31096 14924 31124
rect 14875 31093 14887 31096
rect 14829 31087 14887 31093
rect 14918 31084 14924 31096
rect 14976 31084 14982 31136
rect 15212 31124 15240 31232
rect 15304 31192 15332 31291
rect 15654 31288 15660 31300
rect 15712 31288 15718 31340
rect 15470 31192 15476 31204
rect 15304 31164 15476 31192
rect 15470 31152 15476 31164
rect 15528 31152 15534 31204
rect 15562 31124 15568 31136
rect 15212 31096 15568 31124
rect 15562 31084 15568 31096
rect 15620 31084 15626 31136
rect 15764 31124 15792 31368
rect 23124 31368 23397 31396
rect 19426 31288 19432 31340
rect 19484 31328 19490 31340
rect 19777 31331 19835 31337
rect 19777 31328 19789 31331
rect 19484 31300 19789 31328
rect 19484 31288 19490 31300
rect 19777 31297 19789 31300
rect 19823 31297 19835 31331
rect 22276 31328 22282 31340
rect 22239 31300 22282 31328
rect 19777 31291 19835 31297
rect 22276 31288 22282 31300
rect 22334 31288 22340 31340
rect 22373 31331 22431 31337
rect 22373 31297 22385 31331
rect 22419 31297 22431 31331
rect 22373 31291 22431 31297
rect 19242 31220 19248 31272
rect 19300 31260 19306 31272
rect 19521 31263 19579 31269
rect 19521 31260 19533 31263
rect 19300 31232 19533 31260
rect 19300 31220 19306 31232
rect 19521 31229 19533 31232
rect 19567 31229 19579 31263
rect 19521 31223 19579 31229
rect 20806 31220 20812 31272
rect 20864 31260 20870 31272
rect 22388 31260 22416 31291
rect 22462 31288 22468 31340
rect 22520 31337 22526 31340
rect 22520 31328 22528 31337
rect 22649 31331 22707 31337
rect 22520 31300 22565 31328
rect 22520 31291 22528 31300
rect 22649 31297 22661 31331
rect 22695 31297 22707 31331
rect 22649 31291 22707 31297
rect 22520 31288 22526 31291
rect 20864 31232 22416 31260
rect 20864 31220 20870 31232
rect 22554 31220 22560 31272
rect 22612 31260 22618 31272
rect 22664 31260 22692 31291
rect 22612 31232 22692 31260
rect 22612 31220 22618 31232
rect 15930 31152 15936 31204
rect 15988 31192 15994 31204
rect 23124 31192 23152 31368
rect 23385 31365 23397 31368
rect 23431 31396 23443 31399
rect 24302 31396 24308 31408
rect 23431 31368 24308 31396
rect 23431 31365 23443 31368
rect 23385 31359 23443 31365
rect 24302 31356 24308 31368
rect 24360 31356 24366 31408
rect 27586 31396 27614 31436
rect 29546 31424 29552 31476
rect 29604 31464 29610 31476
rect 29914 31464 29920 31476
rect 29604 31436 29920 31464
rect 29604 31424 29610 31436
rect 29914 31424 29920 31436
rect 29972 31424 29978 31476
rect 30377 31467 30435 31473
rect 30377 31433 30389 31467
rect 30423 31464 30435 31467
rect 32214 31464 32220 31476
rect 30423 31436 32220 31464
rect 30423 31433 30435 31436
rect 30377 31427 30435 31433
rect 32214 31424 32220 31436
rect 32272 31424 32278 31476
rect 36173 31467 36231 31473
rect 36173 31433 36185 31467
rect 36219 31464 36231 31467
rect 36262 31464 36268 31476
rect 36219 31436 36268 31464
rect 36219 31433 36231 31436
rect 36173 31427 36231 31433
rect 36262 31424 36268 31436
rect 36320 31424 36326 31476
rect 30926 31396 30932 31408
rect 27586 31368 30932 31396
rect 30926 31356 30932 31368
rect 30984 31356 30990 31408
rect 31110 31396 31116 31408
rect 31071 31368 31116 31396
rect 31110 31356 31116 31368
rect 31168 31356 31174 31408
rect 33594 31356 33600 31408
rect 33652 31396 33658 31408
rect 35989 31399 36047 31405
rect 35989 31396 36001 31399
rect 33652 31368 36001 31396
rect 33652 31356 33658 31368
rect 35989 31365 36001 31368
rect 36035 31396 36047 31399
rect 38930 31396 38936 31408
rect 36035 31368 38936 31396
rect 36035 31365 36047 31368
rect 35989 31359 36047 31365
rect 38930 31356 38936 31368
rect 38988 31356 38994 31408
rect 23201 31331 23259 31337
rect 23201 31297 23213 31331
rect 23247 31328 23259 31331
rect 23658 31328 23664 31340
rect 23247 31300 23664 31328
rect 23247 31297 23259 31300
rect 23201 31291 23259 31297
rect 23658 31288 23664 31300
rect 23716 31288 23722 31340
rect 29914 31288 29920 31340
rect 29972 31328 29978 31340
rect 30190 31328 30196 31340
rect 29972 31300 30196 31328
rect 29972 31288 29978 31300
rect 30190 31288 30196 31300
rect 30248 31288 30254 31340
rect 30374 31288 30380 31340
rect 30432 31328 30438 31340
rect 31021 31331 31079 31337
rect 31021 31328 31033 31331
rect 30432 31300 31033 31328
rect 30432 31288 30438 31300
rect 31021 31297 31033 31300
rect 31067 31297 31079 31331
rect 31202 31328 31208 31340
rect 31163 31300 31208 31328
rect 31021 31291 31079 31297
rect 30009 31263 30067 31269
rect 30009 31260 30021 31263
rect 15988 31164 19104 31192
rect 15988 31152 15994 31164
rect 16025 31127 16083 31133
rect 16025 31124 16037 31127
rect 15764 31096 16037 31124
rect 16025 31093 16037 31096
rect 16071 31124 16083 31127
rect 16298 31124 16304 31136
rect 16071 31096 16304 31124
rect 16071 31093 16083 31096
rect 16025 31087 16083 31093
rect 16298 31084 16304 31096
rect 16356 31084 16362 31136
rect 18782 31084 18788 31136
rect 18840 31124 18846 31136
rect 18969 31127 19027 31133
rect 18969 31124 18981 31127
rect 18840 31096 18981 31124
rect 18840 31084 18846 31096
rect 18969 31093 18981 31096
rect 19015 31093 19027 31127
rect 19076 31124 19104 31164
rect 20456 31164 23152 31192
rect 29472 31232 30021 31260
rect 20456 31124 20484 31164
rect 29472 31136 29500 31232
rect 30009 31229 30021 31232
rect 30055 31229 30067 31263
rect 31036 31260 31064 31291
rect 31202 31288 31208 31300
rect 31260 31288 31266 31340
rect 31386 31328 31392 31340
rect 31347 31300 31392 31328
rect 31386 31288 31392 31300
rect 31444 31288 31450 31340
rect 32309 31331 32367 31337
rect 32309 31297 32321 31331
rect 32355 31328 32367 31331
rect 33134 31328 33140 31340
rect 32355 31300 33140 31328
rect 32355 31297 32367 31300
rect 32309 31291 32367 31297
rect 33134 31288 33140 31300
rect 33192 31288 33198 31340
rect 35342 31288 35348 31340
rect 35400 31328 35406 31340
rect 35805 31331 35863 31337
rect 35805 31328 35817 31331
rect 35400 31300 35817 31328
rect 35400 31288 35406 31300
rect 35805 31297 35817 31300
rect 35851 31328 35863 31331
rect 37274 31328 37280 31340
rect 35851 31300 37280 31328
rect 35851 31297 35863 31300
rect 35805 31291 35863 31297
rect 37274 31288 37280 31300
rect 37332 31288 37338 31340
rect 33502 31260 33508 31272
rect 31036 31232 33508 31260
rect 30009 31223 30067 31229
rect 33502 31220 33508 31232
rect 33560 31220 33566 31272
rect 30098 31152 30104 31204
rect 30156 31192 30162 31204
rect 32125 31195 32183 31201
rect 32125 31192 32137 31195
rect 30156 31164 32137 31192
rect 30156 31152 30162 31164
rect 32125 31161 32137 31164
rect 32171 31161 32183 31195
rect 32125 31155 32183 31161
rect 20898 31124 20904 31136
rect 19076 31096 20484 31124
rect 20859 31096 20904 31124
rect 18969 31087 19027 31093
rect 20898 31084 20904 31096
rect 20956 31084 20962 31136
rect 22002 31124 22008 31136
rect 21963 31096 22008 31124
rect 22002 31084 22008 31096
rect 22060 31084 22066 31136
rect 23658 31084 23664 31136
rect 23716 31124 23722 31136
rect 23937 31127 23995 31133
rect 23937 31124 23949 31127
rect 23716 31096 23949 31124
rect 23716 31084 23722 31096
rect 23937 31093 23949 31096
rect 23983 31093 23995 31127
rect 23937 31087 23995 31093
rect 25041 31127 25099 31133
rect 25041 31093 25053 31127
rect 25087 31124 25099 31127
rect 25406 31124 25412 31136
rect 25087 31096 25412 31124
rect 25087 31093 25099 31096
rect 25041 31087 25099 31093
rect 25406 31084 25412 31096
rect 25464 31084 25470 31136
rect 29454 31124 29460 31136
rect 29415 31096 29460 31124
rect 29454 31084 29460 31096
rect 29512 31084 29518 31136
rect 30837 31127 30895 31133
rect 30837 31093 30849 31127
rect 30883 31124 30895 31127
rect 31018 31124 31024 31136
rect 30883 31096 31024 31124
rect 30883 31093 30895 31096
rect 30837 31087 30895 31093
rect 31018 31084 31024 31096
rect 31076 31084 31082 31136
rect 31110 31084 31116 31136
rect 31168 31124 31174 31136
rect 31938 31124 31944 31136
rect 31168 31096 31944 31124
rect 31168 31084 31174 31096
rect 31938 31084 31944 31096
rect 31996 31084 32002 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 5902 30920 5908 30932
rect 5863 30892 5908 30920
rect 5902 30880 5908 30892
rect 5960 30880 5966 30932
rect 6365 30923 6423 30929
rect 6365 30889 6377 30923
rect 6411 30920 6423 30923
rect 6454 30920 6460 30932
rect 6411 30892 6460 30920
rect 6411 30889 6423 30892
rect 6365 30883 6423 30889
rect 6454 30880 6460 30892
rect 6512 30880 6518 30932
rect 7926 30880 7932 30932
rect 7984 30920 7990 30932
rect 8021 30923 8079 30929
rect 8021 30920 8033 30923
rect 7984 30892 8033 30920
rect 7984 30880 7990 30892
rect 8021 30889 8033 30892
rect 8067 30889 8079 30923
rect 8021 30883 8079 30889
rect 11790 30880 11796 30932
rect 11848 30920 11854 30932
rect 11885 30923 11943 30929
rect 11885 30920 11897 30923
rect 11848 30892 11897 30920
rect 11848 30880 11854 30892
rect 11885 30889 11897 30892
rect 11931 30920 11943 30923
rect 17034 30920 17040 30932
rect 11931 30892 17040 30920
rect 11931 30889 11943 30892
rect 11885 30883 11943 30889
rect 17034 30880 17040 30892
rect 17092 30920 17098 30932
rect 20254 30920 20260 30932
rect 17092 30892 20260 30920
rect 17092 30880 17098 30892
rect 20254 30880 20260 30892
rect 20312 30880 20318 30932
rect 29546 30920 29552 30932
rect 20364 30892 29552 30920
rect 6822 30852 6828 30864
rect 6656 30824 6828 30852
rect 6656 30784 6684 30824
rect 6822 30812 6828 30824
rect 6880 30812 6886 30864
rect 9033 30855 9091 30861
rect 9033 30852 9045 30855
rect 7668 30824 9045 30852
rect 7558 30784 7564 30796
rect 6656 30756 6776 30784
rect 2593 30719 2651 30725
rect 2593 30685 2605 30719
rect 2639 30716 2651 30719
rect 3786 30716 3792 30728
rect 2639 30688 3792 30716
rect 2639 30685 2651 30688
rect 2593 30679 2651 30685
rect 3786 30676 3792 30688
rect 3844 30676 3850 30728
rect 5537 30719 5595 30725
rect 5537 30685 5549 30719
rect 5583 30716 5595 30719
rect 5626 30716 5632 30728
rect 5583 30688 5632 30716
rect 5583 30685 5595 30688
rect 5537 30679 5595 30685
rect 5626 30676 5632 30688
rect 5684 30676 5690 30728
rect 6638 30716 6644 30728
rect 6551 30688 6644 30716
rect 6638 30676 6644 30688
rect 6696 30676 6702 30728
rect 6748 30725 6776 30756
rect 6840 30756 7564 30784
rect 6840 30725 6868 30756
rect 7558 30744 7564 30756
rect 7616 30744 7622 30796
rect 6733 30719 6791 30725
rect 6733 30685 6745 30719
rect 6779 30685 6791 30719
rect 6733 30679 6791 30685
rect 6825 30719 6883 30725
rect 6825 30685 6837 30719
rect 6871 30685 6883 30719
rect 6825 30679 6883 30685
rect 7009 30719 7067 30725
rect 7009 30685 7021 30719
rect 7055 30716 7067 30719
rect 7098 30716 7104 30728
rect 7055 30688 7104 30716
rect 7055 30685 7067 30688
rect 7009 30679 7067 30685
rect 7098 30676 7104 30688
rect 7156 30716 7162 30728
rect 7668 30716 7696 30824
rect 9033 30821 9045 30824
rect 9079 30852 9091 30855
rect 14185 30855 14243 30861
rect 9079 30824 14044 30852
rect 9079 30821 9091 30824
rect 9033 30815 9091 30821
rect 9674 30784 9680 30796
rect 8128 30756 9680 30784
rect 8128 30725 8156 30756
rect 9674 30744 9680 30756
rect 9732 30784 9738 30796
rect 13446 30784 13452 30796
rect 9732 30756 13452 30784
rect 9732 30744 9738 30756
rect 13446 30744 13452 30756
rect 13504 30744 13510 30796
rect 7156 30688 7696 30716
rect 8113 30719 8171 30725
rect 7156 30676 7162 30688
rect 8113 30685 8125 30719
rect 8159 30685 8171 30719
rect 8113 30679 8171 30685
rect 11054 30676 11060 30728
rect 11112 30716 11118 30728
rect 12621 30719 12679 30725
rect 12621 30716 12633 30719
rect 11112 30688 12633 30716
rect 11112 30676 11118 30688
rect 12621 30685 12633 30688
rect 12667 30685 12679 30719
rect 12894 30716 12900 30728
rect 12855 30688 12900 30716
rect 12621 30679 12679 30685
rect 12894 30676 12900 30688
rect 12952 30676 12958 30728
rect 12986 30676 12992 30728
rect 13044 30725 13050 30728
rect 13044 30719 13071 30725
rect 13059 30685 13071 30719
rect 13044 30679 13071 30685
rect 13044 30676 13050 30679
rect 2774 30608 2780 30660
rect 2832 30648 2838 30660
rect 4890 30648 4896 30660
rect 2832 30620 4896 30648
rect 2832 30608 2838 30620
rect 4890 30608 4896 30620
rect 4948 30608 4954 30660
rect 5721 30651 5779 30657
rect 5721 30617 5733 30651
rect 5767 30648 5779 30651
rect 6270 30648 6276 30660
rect 5767 30620 6276 30648
rect 5767 30617 5779 30620
rect 5721 30611 5779 30617
rect 6270 30608 6276 30620
rect 6328 30608 6334 30660
rect 6656 30648 6684 30676
rect 6914 30648 6920 30660
rect 6656 30620 6920 30648
rect 6914 30608 6920 30620
rect 6972 30608 6978 30660
rect 10413 30651 10471 30657
rect 10413 30617 10425 30651
rect 10459 30648 10471 30651
rect 12434 30648 12440 30660
rect 10459 30620 12440 30648
rect 10459 30617 10471 30620
rect 10413 30611 10471 30617
rect 12434 30608 12440 30620
rect 12492 30608 12498 30660
rect 12526 30608 12532 30660
rect 12584 30648 12590 30660
rect 12805 30651 12863 30657
rect 12805 30648 12817 30651
rect 12584 30620 12817 30648
rect 12584 30608 12590 30620
rect 12805 30617 12817 30620
rect 12851 30617 12863 30651
rect 14016 30648 14044 30824
rect 14185 30821 14197 30855
rect 14231 30852 14243 30855
rect 14274 30852 14280 30864
rect 14231 30824 14280 30852
rect 14231 30821 14243 30824
rect 14185 30815 14243 30821
rect 14274 30812 14280 30824
rect 14332 30812 14338 30864
rect 16758 30812 16764 30864
rect 16816 30852 16822 30864
rect 17310 30852 17316 30864
rect 16816 30824 17316 30852
rect 16816 30812 16822 30824
rect 17310 30812 17316 30824
rect 17368 30812 17374 30864
rect 18322 30812 18328 30864
rect 18380 30852 18386 30864
rect 19242 30852 19248 30864
rect 18380 30824 19248 30852
rect 18380 30812 18386 30824
rect 19242 30812 19248 30824
rect 19300 30812 19306 30864
rect 14090 30744 14096 30796
rect 14148 30784 14154 30796
rect 14826 30784 14832 30796
rect 14148 30756 14832 30784
rect 14148 30744 14154 30756
rect 14826 30744 14832 30756
rect 14884 30744 14890 30796
rect 20364 30784 20392 30892
rect 29546 30880 29552 30892
rect 29604 30920 29610 30932
rect 29641 30923 29699 30929
rect 29641 30920 29653 30923
rect 29604 30892 29653 30920
rect 29604 30880 29610 30892
rect 29641 30889 29653 30892
rect 29687 30889 29699 30923
rect 29641 30883 29699 30889
rect 24394 30852 24400 30864
rect 24355 30824 24400 30852
rect 24394 30812 24400 30824
rect 24452 30852 24458 30864
rect 24452 30824 25445 30852
rect 24452 30812 24458 30824
rect 15856 30756 20392 30784
rect 14918 30676 14924 30728
rect 14976 30716 14982 30728
rect 15085 30719 15143 30725
rect 15085 30716 15097 30719
rect 14976 30688 15097 30716
rect 14976 30676 14982 30688
rect 15085 30685 15097 30688
rect 15131 30685 15143 30719
rect 15085 30679 15143 30685
rect 15856 30648 15884 30756
rect 16482 30676 16488 30728
rect 16540 30716 16546 30728
rect 16853 30719 16911 30725
rect 16853 30716 16865 30719
rect 16540 30688 16865 30716
rect 16540 30676 16546 30688
rect 16853 30685 16865 30688
rect 16899 30685 16911 30719
rect 17034 30716 17040 30728
rect 16995 30688 17040 30716
rect 16853 30679 16911 30685
rect 17034 30676 17040 30688
rect 17092 30676 17098 30728
rect 19705 30719 19763 30725
rect 19705 30716 19717 30719
rect 18340 30688 19717 30716
rect 16666 30648 16672 30660
rect 14016 30620 15884 30648
rect 15939 30620 16672 30648
rect 12805 30611 12863 30617
rect 2409 30583 2467 30589
rect 2409 30549 2421 30583
rect 2455 30580 2467 30583
rect 2590 30580 2596 30592
rect 2455 30552 2596 30580
rect 2455 30549 2467 30552
rect 2409 30543 2467 30549
rect 2590 30540 2596 30552
rect 2648 30540 2654 30592
rect 13173 30583 13231 30589
rect 13173 30549 13185 30583
rect 13219 30580 13231 30583
rect 13998 30580 14004 30592
rect 13219 30552 14004 30580
rect 13219 30549 13231 30552
rect 13173 30543 13231 30549
rect 13998 30540 14004 30552
rect 14056 30540 14062 30592
rect 14918 30540 14924 30592
rect 14976 30580 14982 30592
rect 15939 30580 15967 30620
rect 16666 30608 16672 30620
rect 16724 30608 16730 30660
rect 18340 30657 18368 30688
rect 19705 30685 19717 30688
rect 19751 30716 19763 30719
rect 20257 30719 20315 30725
rect 20257 30716 20269 30719
rect 19751 30688 20269 30716
rect 19751 30685 19763 30688
rect 19705 30679 19763 30685
rect 20257 30685 20269 30688
rect 20303 30716 20315 30719
rect 20438 30716 20444 30728
rect 20303 30688 20444 30716
rect 20303 30685 20315 30688
rect 20257 30679 20315 30685
rect 20438 30676 20444 30688
rect 20496 30676 20502 30728
rect 20533 30719 20591 30725
rect 20533 30685 20545 30719
rect 20579 30685 20591 30719
rect 21726 30716 21732 30728
rect 21687 30688 21732 30716
rect 20533 30679 20591 30685
rect 18325 30651 18383 30657
rect 18325 30617 18337 30651
rect 18371 30617 18383 30651
rect 18506 30648 18512 30660
rect 18467 30620 18512 30648
rect 18325 30611 18383 30617
rect 16206 30580 16212 30592
rect 14976 30552 15967 30580
rect 16167 30552 16212 30580
rect 14976 30540 14982 30552
rect 16206 30540 16212 30552
rect 16264 30540 16270 30592
rect 17310 30540 17316 30592
rect 17368 30580 17374 30592
rect 17773 30583 17831 30589
rect 17773 30580 17785 30583
rect 17368 30552 17785 30580
rect 17368 30540 17374 30552
rect 17773 30549 17785 30552
rect 17819 30580 17831 30583
rect 18340 30580 18368 30611
rect 18506 30608 18512 30620
rect 18564 30608 18570 30660
rect 20548 30648 20576 30679
rect 21726 30676 21732 30688
rect 21784 30676 21790 30728
rect 22002 30725 22008 30728
rect 21996 30716 22008 30725
rect 21963 30688 22008 30716
rect 21996 30679 22008 30688
rect 22002 30676 22008 30679
rect 22060 30676 22066 30728
rect 24670 30676 24676 30728
rect 24728 30716 24734 30728
rect 24949 30719 25007 30725
rect 24949 30716 24961 30719
rect 24728 30688 24961 30716
rect 24728 30676 24734 30688
rect 24949 30685 24961 30688
rect 24995 30685 25007 30719
rect 25130 30716 25136 30728
rect 25091 30688 25136 30716
rect 24949 30679 25007 30685
rect 25130 30676 25136 30688
rect 25188 30676 25194 30728
rect 25231 30676 25237 30728
rect 25289 30725 25295 30728
rect 25417 30725 25445 30824
rect 25593 30787 25651 30793
rect 25593 30753 25605 30787
rect 25639 30784 25651 30787
rect 27522 30784 27528 30796
rect 25639 30756 26464 30784
rect 27483 30756 27528 30784
rect 25639 30753 25651 30756
rect 25593 30747 25651 30753
rect 25289 30719 25302 30725
rect 25290 30716 25302 30719
rect 25363 30719 25445 30725
rect 25290 30688 25334 30716
rect 25290 30685 25302 30688
rect 25289 30679 25302 30685
rect 25363 30685 25375 30719
rect 25409 30688 25445 30719
rect 26436 30716 26464 30756
rect 27522 30744 27528 30756
rect 27580 30744 27586 30796
rect 29656 30784 29684 30883
rect 30926 30880 30932 30932
rect 30984 30920 30990 30932
rect 33778 30920 33784 30932
rect 30984 30892 33784 30920
rect 30984 30880 30990 30892
rect 33778 30880 33784 30892
rect 33836 30880 33842 30932
rect 39301 30923 39359 30929
rect 39301 30920 39313 30923
rect 35268 30892 39313 30920
rect 29656 30756 31248 30784
rect 27258 30719 27316 30725
rect 27258 30716 27270 30719
rect 26436 30688 27270 30716
rect 25409 30685 25421 30688
rect 25363 30679 25421 30685
rect 27258 30685 27270 30688
rect 27304 30685 27316 30719
rect 30374 30716 30380 30728
rect 30335 30688 30380 30716
rect 27258 30679 27316 30685
rect 25289 30676 25295 30679
rect 30374 30676 30380 30688
rect 30432 30676 30438 30728
rect 30745 30719 30803 30725
rect 30745 30685 30757 30719
rect 30791 30716 30803 30719
rect 31110 30716 31116 30728
rect 30791 30688 31116 30716
rect 30791 30685 30803 30688
rect 30745 30679 30803 30685
rect 31110 30676 31116 30688
rect 31168 30676 31174 30728
rect 31220 30725 31248 30756
rect 31294 30744 31300 30796
rect 31352 30784 31358 30796
rect 32306 30784 32312 30796
rect 31352 30756 31524 30784
rect 32267 30756 32312 30784
rect 31352 30744 31358 30756
rect 31496 30725 31524 30756
rect 32306 30744 32312 30756
rect 32364 30744 32370 30796
rect 31205 30719 31263 30725
rect 31205 30685 31217 30719
rect 31251 30685 31263 30719
rect 31205 30679 31263 30685
rect 31389 30719 31447 30725
rect 31389 30685 31401 30719
rect 31435 30685 31447 30719
rect 31389 30679 31447 30685
rect 31481 30719 31539 30725
rect 31481 30685 31493 30719
rect 31527 30685 31539 30719
rect 31481 30679 31539 30685
rect 22094 30648 22100 30660
rect 20548 30620 22100 30648
rect 22094 30608 22100 30620
rect 22152 30608 22158 30660
rect 30006 30608 30012 30660
rect 30064 30648 30070 30660
rect 30469 30651 30527 30657
rect 30469 30648 30481 30651
rect 30064 30620 30481 30648
rect 30064 30608 30070 30620
rect 30469 30617 30481 30620
rect 30515 30617 30527 30651
rect 30469 30611 30527 30617
rect 30561 30651 30619 30657
rect 30561 30617 30573 30651
rect 30607 30648 30619 30651
rect 30607 30620 31248 30648
rect 30607 30617 30619 30620
rect 30561 30611 30619 30617
rect 31220 30592 31248 30620
rect 17819 30552 18368 30580
rect 17819 30549 17831 30552
rect 17773 30543 17831 30549
rect 18598 30540 18604 30592
rect 18656 30580 18662 30592
rect 18693 30583 18751 30589
rect 18693 30580 18705 30583
rect 18656 30552 18705 30580
rect 18656 30540 18662 30552
rect 18693 30549 18705 30552
rect 18739 30549 18751 30583
rect 18693 30543 18751 30549
rect 22186 30540 22192 30592
rect 22244 30580 22250 30592
rect 22922 30580 22928 30592
rect 22244 30552 22928 30580
rect 22244 30540 22250 30552
rect 22922 30540 22928 30552
rect 22980 30580 22986 30592
rect 23109 30583 23167 30589
rect 23109 30580 23121 30583
rect 22980 30552 23121 30580
rect 22980 30540 22986 30552
rect 23109 30549 23121 30552
rect 23155 30549 23167 30583
rect 23658 30580 23664 30592
rect 23619 30552 23664 30580
rect 23109 30543 23167 30549
rect 23658 30540 23664 30552
rect 23716 30540 23722 30592
rect 24946 30540 24952 30592
rect 25004 30580 25010 30592
rect 26145 30583 26203 30589
rect 26145 30580 26157 30583
rect 25004 30552 26157 30580
rect 25004 30540 25010 30552
rect 26145 30549 26157 30552
rect 26191 30549 26203 30583
rect 30190 30580 30196 30592
rect 30151 30552 30196 30580
rect 26145 30543 26203 30549
rect 30190 30540 30196 30552
rect 30248 30540 30254 30592
rect 31202 30540 31208 30592
rect 31260 30540 31266 30592
rect 31404 30580 31432 30679
rect 31570 30676 31576 30728
rect 31628 30716 31634 30728
rect 31628 30688 31673 30716
rect 31628 30676 31634 30688
rect 34606 30676 34612 30728
rect 34664 30716 34670 30728
rect 35268 30725 35296 30892
rect 39301 30889 39313 30892
rect 39347 30889 39359 30923
rect 39301 30883 39359 30889
rect 35710 30744 35716 30796
rect 35768 30784 35774 30796
rect 37001 30787 37059 30793
rect 37001 30784 37013 30787
rect 35768 30756 37013 30784
rect 35768 30744 35774 30756
rect 35253 30719 35311 30725
rect 35253 30716 35265 30719
rect 34664 30688 35265 30716
rect 34664 30676 34670 30688
rect 35253 30685 35265 30688
rect 35299 30685 35311 30719
rect 35894 30716 35900 30728
rect 35855 30688 35900 30716
rect 35253 30679 35311 30685
rect 35894 30676 35900 30688
rect 35952 30676 35958 30728
rect 36280 30725 36308 30756
rect 37001 30753 37013 30756
rect 37047 30753 37059 30787
rect 37001 30747 37059 30753
rect 37550 30744 37556 30796
rect 37608 30784 37614 30796
rect 37921 30787 37979 30793
rect 37921 30784 37933 30787
rect 37608 30756 37933 30784
rect 37608 30744 37614 30756
rect 37921 30753 37933 30756
rect 37967 30753 37979 30787
rect 37921 30747 37979 30753
rect 36081 30716 36139 30722
rect 36081 30682 36093 30716
rect 36127 30682 36139 30716
rect 36081 30676 36139 30682
rect 36176 30716 36234 30722
rect 36176 30682 36188 30716
rect 36222 30682 36234 30716
rect 36176 30676 36234 30682
rect 36265 30719 36323 30725
rect 36265 30685 36277 30719
rect 36311 30685 36323 30719
rect 58158 30716 58164 30728
rect 58119 30688 58164 30716
rect 36265 30679 36323 30685
rect 58158 30676 58164 30688
rect 58216 30676 58222 30728
rect 31849 30651 31907 30657
rect 31849 30617 31861 30651
rect 31895 30648 31907 30651
rect 32554 30651 32612 30657
rect 32554 30648 32566 30651
rect 31895 30620 32566 30648
rect 31895 30617 31907 30620
rect 31849 30611 31907 30617
rect 32554 30617 32566 30620
rect 32600 30617 32612 30651
rect 32554 30611 32612 30617
rect 35069 30651 35127 30657
rect 35069 30617 35081 30651
rect 35115 30648 35127 30651
rect 35342 30648 35348 30660
rect 35115 30620 35348 30648
rect 35115 30617 35127 30620
rect 35069 30611 35127 30617
rect 35342 30608 35348 30620
rect 35400 30608 35406 30660
rect 35437 30651 35495 30657
rect 35437 30617 35449 30651
rect 35483 30648 35495 30651
rect 36096 30648 36124 30676
rect 36191 30648 36219 30676
rect 35483 30620 36124 30648
rect 36188 30620 36219 30648
rect 36541 30651 36599 30657
rect 35483 30617 35495 30620
rect 35437 30611 35495 30617
rect 36188 30592 36216 30620
rect 36541 30617 36553 30651
rect 36587 30648 36599 30651
rect 38166 30651 38224 30657
rect 38166 30648 38178 30651
rect 36587 30620 38178 30648
rect 36587 30617 36599 30620
rect 36541 30611 36599 30617
rect 38166 30617 38178 30620
rect 38212 30617 38224 30651
rect 38166 30611 38224 30617
rect 32306 30580 32312 30592
rect 31404 30552 32312 30580
rect 32306 30540 32312 30552
rect 32364 30540 32370 30592
rect 32398 30540 32404 30592
rect 32456 30580 32462 30592
rect 32950 30580 32956 30592
rect 32456 30552 32956 30580
rect 32456 30540 32462 30552
rect 32950 30540 32956 30552
rect 33008 30580 33014 30592
rect 33689 30583 33747 30589
rect 33689 30580 33701 30583
rect 33008 30552 33701 30580
rect 33008 30540 33014 30552
rect 33689 30549 33701 30552
rect 33735 30549 33747 30583
rect 33689 30543 33747 30549
rect 36170 30540 36176 30592
rect 36228 30540 36234 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 11793 30379 11851 30385
rect 11793 30345 11805 30379
rect 11839 30376 11851 30379
rect 11882 30376 11888 30388
rect 11839 30348 11888 30376
rect 11839 30345 11851 30348
rect 11793 30339 11851 30345
rect 11882 30336 11888 30348
rect 11940 30336 11946 30388
rect 14826 30336 14832 30388
rect 14884 30376 14890 30388
rect 14884 30348 16620 30376
rect 14884 30336 14890 30348
rect 4617 30311 4675 30317
rect 4617 30277 4629 30311
rect 4663 30308 4675 30311
rect 4890 30308 4896 30320
rect 4663 30280 4896 30308
rect 4663 30277 4675 30280
rect 4617 30271 4675 30277
rect 4890 30268 4896 30280
rect 4948 30268 4954 30320
rect 6362 30268 6368 30320
rect 6420 30308 6426 30320
rect 6822 30308 6828 30320
rect 6420 30280 6828 30308
rect 6420 30268 6426 30280
rect 6822 30268 6828 30280
rect 6880 30308 6886 30320
rect 15381 30311 15439 30317
rect 15381 30308 15393 30311
rect 6880 30280 7788 30308
rect 6880 30268 6886 30280
rect 2222 30200 2228 30252
rect 2280 30240 2286 30252
rect 2409 30243 2467 30249
rect 2409 30240 2421 30243
rect 2280 30212 2421 30240
rect 2280 30200 2286 30212
rect 2409 30209 2421 30212
rect 2455 30209 2467 30243
rect 2409 30203 2467 30209
rect 2498 30200 2504 30252
rect 2556 30240 2562 30252
rect 2665 30243 2723 30249
rect 2665 30240 2677 30243
rect 2556 30212 2677 30240
rect 2556 30200 2562 30212
rect 2665 30209 2677 30212
rect 2711 30209 2723 30243
rect 2665 30203 2723 30209
rect 4433 30243 4491 30249
rect 4433 30209 4445 30243
rect 4479 30240 4491 30243
rect 5258 30240 5264 30252
rect 4479 30212 5264 30240
rect 4479 30209 4491 30212
rect 4433 30203 4491 30209
rect 5258 30200 5264 30212
rect 5316 30200 5322 30252
rect 7489 30243 7547 30249
rect 7489 30209 7501 30243
rect 7535 30240 7547 30243
rect 7650 30240 7656 30252
rect 7535 30212 7656 30240
rect 7535 30209 7547 30212
rect 7489 30203 7547 30209
rect 7650 30200 7656 30212
rect 7708 30200 7714 30252
rect 7760 30249 7788 30280
rect 12406 30280 15393 30308
rect 12406 30252 12434 30280
rect 15381 30277 15393 30280
rect 15427 30277 15439 30311
rect 15381 30271 15439 30277
rect 15473 30311 15531 30317
rect 15473 30277 15485 30311
rect 15519 30308 15531 30311
rect 15746 30308 15752 30320
rect 15519 30280 15752 30308
rect 15519 30277 15531 30280
rect 15473 30271 15531 30277
rect 15746 30268 15752 30280
rect 15804 30308 15810 30320
rect 16206 30308 16212 30320
rect 15804 30280 16212 30308
rect 15804 30268 15810 30280
rect 16206 30268 16212 30280
rect 16264 30268 16270 30320
rect 7745 30243 7803 30249
rect 7745 30209 7757 30243
rect 7791 30209 7803 30243
rect 7745 30203 7803 30209
rect 11977 30243 12035 30249
rect 11977 30209 11989 30243
rect 12023 30240 12035 30243
rect 12342 30240 12348 30252
rect 12023 30212 12348 30240
rect 12023 30209 12035 30212
rect 11977 30203 12035 30209
rect 12342 30200 12348 30212
rect 12400 30212 12434 30252
rect 12400 30200 12406 30212
rect 13998 30200 14004 30252
rect 14056 30240 14062 30252
rect 15286 30249 15292 30252
rect 15105 30243 15163 30249
rect 15105 30240 15117 30243
rect 14056 30212 15117 30240
rect 14056 30200 14062 30212
rect 15105 30209 15117 30212
rect 15151 30209 15163 30243
rect 15105 30203 15163 30209
rect 15253 30243 15292 30249
rect 15253 30209 15265 30243
rect 15253 30203 15292 30209
rect 15286 30200 15292 30203
rect 15344 30200 15350 30252
rect 15570 30243 15628 30249
rect 15570 30240 15582 30243
rect 15396 30212 15582 30240
rect 9950 30132 9956 30184
rect 10008 30172 10014 30184
rect 12161 30175 12219 30181
rect 12161 30172 12173 30175
rect 10008 30144 12173 30172
rect 10008 30132 10014 30144
rect 12161 30141 12173 30144
rect 12207 30172 12219 30175
rect 15396 30172 15424 30212
rect 15570 30209 15582 30212
rect 15616 30240 15628 30243
rect 16482 30240 16488 30252
rect 15616 30212 16488 30240
rect 15616 30209 15628 30212
rect 15570 30203 15628 30209
rect 16482 30200 16488 30212
rect 16540 30200 16546 30252
rect 16592 30240 16620 30348
rect 16666 30336 16672 30388
rect 16724 30376 16730 30388
rect 17034 30376 17040 30388
rect 16724 30348 17040 30376
rect 16724 30336 16730 30348
rect 17034 30336 17040 30348
rect 17092 30376 17098 30388
rect 17221 30379 17279 30385
rect 17221 30376 17233 30379
rect 17092 30348 17233 30376
rect 17092 30336 17098 30348
rect 17221 30345 17233 30348
rect 17267 30376 17279 30379
rect 17267 30348 18460 30376
rect 17267 30345 17279 30348
rect 17221 30339 17279 30345
rect 18322 30308 18328 30320
rect 17696 30280 18328 30308
rect 17696 30249 17724 30280
rect 18322 30268 18328 30280
rect 18380 30268 18386 30320
rect 17954 30249 17960 30252
rect 17681 30243 17739 30249
rect 17681 30240 17693 30243
rect 16592 30212 17693 30240
rect 17681 30209 17693 30212
rect 17727 30209 17739 30243
rect 17681 30203 17739 30209
rect 17948 30203 17960 30249
rect 18012 30240 18018 30252
rect 18432 30240 18460 30348
rect 18506 30336 18512 30388
rect 18564 30376 18570 30388
rect 19061 30379 19119 30385
rect 19061 30376 19073 30379
rect 18564 30348 19073 30376
rect 18564 30336 18570 30348
rect 19061 30345 19073 30348
rect 19107 30376 19119 30379
rect 19150 30376 19156 30388
rect 19107 30348 19156 30376
rect 19107 30345 19119 30348
rect 19061 30339 19119 30345
rect 19150 30336 19156 30348
rect 19208 30336 19214 30388
rect 19426 30336 19432 30388
rect 19484 30376 19490 30388
rect 19521 30379 19579 30385
rect 19521 30376 19533 30379
rect 19484 30348 19533 30376
rect 19484 30336 19490 30348
rect 19521 30345 19533 30348
rect 19567 30345 19579 30379
rect 29454 30376 29460 30388
rect 19521 30339 19579 30345
rect 19628 30348 29460 30376
rect 19628 30240 19656 30348
rect 29454 30336 29460 30348
rect 29512 30376 29518 30388
rect 30834 30376 30840 30388
rect 29512 30348 30840 30376
rect 29512 30336 29518 30348
rect 30834 30336 30840 30348
rect 30892 30336 30898 30388
rect 31202 30336 31208 30388
rect 31260 30376 31266 30388
rect 31260 30348 33732 30376
rect 31260 30336 31266 30348
rect 20993 30311 21051 30317
rect 20993 30308 21005 30311
rect 20088 30280 21005 30308
rect 18012 30212 18048 30240
rect 18432 30212 19656 30240
rect 19797 30243 19855 30249
rect 17954 30200 17960 30203
rect 18012 30200 18018 30212
rect 19797 30209 19809 30243
rect 19843 30209 19855 30243
rect 19797 30203 19855 30209
rect 19902 30246 19960 30252
rect 19902 30212 19914 30246
rect 19948 30212 19960 30246
rect 19902 30206 19960 30212
rect 20002 30246 20060 30252
rect 20002 30212 20014 30246
rect 20048 30243 20060 30246
rect 20088 30243 20116 30280
rect 20993 30277 21005 30280
rect 21039 30277 21051 30311
rect 20993 30271 21051 30277
rect 21634 30268 21640 30320
rect 21692 30308 21698 30320
rect 22094 30308 22100 30320
rect 21692 30280 22100 30308
rect 21692 30268 21698 30280
rect 22094 30268 22100 30280
rect 22152 30268 22158 30320
rect 22465 30311 22523 30317
rect 22465 30277 22477 30311
rect 22511 30308 22523 30311
rect 24118 30308 24124 30320
rect 22511 30280 24124 30308
rect 22511 30277 22523 30280
rect 22465 30271 22523 30277
rect 24118 30268 24124 30280
rect 24176 30268 24182 30320
rect 24581 30311 24639 30317
rect 24581 30277 24593 30311
rect 24627 30308 24639 30311
rect 25130 30308 25136 30320
rect 24627 30280 25136 30308
rect 24627 30277 24639 30280
rect 24581 30271 24639 30277
rect 25130 30268 25136 30280
rect 25188 30268 25194 30320
rect 30650 30308 30656 30320
rect 28828 30280 30656 30308
rect 20048 30215 20116 30243
rect 20177 30243 20235 30249
rect 20048 30212 20060 30215
rect 20002 30206 20060 30212
rect 20177 30209 20189 30243
rect 20223 30240 20235 30243
rect 20346 30240 20352 30252
rect 20223 30212 20352 30240
rect 20223 30209 20235 30212
rect 12207 30144 12434 30172
rect 12207 30141 12219 30144
rect 12161 30135 12219 30141
rect 3786 30104 3792 30116
rect 3747 30076 3792 30104
rect 3786 30064 3792 30076
rect 3844 30064 3850 30116
rect 3510 29996 3516 30048
rect 3568 30036 3574 30048
rect 4249 30039 4307 30045
rect 4249 30036 4261 30039
rect 3568 30008 4261 30036
rect 3568 29996 3574 30008
rect 4249 30005 4261 30008
rect 4295 30005 4307 30039
rect 6362 30036 6368 30048
rect 6323 30008 6368 30036
rect 4249 29999 4307 30005
rect 6362 29996 6368 30008
rect 6420 29996 6426 30048
rect 10505 30039 10563 30045
rect 10505 30005 10517 30039
rect 10551 30036 10563 30039
rect 10778 30036 10784 30048
rect 10551 30008 10784 30036
rect 10551 30005 10563 30008
rect 10505 29999 10563 30005
rect 10778 29996 10784 30008
rect 10836 29996 10842 30048
rect 12406 30036 12434 30144
rect 14016 30144 15424 30172
rect 14016 30116 14044 30144
rect 19242 30132 19248 30184
rect 19300 30172 19306 30184
rect 19812 30172 19840 30203
rect 19300 30144 19840 30172
rect 19300 30132 19306 30144
rect 19917 30116 19945 30206
rect 20177 30203 20235 30209
rect 20346 30200 20352 30212
rect 20404 30200 20410 30252
rect 20438 30200 20444 30252
rect 20496 30240 20502 30252
rect 20625 30243 20683 30249
rect 20625 30240 20637 30243
rect 20496 30212 20637 30240
rect 20496 30200 20502 30212
rect 20625 30209 20637 30212
rect 20671 30209 20683 30243
rect 20625 30203 20683 30209
rect 20809 30243 20867 30249
rect 20809 30209 20821 30243
rect 20855 30240 20867 30243
rect 20898 30240 20904 30252
rect 20855 30212 20904 30240
rect 20855 30209 20867 30212
rect 20809 30203 20867 30209
rect 20898 30200 20904 30212
rect 20956 30240 20962 30252
rect 21818 30240 21824 30252
rect 20956 30212 21824 30240
rect 20956 30200 20962 30212
rect 21818 30200 21824 30212
rect 21876 30200 21882 30252
rect 22278 30200 22284 30252
rect 22336 30240 22342 30252
rect 22373 30243 22431 30249
rect 22373 30240 22385 30243
rect 22336 30212 22385 30240
rect 22336 30200 22342 30212
rect 22373 30209 22385 30212
rect 22419 30209 22431 30243
rect 22373 30203 22431 30209
rect 22557 30243 22615 30249
rect 22557 30209 22569 30243
rect 22603 30209 22615 30243
rect 22738 30240 22744 30252
rect 22699 30212 22744 30240
rect 22557 30203 22615 30209
rect 21634 30132 21640 30184
rect 21692 30172 21698 30184
rect 22572 30172 22600 30203
rect 22738 30200 22744 30212
rect 22796 30200 22802 30252
rect 24026 30200 24032 30252
rect 24084 30240 24090 30252
rect 24213 30243 24271 30249
rect 24213 30240 24225 30243
rect 24084 30212 24225 30240
rect 24084 30200 24090 30212
rect 24213 30209 24225 30212
rect 24259 30209 24271 30243
rect 24213 30203 24271 30209
rect 24397 30243 24455 30249
rect 24397 30209 24409 30243
rect 24443 30240 24455 30243
rect 24946 30240 24952 30252
rect 24443 30212 24952 30240
rect 24443 30209 24455 30212
rect 24397 30203 24455 30209
rect 24946 30200 24952 30212
rect 25004 30200 25010 30252
rect 25406 30249 25412 30252
rect 25402 30240 25412 30249
rect 25056 30212 25412 30240
rect 21692 30144 22600 30172
rect 21692 30132 21698 30144
rect 13998 30064 14004 30116
rect 14056 30064 14062 30116
rect 15838 30104 15844 30116
rect 14108 30076 15844 30104
rect 12713 30039 12771 30045
rect 12713 30036 12725 30039
rect 12406 30008 12725 30036
rect 12713 30005 12725 30008
rect 12759 30036 12771 30039
rect 14108 30036 14136 30076
rect 15838 30064 15844 30076
rect 15896 30064 15902 30116
rect 19886 30064 19892 30116
rect 19944 30064 19950 30116
rect 21450 30064 21456 30116
rect 21508 30104 21514 30116
rect 25056 30104 25084 30212
rect 25402 30203 25412 30212
rect 25406 30200 25412 30203
rect 25464 30200 25470 30252
rect 25498 30200 25504 30252
rect 25556 30240 25562 30252
rect 26145 30243 26203 30249
rect 26145 30240 26157 30243
rect 25556 30212 26157 30240
rect 25556 30200 25562 30212
rect 26145 30209 26157 30212
rect 26191 30209 26203 30243
rect 26145 30203 26203 30209
rect 27890 30200 27896 30252
rect 27948 30240 27954 30252
rect 28626 30240 28632 30252
rect 27948 30212 28632 30240
rect 27948 30200 27954 30212
rect 28626 30200 28632 30212
rect 28684 30240 28690 30252
rect 28828 30249 28856 30280
rect 30650 30268 30656 30280
rect 30708 30268 30714 30320
rect 32214 30308 32220 30320
rect 32175 30280 32220 30308
rect 32214 30268 32220 30280
rect 32272 30268 32278 30320
rect 32306 30268 32312 30320
rect 32364 30308 32370 30320
rect 32585 30311 32643 30317
rect 32585 30308 32597 30311
rect 32364 30280 32597 30308
rect 32364 30268 32370 30280
rect 32585 30277 32597 30280
rect 32631 30277 32643 30311
rect 33594 30308 33600 30320
rect 33555 30280 33600 30308
rect 32585 30271 32643 30277
rect 33594 30268 33600 30280
rect 33652 30268 33658 30320
rect 33704 30317 33732 30348
rect 34422 30336 34428 30388
rect 34480 30376 34486 30388
rect 35345 30379 35403 30385
rect 35345 30376 35357 30379
rect 34480 30348 35357 30376
rect 34480 30336 34486 30348
rect 35345 30345 35357 30348
rect 35391 30345 35403 30379
rect 37645 30379 37703 30385
rect 37645 30376 37657 30379
rect 35345 30339 35403 30345
rect 36004 30348 37657 30376
rect 33689 30311 33747 30317
rect 33689 30277 33701 30311
rect 33735 30308 33747 30311
rect 33962 30308 33968 30320
rect 33735 30280 33968 30308
rect 33735 30277 33747 30280
rect 33689 30271 33747 30277
rect 33962 30268 33968 30280
rect 34020 30268 34026 30320
rect 34606 30308 34612 30320
rect 34567 30280 34612 30308
rect 34606 30268 34612 30280
rect 34664 30268 34670 30320
rect 28721 30243 28779 30249
rect 28721 30240 28733 30243
rect 28684 30212 28733 30240
rect 28684 30200 28690 30212
rect 28721 30209 28733 30212
rect 28767 30209 28779 30243
rect 28721 30203 28779 30209
rect 28813 30243 28871 30249
rect 28813 30209 28825 30243
rect 28859 30209 28871 30243
rect 28813 30203 28871 30209
rect 28902 30200 28908 30252
rect 28960 30240 28966 30252
rect 29089 30243 29147 30249
rect 28960 30212 29005 30240
rect 28960 30200 28966 30212
rect 29089 30209 29101 30243
rect 29135 30240 29147 30243
rect 30282 30240 30288 30252
rect 29135 30212 30288 30240
rect 29135 30209 29147 30212
rect 29089 30203 29147 30209
rect 30282 30200 30288 30212
rect 30340 30200 30346 30252
rect 30469 30243 30527 30249
rect 30469 30209 30481 30243
rect 30515 30240 30527 30243
rect 30558 30240 30564 30252
rect 30515 30212 30564 30240
rect 30515 30209 30527 30212
rect 30469 30203 30527 30209
rect 30558 30200 30564 30212
rect 30616 30200 30622 30252
rect 32398 30240 32404 30252
rect 32359 30212 32404 30240
rect 32398 30200 32404 30212
rect 32456 30200 32462 30252
rect 33502 30200 33508 30252
rect 33560 30240 33566 30252
rect 33870 30240 33876 30252
rect 33560 30212 33605 30240
rect 33831 30212 33876 30240
rect 33560 30200 33566 30212
rect 33870 30200 33876 30212
rect 33928 30200 33934 30252
rect 34330 30200 34336 30252
rect 34388 30240 34394 30252
rect 34517 30243 34575 30249
rect 34517 30240 34529 30243
rect 34388 30212 34529 30240
rect 34388 30200 34394 30212
rect 34517 30209 34529 30212
rect 34563 30209 34575 30243
rect 34517 30203 34575 30209
rect 34701 30243 34759 30249
rect 34701 30209 34713 30243
rect 34747 30209 34759 30243
rect 34701 30203 34759 30209
rect 27430 30172 27436 30184
rect 25240 30144 27436 30172
rect 25240 30113 25268 30144
rect 27430 30132 27436 30144
rect 27488 30132 27494 30184
rect 30006 30132 30012 30184
rect 30064 30172 30070 30184
rect 30193 30175 30251 30181
rect 30193 30172 30205 30175
rect 30064 30144 30205 30172
rect 30064 30132 30070 30144
rect 30193 30141 30205 30144
rect 30239 30141 30251 30175
rect 30193 30135 30251 30141
rect 34054 30132 34060 30184
rect 34112 30172 34118 30184
rect 34716 30172 34744 30203
rect 34790 30200 34796 30252
rect 34848 30240 34854 30252
rect 34885 30243 34943 30249
rect 34885 30240 34897 30243
rect 34848 30212 34897 30240
rect 34848 30200 34854 30212
rect 34885 30209 34897 30212
rect 34931 30209 34943 30243
rect 34885 30203 34943 30209
rect 34112 30144 34744 30172
rect 34112 30132 34118 30144
rect 21508 30076 25084 30104
rect 25225 30107 25283 30113
rect 21508 30064 21514 30076
rect 25225 30073 25237 30107
rect 25271 30073 25283 30107
rect 25958 30104 25964 30116
rect 25919 30076 25964 30104
rect 25225 30067 25283 30073
rect 25958 30064 25964 30076
rect 26016 30064 26022 30116
rect 28258 30064 28264 30116
rect 28316 30104 28322 30116
rect 31481 30107 31539 30113
rect 31481 30104 31493 30107
rect 28316 30076 31493 30104
rect 28316 30064 28322 30076
rect 31481 30073 31493 30076
rect 31527 30104 31539 30107
rect 31570 30104 31576 30116
rect 31527 30076 31576 30104
rect 31527 30073 31539 30076
rect 31481 30067 31539 30073
rect 31570 30064 31576 30076
rect 31628 30104 31634 30116
rect 32214 30104 32220 30116
rect 31628 30076 32220 30104
rect 31628 30064 31634 30076
rect 32214 30064 32220 30076
rect 32272 30064 32278 30116
rect 12759 30008 14136 30036
rect 15749 30039 15807 30045
rect 12759 30005 12771 30008
rect 12713 29999 12771 30005
rect 15749 30005 15761 30039
rect 15795 30036 15807 30039
rect 16390 30036 16396 30048
rect 15795 30008 16396 30036
rect 15795 30005 15807 30008
rect 15749 29999 15807 30005
rect 16390 29996 16396 30008
rect 16448 29996 16454 30048
rect 22189 30039 22247 30045
rect 22189 30005 22201 30039
rect 22235 30036 22247 30039
rect 22370 30036 22376 30048
rect 22235 30008 22376 30036
rect 22235 30005 22247 30008
rect 22189 29999 22247 30005
rect 22370 29996 22376 30008
rect 22428 29996 22434 30048
rect 25498 29996 25504 30048
rect 25556 30036 25562 30048
rect 26973 30039 27031 30045
rect 26973 30036 26985 30039
rect 25556 30008 26985 30036
rect 25556 29996 25562 30008
rect 26973 30005 26985 30008
rect 27019 30005 27031 30039
rect 27890 30036 27896 30048
rect 27851 30008 27896 30036
rect 26973 29999 27031 30005
rect 27890 29996 27896 30008
rect 27948 29996 27954 30048
rect 28442 30036 28448 30048
rect 28403 30008 28448 30036
rect 28442 29996 28448 30008
rect 28500 29996 28506 30048
rect 33321 30039 33379 30045
rect 33321 30005 33333 30039
rect 33367 30036 33379 30039
rect 33594 30036 33600 30048
rect 33367 30008 33600 30036
rect 33367 30005 33379 30008
rect 33321 29999 33379 30005
rect 33594 29996 33600 30008
rect 33652 29996 33658 30048
rect 34330 30036 34336 30048
rect 34291 30008 34336 30036
rect 34330 29996 34336 30008
rect 34388 29996 34394 30048
rect 35360 30036 35388 30339
rect 35894 30240 35900 30252
rect 35855 30212 35900 30240
rect 35894 30200 35900 30212
rect 35952 30200 35958 30252
rect 36004 30246 36032 30348
rect 37645 30345 37657 30348
rect 37691 30345 37703 30379
rect 37645 30339 37703 30345
rect 37274 30308 37280 30320
rect 37235 30280 37280 30308
rect 37274 30268 37280 30280
rect 37332 30268 37338 30320
rect 36060 30249 36118 30255
rect 36060 30246 36072 30249
rect 36004 30218 36072 30246
rect 36060 30215 36072 30218
rect 36106 30215 36118 30249
rect 36060 30209 36118 30215
rect 36170 30200 36176 30252
rect 36228 30240 36234 30252
rect 36354 30249 36360 30252
rect 36311 30243 36360 30249
rect 36228 30212 36273 30240
rect 36228 30200 36234 30212
rect 36311 30209 36323 30243
rect 36357 30209 36360 30243
rect 36311 30203 36360 30209
rect 36354 30200 36360 30203
rect 36412 30200 36418 30252
rect 37458 30240 37464 30252
rect 37419 30212 37464 30240
rect 37458 30200 37464 30212
rect 37516 30200 37522 30252
rect 36354 30036 36360 30048
rect 35360 30008 36360 30036
rect 36354 29996 36360 30008
rect 36412 29996 36418 30048
rect 36541 30039 36599 30045
rect 36541 30005 36553 30039
rect 36587 30036 36599 30039
rect 39666 30036 39672 30048
rect 36587 30008 39672 30036
rect 36587 30005 36599 30008
rect 36541 29999 36599 30005
rect 39666 29996 39672 30008
rect 39724 29996 39730 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 2133 29835 2191 29841
rect 2133 29801 2145 29835
rect 2179 29832 2191 29835
rect 2498 29832 2504 29844
rect 2179 29804 2504 29832
rect 2179 29801 2191 29804
rect 2133 29795 2191 29801
rect 2498 29792 2504 29804
rect 2556 29792 2562 29844
rect 8938 29792 8944 29844
rect 8996 29832 9002 29844
rect 9125 29835 9183 29841
rect 9125 29832 9137 29835
rect 8996 29804 9137 29832
rect 8996 29792 9002 29804
rect 9125 29801 9137 29804
rect 9171 29801 9183 29835
rect 9125 29795 9183 29801
rect 11698 29792 11704 29844
rect 11756 29832 11762 29844
rect 11974 29832 11980 29844
rect 11756 29804 11980 29832
rect 11756 29792 11762 29804
rect 11974 29792 11980 29804
rect 12032 29792 12038 29844
rect 15470 29832 15476 29844
rect 15431 29804 15476 29832
rect 15470 29792 15476 29804
rect 15528 29792 15534 29844
rect 17954 29792 17960 29844
rect 18012 29832 18018 29844
rect 18049 29835 18107 29841
rect 18049 29832 18061 29835
rect 18012 29804 18061 29832
rect 18012 29792 18018 29804
rect 18049 29801 18061 29804
rect 18095 29801 18107 29835
rect 18049 29795 18107 29801
rect 19429 29835 19487 29841
rect 19429 29801 19441 29835
rect 19475 29832 19487 29835
rect 20346 29832 20352 29844
rect 19475 29804 20352 29832
rect 19475 29801 19487 29804
rect 19429 29795 19487 29801
rect 2590 29724 2596 29776
rect 2648 29764 2654 29776
rect 2648 29736 2728 29764
rect 2648 29724 2654 29736
rect 2314 29588 2320 29640
rect 2372 29637 2378 29640
rect 2372 29631 2421 29637
rect 2372 29597 2375 29631
rect 2409 29597 2421 29631
rect 2372 29591 2421 29597
rect 2482 29628 2540 29634
rect 2482 29594 2494 29628
rect 2528 29594 2540 29628
rect 2372 29588 2378 29591
rect 2482 29588 2540 29594
rect 2593 29631 2651 29637
rect 2593 29597 2605 29631
rect 2639 29628 2651 29631
rect 2700 29628 2728 29736
rect 14182 29724 14188 29776
rect 14240 29764 14246 29776
rect 16945 29767 17003 29773
rect 16945 29764 16957 29767
rect 14240 29736 16957 29764
rect 14240 29724 14246 29736
rect 16945 29733 16957 29736
rect 16991 29733 17003 29767
rect 16945 29727 17003 29733
rect 4706 29696 4712 29708
rect 4448 29668 4712 29696
rect 2639 29600 2728 29628
rect 2639 29597 2651 29600
rect 2593 29591 2651 29597
rect 2774 29588 2780 29640
rect 2832 29628 2838 29640
rect 3418 29628 3424 29640
rect 2832 29600 3424 29628
rect 2832 29588 2838 29600
rect 3418 29588 3424 29600
rect 3476 29588 3482 29640
rect 3602 29588 3608 29640
rect 3660 29628 3666 29640
rect 4448 29637 4476 29668
rect 4706 29656 4712 29668
rect 4764 29656 4770 29708
rect 9493 29699 9551 29705
rect 9493 29665 9505 29699
rect 9539 29696 9551 29699
rect 9950 29696 9956 29708
rect 9539 29668 9956 29696
rect 9539 29665 9551 29668
rect 9493 29659 9551 29665
rect 9950 29656 9956 29668
rect 10008 29656 10014 29708
rect 16960 29640 16988 29727
rect 4157 29631 4215 29637
rect 4157 29628 4169 29631
rect 3660 29600 4169 29628
rect 3660 29588 3666 29600
rect 4157 29597 4169 29600
rect 4203 29597 4215 29631
rect 4157 29591 4215 29597
rect 4433 29631 4491 29637
rect 4433 29597 4445 29631
rect 4479 29597 4491 29631
rect 4433 29591 4491 29597
rect 4525 29631 4583 29637
rect 4525 29597 4537 29631
rect 4571 29628 4583 29631
rect 5626 29628 5632 29640
rect 4571 29600 5632 29628
rect 4571 29597 4583 29600
rect 4525 29591 4583 29597
rect 5626 29588 5632 29600
rect 5684 29588 5690 29640
rect 9306 29628 9312 29640
rect 9267 29600 9312 29628
rect 9306 29588 9312 29600
rect 9364 29588 9370 29640
rect 10597 29631 10655 29637
rect 10597 29597 10609 29631
rect 10643 29628 10655 29631
rect 12158 29628 12164 29640
rect 10643 29600 12164 29628
rect 10643 29597 10655 29600
rect 10597 29591 10655 29597
rect 12158 29588 12164 29600
rect 12216 29588 12222 29640
rect 13170 29588 13176 29640
rect 13228 29628 13234 29640
rect 14918 29628 14924 29640
rect 13228 29600 14924 29628
rect 13228 29588 13234 29600
rect 14918 29588 14924 29600
rect 14976 29628 14982 29640
rect 15105 29631 15163 29637
rect 15105 29628 15117 29631
rect 14976 29600 15117 29628
rect 14976 29588 14982 29600
rect 15105 29597 15117 29600
rect 15151 29597 15163 29631
rect 15105 29591 15163 29597
rect 15289 29631 15347 29637
rect 15289 29597 15301 29631
rect 15335 29628 15347 29631
rect 15746 29628 15752 29640
rect 15335 29600 15752 29628
rect 15335 29597 15347 29600
rect 15289 29591 15347 29597
rect 15746 29588 15752 29600
rect 15804 29588 15810 29640
rect 16942 29628 16948 29640
rect 16855 29600 16948 29628
rect 16942 29588 16948 29600
rect 17000 29628 17006 29640
rect 18325 29631 18383 29637
rect 18325 29628 18337 29631
rect 17000 29600 18337 29628
rect 17000 29588 17006 29600
rect 18325 29597 18337 29600
rect 18371 29597 18383 29631
rect 18325 29591 18383 29597
rect 18417 29631 18475 29637
rect 18417 29597 18429 29631
rect 18463 29597 18475 29631
rect 18417 29591 18475 29597
rect 18509 29631 18567 29637
rect 18509 29597 18521 29631
rect 18555 29628 18567 29631
rect 18598 29628 18604 29640
rect 18555 29600 18604 29628
rect 18555 29597 18567 29600
rect 18509 29591 18567 29597
rect 2497 29560 2525 29588
rect 3234 29560 3240 29572
rect 2497 29532 3240 29560
rect 3234 29520 3240 29532
rect 3292 29520 3298 29572
rect 4338 29560 4344 29572
rect 4299 29532 4344 29560
rect 4338 29520 4344 29532
rect 4396 29520 4402 29572
rect 7742 29520 7748 29572
rect 7800 29560 7806 29572
rect 10686 29560 10692 29572
rect 7800 29532 10692 29560
rect 7800 29520 7806 29532
rect 10686 29520 10692 29532
rect 10744 29520 10750 29572
rect 10864 29563 10922 29569
rect 10864 29529 10876 29563
rect 10910 29560 10922 29563
rect 10962 29560 10968 29572
rect 10910 29532 10968 29560
rect 10910 29529 10922 29532
rect 10864 29523 10922 29529
rect 10962 29520 10968 29532
rect 11020 29520 11026 29572
rect 12618 29520 12624 29572
rect 12676 29560 12682 29572
rect 17497 29563 17555 29569
rect 17497 29560 17509 29563
rect 12676 29532 17509 29560
rect 12676 29520 12682 29532
rect 17497 29529 17509 29532
rect 17543 29560 17555 29563
rect 18432 29560 18460 29591
rect 18598 29588 18604 29600
rect 18656 29588 18662 29640
rect 18693 29631 18751 29637
rect 18693 29597 18705 29631
rect 18739 29628 18751 29631
rect 18874 29628 18880 29640
rect 18739 29600 18880 29628
rect 18739 29597 18751 29600
rect 18693 29591 18751 29597
rect 18874 29588 18880 29600
rect 18932 29628 18938 29640
rect 19444 29628 19472 29795
rect 20346 29792 20352 29804
rect 20404 29832 20410 29844
rect 20717 29835 20775 29841
rect 20717 29832 20729 29835
rect 20404 29804 20729 29832
rect 20404 29792 20410 29804
rect 20717 29801 20729 29804
rect 20763 29801 20775 29835
rect 21542 29832 21548 29844
rect 21503 29804 21548 29832
rect 20717 29795 20775 29801
rect 21542 29792 21548 29804
rect 21600 29792 21606 29844
rect 23290 29792 23296 29844
rect 23348 29832 23354 29844
rect 23845 29835 23903 29841
rect 23845 29832 23857 29835
rect 23348 29804 23857 29832
rect 23348 29792 23354 29804
rect 23845 29801 23857 29804
rect 23891 29832 23903 29835
rect 23891 29804 25084 29832
rect 23891 29801 23903 29804
rect 23845 29795 23903 29801
rect 20165 29767 20223 29773
rect 20165 29733 20177 29767
rect 20211 29764 20223 29767
rect 20806 29764 20812 29776
rect 20211 29736 20812 29764
rect 20211 29733 20223 29736
rect 20165 29727 20223 29733
rect 20806 29724 20812 29736
rect 20864 29724 20870 29776
rect 24854 29764 24860 29776
rect 24504 29736 24860 29764
rect 18932 29600 19472 29628
rect 20809 29631 20867 29637
rect 18932 29588 18938 29600
rect 20809 29597 20821 29631
rect 20855 29628 20867 29631
rect 21174 29628 21180 29640
rect 20855 29600 21180 29628
rect 20855 29597 20867 29600
rect 20809 29591 20867 29597
rect 18782 29560 18788 29572
rect 17543 29532 18788 29560
rect 17543 29529 17555 29532
rect 17497 29523 17555 29529
rect 18782 29520 18788 29532
rect 18840 29560 18846 29572
rect 19426 29560 19432 29572
rect 18840 29532 19432 29560
rect 18840 29520 18846 29532
rect 19426 29520 19432 29532
rect 19484 29560 19490 29572
rect 19886 29560 19892 29572
rect 19484 29532 19892 29560
rect 19484 29520 19490 29532
rect 19886 29520 19892 29532
rect 19944 29560 19950 29572
rect 19981 29563 20039 29569
rect 19981 29560 19993 29563
rect 19944 29532 19993 29560
rect 19944 29520 19950 29532
rect 19981 29529 19993 29532
rect 20027 29529 20039 29563
rect 19981 29523 20039 29529
rect 20346 29520 20352 29572
rect 20404 29560 20410 29572
rect 20824 29560 20852 29591
rect 21174 29588 21180 29600
rect 21232 29588 21238 29640
rect 21361 29631 21419 29637
rect 21361 29597 21373 29631
rect 21407 29628 21419 29631
rect 21450 29628 21456 29640
rect 21407 29600 21456 29628
rect 21407 29597 21419 29600
rect 21361 29591 21419 29597
rect 21450 29588 21456 29600
rect 21508 29588 21514 29640
rect 22186 29628 22192 29640
rect 22147 29600 22192 29628
rect 22186 29588 22192 29600
rect 22244 29588 22250 29640
rect 22278 29588 22284 29640
rect 22336 29628 22342 29640
rect 22557 29631 22615 29637
rect 22557 29628 22569 29631
rect 22336 29600 22569 29628
rect 22336 29588 22342 29600
rect 22557 29597 22569 29600
rect 22603 29597 22615 29631
rect 22557 29591 22615 29597
rect 20404 29532 20852 29560
rect 20404 29520 20410 29532
rect 21634 29520 21640 29572
rect 21692 29560 21698 29572
rect 22373 29563 22431 29569
rect 22373 29560 22385 29563
rect 21692 29532 22385 29560
rect 21692 29520 21698 29532
rect 22373 29529 22385 29532
rect 22419 29529 22431 29563
rect 22373 29523 22431 29529
rect 22465 29563 22523 29569
rect 22465 29529 22477 29563
rect 22511 29560 22523 29563
rect 24504 29560 24532 29736
rect 24854 29724 24860 29736
rect 24912 29724 24918 29776
rect 24670 29628 24676 29640
rect 24631 29600 24676 29628
rect 24670 29588 24676 29600
rect 24728 29588 24734 29640
rect 24854 29628 24860 29640
rect 24815 29600 24860 29628
rect 24854 29588 24860 29600
rect 24912 29588 24918 29640
rect 25056 29637 25084 29804
rect 25406 29792 25412 29844
rect 25464 29832 25470 29844
rect 28350 29832 28356 29844
rect 25464 29804 28356 29832
rect 25464 29792 25470 29804
rect 28350 29792 28356 29804
rect 28408 29792 28414 29844
rect 28902 29792 28908 29844
rect 28960 29832 28966 29844
rect 28997 29835 29055 29841
rect 28997 29832 29009 29835
rect 28960 29804 29009 29832
rect 28960 29792 28966 29804
rect 28997 29801 29009 29804
rect 29043 29801 29055 29835
rect 28997 29795 29055 29801
rect 30653 29835 30711 29841
rect 30653 29801 30665 29835
rect 30699 29832 30711 29835
rect 31294 29832 31300 29844
rect 30699 29804 31300 29832
rect 30699 29801 30711 29804
rect 30653 29795 30711 29801
rect 31294 29792 31300 29804
rect 31352 29792 31358 29844
rect 34238 29792 34244 29844
rect 34296 29832 34302 29844
rect 34885 29835 34943 29841
rect 34296 29804 34836 29832
rect 34296 29792 34302 29804
rect 33134 29724 33140 29776
rect 33192 29764 33198 29776
rect 33192 29736 34744 29764
rect 33192 29724 33198 29736
rect 27157 29699 27215 29705
rect 27157 29665 27169 29699
rect 27203 29696 27215 29699
rect 27522 29696 27528 29708
rect 27203 29668 27528 29696
rect 27203 29665 27215 29668
rect 27157 29659 27215 29665
rect 27522 29656 27528 29668
rect 27580 29656 27586 29708
rect 29086 29696 29092 29708
rect 28828 29668 29092 29696
rect 24949 29631 25007 29637
rect 24949 29597 24961 29631
rect 24995 29597 25007 29631
rect 24949 29591 25007 29597
rect 25041 29631 25099 29637
rect 25041 29597 25053 29631
rect 25087 29628 25099 29631
rect 28258 29628 28264 29640
rect 25087 29600 28264 29628
rect 25087 29597 25099 29600
rect 25041 29591 25099 29597
rect 22511 29532 24532 29560
rect 24964 29560 24992 29591
rect 28258 29588 28264 29600
rect 28316 29588 28322 29640
rect 28534 29588 28540 29640
rect 28592 29628 28598 29640
rect 28828 29637 28856 29668
rect 29086 29656 29092 29668
rect 29144 29696 29150 29708
rect 29144 29668 30144 29696
rect 29144 29656 29150 29668
rect 28629 29631 28687 29637
rect 28629 29628 28641 29631
rect 28592 29600 28641 29628
rect 28592 29588 28598 29600
rect 28629 29597 28641 29600
rect 28675 29597 28687 29631
rect 28629 29591 28687 29597
rect 28813 29631 28871 29637
rect 28813 29597 28825 29631
rect 28859 29597 28871 29631
rect 29730 29628 29736 29640
rect 29691 29600 29736 29628
rect 28813 29591 28871 29597
rect 29730 29588 29736 29600
rect 29788 29588 29794 29640
rect 29822 29588 29828 29640
rect 29880 29628 29886 29640
rect 30116 29637 30144 29668
rect 30101 29631 30159 29637
rect 29880 29600 29925 29628
rect 29880 29588 29886 29600
rect 30101 29597 30113 29631
rect 30147 29597 30159 29631
rect 30101 29591 30159 29597
rect 30561 29631 30619 29637
rect 30561 29597 30573 29631
rect 30607 29597 30619 29631
rect 30742 29628 30748 29640
rect 30703 29600 30748 29628
rect 30561 29591 30619 29597
rect 25222 29560 25228 29572
rect 24964 29532 25228 29560
rect 22511 29529 22523 29532
rect 22465 29523 22523 29529
rect 25056 29504 25084 29532
rect 25222 29520 25228 29532
rect 25280 29520 25286 29572
rect 25317 29563 25375 29569
rect 25317 29529 25329 29563
rect 25363 29560 25375 29563
rect 26890 29563 26948 29569
rect 26890 29560 26902 29563
rect 25363 29532 26902 29560
rect 25363 29529 25375 29532
rect 25317 29523 25375 29529
rect 26890 29529 26902 29532
rect 26936 29529 26948 29563
rect 29914 29560 29920 29572
rect 29875 29532 29920 29560
rect 26890 29523 26948 29529
rect 29914 29520 29920 29532
rect 29972 29560 29978 29572
rect 30374 29560 30380 29572
rect 29972 29532 30380 29560
rect 29972 29520 29978 29532
rect 30374 29520 30380 29532
rect 30432 29560 30438 29572
rect 30576 29560 30604 29591
rect 30742 29588 30748 29600
rect 30800 29628 30806 29640
rect 31205 29631 31263 29637
rect 31205 29628 31217 29631
rect 30800 29600 31217 29628
rect 30800 29588 30806 29600
rect 31205 29597 31217 29600
rect 31251 29597 31263 29631
rect 31205 29591 31263 29597
rect 33502 29588 33508 29640
rect 33560 29628 33566 29640
rect 33781 29631 33839 29637
rect 33781 29628 33793 29631
rect 33560 29600 33793 29628
rect 33560 29588 33566 29600
rect 33781 29597 33793 29600
rect 33827 29597 33839 29631
rect 33962 29628 33968 29640
rect 33923 29600 33968 29628
rect 33781 29591 33839 29597
rect 33962 29588 33968 29600
rect 34020 29588 34026 29640
rect 34149 29631 34207 29637
rect 34149 29597 34161 29631
rect 34195 29628 34207 29631
rect 34514 29628 34520 29640
rect 34195 29600 34520 29628
rect 34195 29597 34207 29600
rect 34149 29591 34207 29597
rect 34514 29588 34520 29600
rect 34572 29588 34578 29640
rect 34716 29637 34744 29736
rect 34808 29696 34836 29804
rect 34885 29801 34897 29835
rect 34931 29832 34943 29835
rect 35342 29832 35348 29844
rect 34931 29804 35348 29832
rect 34931 29801 34943 29804
rect 34885 29795 34943 29801
rect 35342 29792 35348 29804
rect 35400 29792 35406 29844
rect 35434 29724 35440 29776
rect 35492 29764 35498 29776
rect 37921 29767 37979 29773
rect 37921 29764 37933 29767
rect 35492 29736 37933 29764
rect 35492 29724 35498 29736
rect 37921 29733 37933 29736
rect 37967 29733 37979 29767
rect 37921 29727 37979 29733
rect 35345 29699 35403 29705
rect 35345 29696 35357 29699
rect 34808 29668 35357 29696
rect 35345 29665 35357 29668
rect 35391 29665 35403 29699
rect 35345 29659 35403 29665
rect 35621 29699 35679 29705
rect 35621 29665 35633 29699
rect 35667 29696 35679 29699
rect 36170 29696 36176 29708
rect 35667 29668 36176 29696
rect 35667 29665 35679 29668
rect 35621 29659 35679 29665
rect 36170 29656 36176 29668
rect 36228 29656 36234 29708
rect 34701 29631 34759 29637
rect 34701 29597 34713 29631
rect 34747 29597 34759 29631
rect 37458 29628 37464 29640
rect 34701 29591 34759 29597
rect 36648 29600 37464 29628
rect 30432 29532 30604 29560
rect 33873 29563 33931 29569
rect 30432 29520 30438 29532
rect 33873 29529 33885 29563
rect 33919 29560 33931 29563
rect 36648 29560 36676 29600
rect 37458 29588 37464 29600
rect 37516 29588 37522 29640
rect 39298 29628 39304 29640
rect 39259 29600 39304 29628
rect 39298 29588 39304 29600
rect 39356 29588 39362 29640
rect 58158 29628 58164 29640
rect 58119 29600 58164 29628
rect 58158 29588 58164 29600
rect 58216 29588 58222 29640
rect 33919 29532 36676 29560
rect 33919 29529 33931 29532
rect 33873 29523 33931 29529
rect 36722 29520 36728 29572
rect 36780 29560 36786 29572
rect 39034 29563 39092 29569
rect 39034 29560 39046 29563
rect 36780 29532 39046 29560
rect 36780 29520 36786 29532
rect 39034 29529 39046 29532
rect 39080 29529 39092 29563
rect 39034 29523 39092 29529
rect 4709 29495 4767 29501
rect 4709 29461 4721 29495
rect 4755 29492 4767 29495
rect 4890 29492 4896 29504
rect 4755 29464 4896 29492
rect 4755 29461 4767 29464
rect 4709 29455 4767 29461
rect 4890 29452 4896 29464
rect 4948 29452 4954 29504
rect 6914 29452 6920 29504
rect 6972 29492 6978 29504
rect 7193 29495 7251 29501
rect 7193 29492 7205 29495
rect 6972 29464 7205 29492
rect 6972 29452 6978 29464
rect 7193 29461 7205 29464
rect 7239 29492 7251 29495
rect 8018 29492 8024 29504
rect 7239 29464 8024 29492
rect 7239 29461 7251 29464
rect 7193 29455 7251 29461
rect 8018 29452 8024 29464
rect 8076 29452 8082 29504
rect 14182 29492 14188 29504
rect 14143 29464 14188 29492
rect 14182 29452 14188 29464
rect 14240 29452 14246 29504
rect 22741 29495 22799 29501
rect 22741 29461 22753 29495
rect 22787 29492 22799 29495
rect 22922 29492 22928 29504
rect 22787 29464 22928 29492
rect 22787 29461 22799 29464
rect 22741 29455 22799 29461
rect 22922 29452 22928 29464
rect 22980 29452 22986 29504
rect 25038 29452 25044 29504
rect 25096 29452 25102 29504
rect 25774 29492 25780 29504
rect 25735 29464 25780 29492
rect 25774 29452 25780 29464
rect 25832 29452 25838 29504
rect 29546 29492 29552 29504
rect 29507 29464 29552 29492
rect 29546 29452 29552 29464
rect 29604 29452 29610 29504
rect 33410 29452 33416 29504
rect 33468 29492 33474 29504
rect 33597 29495 33655 29501
rect 33597 29492 33609 29495
rect 33468 29464 33609 29492
rect 33468 29452 33474 29464
rect 33597 29461 33609 29464
rect 33643 29461 33655 29495
rect 33597 29455 33655 29461
rect 34146 29452 34152 29504
rect 34204 29492 34210 29504
rect 36630 29492 36636 29504
rect 34204 29464 36636 29492
rect 34204 29452 34210 29464
rect 36630 29452 36636 29464
rect 36688 29452 36694 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 9306 29288 9312 29300
rect 5368 29260 9312 29288
rect 3510 29220 3516 29232
rect 3344 29192 3516 29220
rect 2958 29112 2964 29164
rect 3016 29161 3022 29164
rect 3016 29155 3065 29161
rect 3016 29121 3019 29155
rect 3053 29121 3065 29155
rect 3142 29152 3148 29164
rect 3103 29124 3148 29152
rect 3016 29115 3065 29121
rect 3016 29112 3022 29115
rect 3142 29112 3148 29124
rect 3200 29112 3206 29164
rect 3258 29161 3316 29167
rect 3258 29127 3270 29161
rect 3304 29158 3316 29161
rect 3344 29158 3372 29192
rect 3510 29180 3516 29192
rect 3568 29180 3574 29232
rect 4338 29180 4344 29232
rect 4396 29220 4402 29232
rect 4433 29223 4491 29229
rect 4433 29220 4445 29223
rect 4396 29192 4445 29220
rect 4396 29180 4402 29192
rect 4433 29189 4445 29192
rect 4479 29220 4491 29223
rect 5368 29220 5396 29260
rect 9306 29248 9312 29260
rect 9364 29248 9370 29300
rect 10962 29288 10968 29300
rect 9416 29260 10824 29288
rect 10923 29260 10968 29288
rect 5534 29220 5540 29232
rect 4479 29192 5396 29220
rect 5495 29192 5540 29220
rect 4479 29189 4491 29192
rect 4433 29183 4491 29189
rect 3304 29130 3372 29158
rect 3304 29127 3316 29130
rect 3258 29121 3316 29127
rect 3418 29112 3424 29164
rect 3476 29152 3482 29164
rect 3476 29124 3521 29152
rect 3476 29112 3482 29124
rect 3786 29112 3792 29164
rect 3844 29152 3850 29164
rect 4249 29155 4307 29161
rect 4249 29152 4261 29155
rect 3844 29124 4261 29152
rect 3844 29112 3850 29124
rect 4249 29121 4261 29124
rect 4295 29121 4307 29155
rect 4249 29115 4307 29121
rect 4525 29155 4583 29161
rect 4525 29121 4537 29155
rect 4571 29121 4583 29155
rect 4525 29115 4583 29121
rect 4617 29155 4675 29161
rect 4617 29121 4629 29155
rect 4663 29121 4675 29155
rect 5258 29152 5264 29164
rect 5219 29124 5264 29152
rect 4617 29115 4675 29121
rect 1946 29044 1952 29096
rect 2004 29084 2010 29096
rect 4540 29084 4568 29115
rect 2004 29056 2774 29084
rect 2004 29044 2010 29056
rect 2746 29016 2774 29056
rect 3804 29056 4568 29084
rect 4632 29084 4660 29115
rect 5258 29112 5264 29124
rect 5316 29112 5322 29164
rect 5368 29152 5396 29192
rect 5534 29180 5540 29192
rect 5592 29180 5598 29232
rect 8386 29180 8392 29232
rect 8444 29220 8450 29232
rect 9416 29220 9444 29260
rect 8444 29192 9444 29220
rect 8444 29180 8450 29192
rect 9674 29180 9680 29232
rect 9732 29220 9738 29232
rect 10796 29220 10824 29260
rect 10962 29248 10968 29260
rect 11020 29248 11026 29300
rect 18782 29288 18788 29300
rect 18695 29260 18788 29288
rect 18782 29248 18788 29260
rect 18840 29288 18846 29300
rect 19242 29288 19248 29300
rect 18840 29260 19248 29288
rect 18840 29248 18846 29260
rect 19242 29248 19248 29260
rect 19300 29248 19306 29300
rect 20438 29288 20444 29300
rect 20399 29260 20444 29288
rect 20438 29248 20444 29260
rect 20496 29248 20502 29300
rect 21269 29291 21327 29297
rect 21269 29257 21281 29291
rect 21315 29288 21327 29291
rect 21450 29288 21456 29300
rect 21315 29260 21456 29288
rect 21315 29257 21327 29260
rect 21269 29251 21327 29257
rect 21450 29248 21456 29260
rect 21508 29248 21514 29300
rect 24397 29291 24455 29297
rect 24397 29257 24409 29291
rect 24443 29288 24455 29291
rect 24854 29288 24860 29300
rect 24443 29260 24860 29288
rect 24443 29257 24455 29260
rect 24397 29251 24455 29257
rect 24854 29248 24860 29260
rect 24912 29248 24918 29300
rect 24949 29291 25007 29297
rect 24949 29257 24961 29291
rect 24995 29288 25007 29291
rect 26050 29288 26056 29300
rect 24995 29260 26056 29288
rect 24995 29257 25007 29260
rect 24949 29251 25007 29257
rect 26050 29248 26056 29260
rect 26108 29288 26114 29300
rect 26108 29260 27568 29288
rect 26108 29248 26114 29260
rect 13262 29220 13268 29232
rect 9732 29192 10640 29220
rect 10796 29192 13268 29220
rect 9732 29180 9738 29192
rect 5445 29155 5503 29161
rect 5445 29152 5457 29155
rect 5368 29124 5457 29152
rect 5445 29121 5457 29124
rect 5491 29121 5503 29155
rect 5626 29152 5632 29164
rect 5587 29124 5632 29152
rect 5445 29115 5503 29121
rect 5626 29112 5632 29124
rect 5684 29112 5690 29164
rect 6822 29112 6828 29164
rect 6880 29152 6886 29164
rect 7837 29155 7895 29161
rect 7837 29152 7849 29155
rect 6880 29124 7849 29152
rect 6880 29112 6886 29124
rect 7837 29121 7849 29124
rect 7883 29121 7895 29155
rect 7837 29115 7895 29121
rect 8104 29155 8162 29161
rect 8104 29121 8116 29155
rect 8150 29152 8162 29155
rect 9030 29152 9036 29164
rect 8150 29124 9036 29152
rect 8150 29121 8162 29124
rect 8104 29115 8162 29121
rect 9030 29112 9036 29124
rect 9088 29112 9094 29164
rect 9858 29112 9864 29164
rect 9916 29152 9922 29164
rect 10327 29155 10385 29161
rect 10500 29158 10558 29164
rect 10612 29161 10640 29192
rect 13262 29180 13268 29192
rect 13320 29220 13326 29232
rect 14918 29220 14924 29232
rect 13320 29192 13584 29220
rect 14879 29192 14924 29220
rect 13320 29180 13326 29192
rect 10244 29152 10339 29155
rect 9916 29127 10339 29152
rect 9916 29124 10272 29127
rect 9916 29112 9922 29124
rect 10327 29121 10339 29127
rect 10373 29121 10385 29155
rect 10327 29115 10385 29121
rect 10428 29130 10512 29158
rect 5644 29084 5672 29112
rect 10428 29096 10456 29130
rect 10500 29124 10512 29130
rect 10546 29124 10558 29158
rect 10500 29118 10558 29124
rect 10597 29155 10655 29161
rect 10597 29121 10609 29155
rect 10643 29121 10655 29155
rect 10597 29115 10655 29121
rect 10689 29155 10747 29161
rect 10689 29121 10701 29155
rect 10735 29127 10824 29155
rect 13446 29152 13452 29164
rect 10735 29121 10747 29127
rect 10689 29115 10747 29121
rect 4632 29056 5672 29084
rect 2746 28988 3648 29016
rect 2774 28908 2780 28960
rect 2832 28948 2838 28960
rect 3620 28948 3648 28988
rect 3804 28948 3832 29056
rect 10410 29044 10416 29096
rect 10468 29044 10474 29096
rect 4801 29019 4859 29025
rect 4801 28985 4813 29019
rect 4847 29016 4859 29019
rect 4982 29016 4988 29028
rect 4847 28988 4988 29016
rect 4847 28985 4859 28988
rect 4801 28979 4859 28985
rect 4982 28976 4988 28988
rect 5040 28976 5046 29028
rect 10796 29016 10824 29127
rect 13407 29124 13452 29152
rect 13446 29112 13452 29124
rect 13504 29112 13510 29164
rect 13556 29161 13584 29192
rect 14918 29180 14924 29192
rect 14976 29180 14982 29232
rect 15378 29180 15384 29232
rect 15436 29220 15442 29232
rect 23290 29220 23296 29232
rect 15436 29192 23296 29220
rect 15436 29180 15442 29192
rect 23290 29180 23296 29192
rect 23348 29180 23354 29232
rect 23382 29180 23388 29232
rect 23440 29220 23446 29232
rect 24213 29223 24271 29229
rect 24213 29220 24225 29223
rect 23440 29192 24225 29220
rect 23440 29180 23446 29192
rect 24213 29189 24225 29192
rect 24259 29220 24271 29223
rect 25774 29220 25780 29232
rect 24259 29192 25780 29220
rect 24259 29189 24271 29192
rect 24213 29183 24271 29189
rect 25774 29180 25780 29192
rect 25832 29180 25838 29232
rect 27540 29220 27568 29260
rect 28994 29248 29000 29300
rect 29052 29288 29058 29300
rect 29917 29291 29975 29297
rect 29917 29288 29929 29291
rect 29052 29260 29929 29288
rect 29052 29248 29058 29260
rect 29917 29257 29929 29260
rect 29963 29288 29975 29291
rect 30098 29288 30104 29300
rect 29963 29260 30104 29288
rect 29963 29257 29975 29260
rect 29917 29251 29975 29257
rect 30098 29248 30104 29260
rect 30156 29248 30162 29300
rect 31205 29291 31263 29297
rect 31205 29257 31217 29291
rect 31251 29288 31263 29291
rect 33134 29288 33140 29300
rect 31251 29260 33140 29288
rect 31251 29257 31263 29260
rect 31205 29251 31263 29257
rect 33134 29248 33140 29260
rect 33192 29248 33198 29300
rect 36722 29288 36728 29300
rect 36683 29260 36728 29288
rect 36722 29248 36728 29260
rect 36780 29248 36786 29300
rect 37458 29248 37464 29300
rect 37516 29288 37522 29300
rect 38565 29291 38623 29297
rect 38565 29288 38577 29291
rect 37516 29260 38577 29288
rect 37516 29248 37522 29260
rect 38565 29257 38577 29260
rect 38611 29257 38623 29291
rect 38565 29251 38623 29257
rect 34422 29220 34428 29232
rect 27540 29192 34428 29220
rect 34422 29180 34428 29192
rect 34480 29180 34486 29232
rect 35434 29220 35440 29232
rect 35395 29192 35440 29220
rect 35434 29180 35440 29192
rect 35492 29180 35498 29232
rect 35621 29223 35679 29229
rect 35621 29189 35633 29223
rect 35667 29220 35679 29223
rect 35667 29192 36308 29220
rect 35667 29189 35679 29192
rect 35621 29183 35679 29189
rect 13541 29155 13599 29161
rect 13541 29121 13553 29155
rect 13587 29121 13599 29155
rect 13541 29115 13599 29121
rect 13633 29155 13691 29161
rect 13633 29121 13645 29155
rect 13679 29121 13691 29155
rect 13633 29115 13691 29121
rect 13648 29084 13676 29115
rect 13722 29112 13728 29164
rect 13780 29152 13786 29164
rect 13817 29155 13875 29161
rect 13817 29152 13829 29155
rect 13780 29124 13829 29152
rect 13780 29112 13786 29124
rect 13817 29121 13829 29124
rect 13863 29121 13875 29155
rect 15102 29152 15108 29164
rect 15063 29124 15108 29152
rect 13817 29115 13875 29121
rect 15102 29112 15108 29124
rect 15160 29112 15166 29164
rect 19150 29112 19156 29164
rect 19208 29152 19214 29164
rect 19245 29155 19303 29161
rect 19245 29152 19257 29155
rect 19208 29124 19257 29152
rect 19208 29112 19214 29124
rect 19245 29121 19257 29124
rect 19291 29121 19303 29155
rect 19245 29115 19303 29121
rect 19334 29112 19340 29164
rect 19392 29152 19398 29164
rect 19429 29155 19487 29161
rect 19429 29152 19441 29155
rect 19392 29124 19441 29152
rect 19392 29112 19398 29124
rect 19429 29121 19441 29124
rect 19475 29121 19487 29155
rect 19429 29115 19487 29121
rect 19521 29155 19579 29161
rect 19521 29121 19533 29155
rect 19567 29121 19579 29155
rect 19521 29115 19579 29121
rect 19613 29155 19671 29161
rect 19613 29121 19625 29155
rect 19659 29152 19671 29155
rect 20070 29152 20076 29164
rect 19659 29124 20076 29152
rect 19659 29121 19671 29124
rect 19613 29115 19671 29121
rect 14458 29084 14464 29096
rect 13648 29056 14464 29084
rect 14458 29044 14464 29056
rect 14516 29044 14522 29096
rect 19536 29084 19564 29115
rect 20070 29112 20076 29124
rect 20128 29112 20134 29164
rect 21634 29112 21640 29164
rect 21692 29152 21698 29164
rect 22557 29155 22615 29161
rect 22557 29152 22569 29155
rect 21692 29124 22569 29152
rect 21692 29112 21698 29124
rect 22557 29121 22569 29124
rect 22603 29121 22615 29155
rect 24026 29152 24032 29164
rect 23987 29124 24032 29152
rect 22557 29115 22615 29121
rect 24026 29112 24032 29124
rect 24084 29112 24090 29164
rect 25133 29155 25191 29161
rect 25133 29121 25145 29155
rect 25179 29121 25191 29155
rect 25133 29115 25191 29121
rect 24946 29084 24952 29096
rect 19536 29056 24952 29084
rect 24946 29044 24952 29056
rect 25004 29044 25010 29096
rect 25148 29084 25176 29115
rect 25498 29112 25504 29164
rect 25556 29152 25562 29164
rect 25869 29155 25927 29161
rect 25869 29152 25881 29155
rect 25556 29124 25881 29152
rect 25556 29112 25562 29124
rect 25869 29121 25881 29124
rect 25915 29121 25927 29155
rect 28629 29155 28687 29161
rect 28629 29152 28641 29155
rect 25869 29115 25927 29121
rect 28092 29124 28641 29152
rect 25148 29056 26464 29084
rect 13170 29016 13176 29028
rect 10428 28988 10824 29016
rect 13131 28988 13176 29016
rect 10428 28960 10456 28988
rect 13170 28976 13176 28988
rect 13228 28976 13234 29028
rect 13446 28976 13452 29028
rect 13504 29016 13510 29028
rect 14182 29016 14188 29028
rect 13504 28988 14188 29016
rect 13504 28976 13510 28988
rect 14182 28976 14188 28988
rect 14240 29016 14246 29028
rect 14369 29019 14427 29025
rect 14369 29016 14381 29019
rect 14240 28988 14381 29016
rect 14240 28976 14246 28988
rect 14369 28985 14381 28988
rect 14415 29016 14427 29019
rect 15378 29016 15384 29028
rect 14415 28988 15384 29016
rect 14415 28985 14427 28988
rect 14369 28979 14427 28985
rect 15378 28976 15384 28988
rect 15436 28976 15442 29028
rect 18233 29019 18291 29025
rect 18233 28985 18245 29019
rect 18279 29016 18291 29019
rect 18874 29016 18880 29028
rect 18279 28988 18880 29016
rect 18279 28985 18291 28988
rect 18233 28979 18291 28985
rect 18874 28976 18880 28988
rect 18932 28976 18938 29028
rect 19797 29019 19855 29025
rect 19797 28985 19809 29019
rect 19843 29016 19855 29019
rect 20346 29016 20352 29028
rect 19843 28988 20352 29016
rect 19843 28985 19855 28988
rect 19797 28979 19855 28985
rect 20346 28976 20352 28988
rect 20404 28976 20410 29028
rect 22554 28976 22560 29028
rect 22612 29016 22618 29028
rect 22741 29019 22799 29025
rect 22741 29016 22753 29019
rect 22612 28988 22753 29016
rect 22612 28976 22618 28988
rect 22741 28985 22753 28988
rect 22787 29016 22799 29019
rect 22830 29016 22836 29028
rect 22787 28988 22836 29016
rect 22787 28985 22799 28988
rect 22741 28979 22799 28985
rect 22830 28976 22836 28988
rect 22888 28976 22894 29028
rect 25682 29016 25688 29028
rect 25643 28988 25688 29016
rect 25682 28976 25688 28988
rect 25740 28976 25746 29028
rect 26436 28960 26464 29056
rect 27614 28976 27620 29028
rect 27672 29016 27678 29028
rect 28092 29025 28120 29124
rect 28629 29121 28641 29124
rect 28675 29121 28687 29155
rect 28629 29115 28687 29121
rect 29730 29112 29736 29164
rect 29788 29152 29794 29164
rect 31021 29155 31079 29161
rect 31021 29152 31033 29155
rect 29788 29124 31033 29152
rect 29788 29112 29794 29124
rect 31021 29121 31033 29124
rect 31067 29121 31079 29155
rect 33502 29152 33508 29164
rect 33463 29124 33508 29152
rect 31021 29115 31079 29121
rect 33502 29112 33508 29124
rect 33560 29112 33566 29164
rect 35253 29155 35311 29161
rect 35253 29121 35265 29155
rect 35299 29152 35311 29155
rect 35342 29152 35348 29164
rect 35299 29124 35348 29152
rect 35299 29121 35311 29124
rect 35253 29115 35311 29121
rect 35342 29112 35348 29124
rect 35400 29112 35406 29164
rect 36078 29112 36084 29164
rect 36136 29152 36142 29164
rect 36280 29161 36308 29192
rect 39666 29180 39672 29232
rect 39724 29229 39730 29232
rect 39724 29220 39736 29229
rect 39724 29192 39769 29220
rect 39724 29183 39736 29192
rect 39724 29180 39730 29183
rect 36265 29155 36323 29161
rect 36136 29124 36181 29152
rect 36136 29112 36142 29124
rect 36265 29121 36277 29155
rect 36311 29121 36323 29155
rect 36265 29115 36323 29121
rect 36357 29155 36415 29161
rect 36357 29121 36369 29155
rect 36403 29121 36415 29155
rect 36357 29115 36415 29121
rect 36495 29155 36553 29161
rect 36495 29121 36507 29155
rect 36541 29152 36553 29155
rect 36630 29152 36636 29164
rect 36541 29124 36636 29152
rect 36541 29121 36553 29124
rect 36495 29115 36553 29121
rect 30834 29084 30840 29096
rect 30795 29056 30840 29084
rect 30834 29044 30840 29056
rect 30892 29044 30898 29096
rect 33781 29087 33839 29093
rect 33781 29053 33793 29087
rect 33827 29084 33839 29087
rect 34146 29084 34152 29096
rect 33827 29056 34152 29084
rect 33827 29053 33839 29056
rect 33781 29047 33839 29053
rect 34146 29044 34152 29056
rect 34204 29044 34210 29096
rect 36170 29044 36176 29096
rect 36228 29084 36234 29096
rect 36372 29084 36400 29115
rect 36630 29112 36636 29124
rect 36688 29112 36694 29164
rect 36228 29056 36400 29084
rect 39945 29087 40003 29093
rect 36228 29044 36234 29056
rect 39945 29053 39957 29087
rect 39991 29053 40003 29087
rect 39945 29047 40003 29053
rect 28077 29019 28135 29025
rect 28077 29016 28089 29019
rect 27672 28988 28089 29016
rect 27672 28976 27678 28988
rect 28077 28985 28089 28988
rect 28123 28985 28135 29019
rect 28077 28979 28135 28985
rect 30282 28976 30288 29028
rect 30340 29016 30346 29028
rect 31754 29016 31760 29028
rect 30340 28988 31760 29016
rect 30340 28976 30346 28988
rect 31754 28976 31760 28988
rect 31812 28976 31818 29028
rect 2832 28920 2877 28948
rect 3620 28920 3832 28948
rect 5813 28951 5871 28957
rect 2832 28908 2838 28920
rect 5813 28917 5825 28951
rect 5859 28948 5871 28951
rect 6638 28948 6644 28960
rect 5859 28920 6644 28948
rect 5859 28917 5871 28920
rect 5813 28911 5871 28917
rect 6638 28908 6644 28920
rect 6696 28908 6702 28960
rect 9214 28948 9220 28960
rect 9175 28920 9220 28948
rect 9214 28908 9220 28920
rect 9272 28908 9278 28960
rect 9861 28951 9919 28957
rect 9861 28917 9873 28951
rect 9907 28948 9919 28951
rect 10410 28948 10416 28960
rect 9907 28920 10416 28948
rect 9907 28917 9919 28920
rect 9861 28911 9919 28917
rect 10410 28908 10416 28920
rect 10468 28908 10474 28960
rect 15286 28948 15292 28960
rect 15247 28920 15292 28948
rect 15286 28908 15292 28920
rect 15344 28908 15350 28960
rect 16025 28951 16083 28957
rect 16025 28917 16037 28951
rect 16071 28948 16083 28951
rect 16206 28948 16212 28960
rect 16071 28920 16212 28948
rect 16071 28917 16083 28920
rect 16025 28911 16083 28917
rect 16206 28908 16212 28920
rect 16264 28908 16270 28960
rect 19334 28908 19340 28960
rect 19392 28948 19398 28960
rect 21634 28948 21640 28960
rect 19392 28920 21640 28948
rect 19392 28908 19398 28920
rect 21634 28908 21640 28920
rect 21692 28908 21698 28960
rect 26418 28948 26424 28960
rect 26379 28920 26424 28948
rect 26418 28908 26424 28920
rect 26476 28908 26482 28960
rect 38746 28908 38752 28960
rect 38804 28948 38810 28960
rect 39298 28948 39304 28960
rect 38804 28920 39304 28948
rect 38804 28908 38810 28920
rect 39298 28908 39304 28920
rect 39356 28948 39362 28960
rect 39960 28948 39988 29047
rect 39356 28920 39988 28948
rect 39356 28908 39362 28920
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 2314 28704 2320 28756
rect 2372 28744 2378 28756
rect 2866 28744 2872 28756
rect 2372 28716 2872 28744
rect 2372 28704 2378 28716
rect 2866 28704 2872 28716
rect 2924 28704 2930 28756
rect 9030 28744 9036 28756
rect 8991 28716 9036 28744
rect 9030 28704 9036 28716
rect 9088 28704 9094 28756
rect 13541 28747 13599 28753
rect 13541 28713 13553 28747
rect 13587 28744 13599 28747
rect 13722 28744 13728 28756
rect 13587 28716 13728 28744
rect 13587 28713 13599 28716
rect 13541 28707 13599 28713
rect 13722 28704 13728 28716
rect 13780 28704 13786 28756
rect 14458 28744 14464 28756
rect 14419 28716 14464 28744
rect 14458 28704 14464 28716
rect 14516 28704 14522 28756
rect 15654 28744 15660 28756
rect 14936 28716 15660 28744
rect 5626 28636 5632 28688
rect 5684 28676 5690 28688
rect 11698 28676 11704 28688
rect 5684 28648 11704 28676
rect 5684 28636 5690 28648
rect 8128 28549 8156 28648
rect 11698 28636 11704 28648
rect 11756 28636 11762 28688
rect 8386 28608 8392 28620
rect 8347 28580 8392 28608
rect 8386 28568 8392 28580
rect 8444 28568 8450 28620
rect 9582 28568 9588 28620
rect 9640 28608 9646 28620
rect 9640 28580 12480 28608
rect 9640 28568 9646 28580
rect 8113 28543 8171 28549
rect 8113 28509 8125 28543
rect 8159 28509 8171 28543
rect 8294 28540 8300 28552
rect 8255 28512 8300 28540
rect 8113 28503 8171 28509
rect 8294 28500 8300 28512
rect 8352 28500 8358 28552
rect 9263 28543 9321 28549
rect 9263 28509 9275 28543
rect 9309 28509 9321 28543
rect 9398 28540 9404 28552
rect 9359 28512 9404 28540
rect 9263 28503 9321 28509
rect 7561 28475 7619 28481
rect 7561 28441 7573 28475
rect 7607 28472 7619 28475
rect 8312 28472 8340 28500
rect 7607 28444 8340 28472
rect 7607 28441 7619 28444
rect 7561 28435 7619 28441
rect 2958 28364 2964 28416
rect 3016 28404 3022 28416
rect 3881 28407 3939 28413
rect 3881 28404 3893 28407
rect 3016 28376 3893 28404
rect 3016 28364 3022 28376
rect 3881 28373 3893 28376
rect 3927 28404 3939 28407
rect 4614 28404 4620 28416
rect 3927 28376 4620 28404
rect 3927 28373 3939 28376
rect 3881 28367 3939 28373
rect 4614 28364 4620 28376
rect 4672 28364 4678 28416
rect 9278 28404 9306 28503
rect 9398 28500 9404 28512
rect 9456 28500 9462 28552
rect 9490 28500 9496 28552
rect 9548 28540 9554 28552
rect 9677 28543 9735 28549
rect 9548 28512 9593 28540
rect 9548 28500 9554 28512
rect 9677 28509 9689 28543
rect 9723 28540 9735 28543
rect 10778 28540 10784 28552
rect 9723 28512 10784 28540
rect 9723 28509 9735 28512
rect 9677 28503 9735 28509
rect 10778 28500 10784 28512
rect 10836 28500 10842 28552
rect 12452 28549 12480 28580
rect 14936 28552 14964 28716
rect 15654 28704 15660 28716
rect 15712 28704 15718 28756
rect 19426 28704 19432 28756
rect 19484 28744 19490 28756
rect 19705 28747 19763 28753
rect 19705 28744 19717 28747
rect 19484 28716 19717 28744
rect 19484 28704 19490 28716
rect 19705 28713 19717 28716
rect 19751 28713 19763 28747
rect 20438 28744 20444 28756
rect 20399 28716 20444 28744
rect 19705 28707 19763 28713
rect 20438 28704 20444 28716
rect 20496 28704 20502 28756
rect 24762 28744 24768 28756
rect 24723 28716 24768 28744
rect 24762 28704 24768 28716
rect 24820 28704 24826 28756
rect 26970 28744 26976 28756
rect 26931 28716 26976 28744
rect 26970 28704 26976 28716
rect 27028 28704 27034 28756
rect 28997 28747 29055 28753
rect 28997 28713 29009 28747
rect 29043 28744 29055 28747
rect 29086 28744 29092 28756
rect 29043 28716 29092 28744
rect 29043 28713 29055 28716
rect 28997 28707 29055 28713
rect 29086 28704 29092 28716
rect 29144 28704 29150 28756
rect 30834 28704 30840 28756
rect 30892 28744 30898 28756
rect 31389 28747 31447 28753
rect 31389 28744 31401 28747
rect 30892 28716 31401 28744
rect 30892 28704 30898 28716
rect 31389 28713 31401 28716
rect 31435 28713 31447 28747
rect 31389 28707 31447 28713
rect 15286 28636 15292 28688
rect 15344 28636 15350 28688
rect 36170 28636 36176 28688
rect 36228 28636 36234 28688
rect 15304 28608 15332 28636
rect 30374 28608 30380 28620
rect 15120 28580 15332 28608
rect 30335 28580 30380 28608
rect 12437 28543 12495 28549
rect 12437 28509 12449 28543
rect 12483 28509 12495 28543
rect 12437 28503 12495 28509
rect 12526 28500 12532 28552
rect 12584 28540 12590 28552
rect 12621 28543 12679 28549
rect 12621 28540 12633 28543
rect 12584 28512 12633 28540
rect 12584 28500 12590 28512
rect 12621 28509 12633 28512
rect 12667 28509 12679 28543
rect 12802 28540 12808 28552
rect 12763 28512 12808 28540
rect 12621 28503 12679 28509
rect 12802 28500 12808 28512
rect 12860 28500 12866 28552
rect 14277 28543 14335 28549
rect 14277 28540 14289 28543
rect 13556 28512 14289 28540
rect 10229 28407 10287 28413
rect 10229 28404 10241 28407
rect 9278 28376 10241 28404
rect 10229 28373 10241 28376
rect 10275 28404 10287 28407
rect 10410 28404 10416 28416
rect 10275 28376 10416 28404
rect 10275 28373 10287 28376
rect 10229 28367 10287 28373
rect 10410 28364 10416 28376
rect 10468 28364 10474 28416
rect 10796 28413 10824 28500
rect 13556 28484 13584 28512
rect 14277 28509 14289 28512
rect 14323 28509 14335 28543
rect 14918 28540 14924 28552
rect 14879 28512 14924 28540
rect 14277 28503 14335 28509
rect 14918 28500 14924 28512
rect 14976 28500 14982 28552
rect 15120 28549 15148 28580
rect 30374 28568 30380 28580
rect 30432 28568 30438 28620
rect 33505 28611 33563 28617
rect 33505 28577 33517 28611
rect 33551 28608 33563 28611
rect 33962 28608 33968 28620
rect 33551 28580 33968 28608
rect 33551 28577 33563 28580
rect 33505 28571 33563 28577
rect 33962 28568 33968 28580
rect 34020 28568 34026 28620
rect 35434 28608 35440 28620
rect 34992 28580 35440 28608
rect 15105 28543 15163 28549
rect 15105 28509 15117 28543
rect 15151 28509 15163 28543
rect 15105 28503 15163 28509
rect 15197 28543 15255 28549
rect 15197 28509 15209 28543
rect 15243 28509 15255 28543
rect 15197 28503 15255 28509
rect 15289 28543 15347 28549
rect 15289 28509 15301 28543
rect 15335 28540 15347 28543
rect 15378 28540 15384 28552
rect 15335 28512 15384 28540
rect 15335 28509 15347 28512
rect 15289 28503 15347 28509
rect 12713 28475 12771 28481
rect 12713 28441 12725 28475
rect 12759 28472 12771 28475
rect 13538 28472 13544 28484
rect 12759 28444 13544 28472
rect 12759 28441 12771 28444
rect 12713 28435 12771 28441
rect 13538 28432 13544 28444
rect 13596 28432 13602 28484
rect 14093 28475 14151 28481
rect 14093 28441 14105 28475
rect 14139 28441 14151 28475
rect 15212 28472 15240 28503
rect 15378 28500 15384 28512
rect 15436 28500 15442 28552
rect 15562 28500 15568 28552
rect 15620 28500 15626 28552
rect 21450 28500 21456 28552
rect 21508 28540 21514 28552
rect 21634 28540 21640 28552
rect 21508 28512 21553 28540
rect 21595 28512 21640 28540
rect 21508 28500 21514 28512
rect 21634 28500 21640 28512
rect 21692 28500 21698 28552
rect 21818 28500 21824 28552
rect 21876 28540 21882 28552
rect 24949 28543 25007 28549
rect 21876 28512 21921 28540
rect 21876 28500 21882 28512
rect 24949 28509 24961 28543
rect 24995 28509 25007 28543
rect 26418 28540 26424 28552
rect 26331 28512 26424 28540
rect 24949 28503 25007 28509
rect 15580 28472 15608 28500
rect 16206 28472 16212 28484
rect 15212 28444 15608 28472
rect 16167 28444 16212 28472
rect 14093 28435 14151 28441
rect 10781 28407 10839 28413
rect 10781 28373 10793 28407
rect 10827 28404 10839 28407
rect 11514 28404 11520 28416
rect 10827 28376 11520 28404
rect 10827 28373 10839 28376
rect 10781 28367 10839 28373
rect 11514 28364 11520 28376
rect 11572 28364 11578 28416
rect 12986 28404 12992 28416
rect 12947 28376 12992 28404
rect 12986 28364 12992 28376
rect 13044 28364 13050 28416
rect 13078 28364 13084 28416
rect 13136 28404 13142 28416
rect 14108 28404 14136 28435
rect 16206 28432 16212 28444
rect 16264 28432 16270 28484
rect 16393 28475 16451 28481
rect 16393 28441 16405 28475
rect 16439 28472 16451 28475
rect 18230 28472 18236 28484
rect 16439 28444 18236 28472
rect 16439 28441 16451 28444
rect 16393 28435 16451 28441
rect 18230 28432 18236 28444
rect 18288 28472 18294 28484
rect 18414 28472 18420 28484
rect 18288 28444 18420 28472
rect 18288 28432 18294 28444
rect 18414 28432 18420 28444
rect 18472 28432 18478 28484
rect 21545 28475 21603 28481
rect 21545 28472 21557 28475
rect 21468 28444 21557 28472
rect 15562 28404 15568 28416
rect 13136 28376 14136 28404
rect 15523 28376 15568 28404
rect 13136 28364 13142 28376
rect 15562 28364 15568 28376
rect 15620 28364 15626 28416
rect 20990 28364 20996 28416
rect 21048 28404 21054 28416
rect 21269 28407 21327 28413
rect 21269 28404 21281 28407
rect 21048 28376 21281 28404
rect 21048 28364 21054 28376
rect 21269 28373 21281 28376
rect 21315 28373 21327 28407
rect 21468 28404 21496 28444
rect 21545 28441 21557 28444
rect 21591 28441 21603 28475
rect 21545 28435 21603 28441
rect 23566 28432 23572 28484
rect 23624 28472 23630 28484
rect 23845 28475 23903 28481
rect 23845 28472 23857 28475
rect 23624 28444 23857 28472
rect 23624 28432 23630 28444
rect 23845 28441 23857 28444
rect 23891 28472 23903 28475
rect 24964 28472 24992 28503
rect 26418 28500 26424 28512
rect 26476 28540 26482 28552
rect 27154 28540 27160 28552
rect 26476 28512 27160 28540
rect 26476 28500 26482 28512
rect 27154 28500 27160 28512
rect 27212 28500 27218 28552
rect 27614 28540 27620 28552
rect 27575 28512 27620 28540
rect 27614 28500 27620 28512
rect 27672 28500 27678 28552
rect 27884 28543 27942 28549
rect 27884 28509 27896 28543
rect 27930 28540 27942 28543
rect 28442 28540 28448 28552
rect 27930 28512 28448 28540
rect 27930 28509 27942 28512
rect 27884 28503 27942 28509
rect 28442 28500 28448 28512
rect 28500 28500 28506 28552
rect 30101 28543 30159 28549
rect 30101 28540 30113 28543
rect 29564 28512 30113 28540
rect 27062 28472 27068 28484
rect 23891 28444 27068 28472
rect 23891 28441 23903 28444
rect 23845 28435 23903 28441
rect 27062 28432 27068 28444
rect 27120 28432 27126 28484
rect 23382 28404 23388 28416
rect 21468 28376 23388 28404
rect 21269 28367 21327 28373
rect 23382 28364 23388 28376
rect 23440 28364 23446 28416
rect 25498 28404 25504 28416
rect 25459 28376 25504 28404
rect 25498 28364 25504 28376
rect 25556 28364 25562 28416
rect 26694 28364 26700 28416
rect 26752 28404 26758 28416
rect 29564 28413 29592 28512
rect 30101 28509 30113 28512
rect 30147 28540 30159 28543
rect 31570 28540 31576 28552
rect 30147 28512 31576 28540
rect 30147 28509 30159 28512
rect 30101 28503 30159 28509
rect 31570 28500 31576 28512
rect 31628 28500 31634 28552
rect 33781 28543 33839 28549
rect 33781 28509 33793 28543
rect 33827 28509 33839 28543
rect 33781 28503 33839 28509
rect 33796 28472 33824 28503
rect 34146 28500 34152 28552
rect 34204 28540 34210 28552
rect 34992 28549 35020 28580
rect 35434 28568 35440 28580
rect 35492 28568 35498 28620
rect 36188 28608 36216 28636
rect 36188 28580 36492 28608
rect 34885 28543 34943 28549
rect 34885 28540 34897 28543
rect 34204 28512 34897 28540
rect 34204 28500 34210 28512
rect 34885 28509 34897 28512
rect 34931 28509 34943 28543
rect 34885 28503 34943 28509
rect 34977 28543 35035 28549
rect 34977 28509 34989 28543
rect 35023 28509 35035 28543
rect 34977 28503 35035 28509
rect 35253 28543 35311 28549
rect 35253 28509 35265 28543
rect 35299 28540 35311 28543
rect 35526 28540 35532 28552
rect 35299 28512 35532 28540
rect 35299 28509 35311 28512
rect 35253 28503 35311 28509
rect 35526 28500 35532 28512
rect 35584 28500 35590 28552
rect 36078 28500 36084 28552
rect 36136 28540 36142 28552
rect 36173 28543 36231 28549
rect 36173 28540 36185 28543
rect 36136 28512 36185 28540
rect 36136 28500 36142 28512
rect 36173 28509 36185 28512
rect 36219 28509 36231 28543
rect 36354 28540 36360 28552
rect 36315 28512 36360 28540
rect 36173 28503 36231 28509
rect 36354 28500 36360 28512
rect 36412 28500 36418 28552
rect 36464 28549 36492 28580
rect 36449 28543 36507 28549
rect 36449 28509 36461 28543
rect 36495 28509 36507 28543
rect 36449 28503 36507 28509
rect 36541 28543 36599 28549
rect 36541 28509 36553 28543
rect 36587 28509 36599 28543
rect 38746 28540 38752 28552
rect 38707 28512 38752 28540
rect 36541 28503 36599 28509
rect 34422 28472 34428 28484
rect 33796 28444 34428 28472
rect 34422 28432 34428 28444
rect 34480 28472 34486 28484
rect 35069 28475 35127 28481
rect 35069 28472 35081 28475
rect 34480 28444 35081 28472
rect 34480 28432 34486 28444
rect 35069 28441 35081 28444
rect 35115 28441 35127 28475
rect 35069 28435 35127 28441
rect 35986 28432 35992 28484
rect 36044 28472 36050 28484
rect 36556 28472 36584 28503
rect 38746 28500 38752 28512
rect 38804 28500 38810 28552
rect 36044 28444 36584 28472
rect 36817 28475 36875 28481
rect 36044 28432 36050 28444
rect 36817 28441 36829 28475
rect 36863 28472 36875 28475
rect 38482 28475 38540 28481
rect 38482 28472 38494 28475
rect 36863 28444 38494 28472
rect 36863 28441 36875 28444
rect 36817 28435 36875 28441
rect 38482 28441 38494 28444
rect 38528 28441 38540 28475
rect 38482 28435 38540 28441
rect 29549 28407 29607 28413
rect 29549 28404 29561 28407
rect 26752 28376 29561 28404
rect 26752 28364 26758 28376
rect 29549 28373 29561 28376
rect 29595 28373 29607 28407
rect 29549 28367 29607 28373
rect 34606 28364 34612 28416
rect 34664 28404 34670 28416
rect 34701 28407 34759 28413
rect 34701 28404 34713 28407
rect 34664 28376 34713 28404
rect 34664 28364 34670 28376
rect 34701 28373 34713 28376
rect 34747 28373 34759 28407
rect 34701 28367 34759 28373
rect 36170 28364 36176 28416
rect 36228 28404 36234 28416
rect 37369 28407 37427 28413
rect 37369 28404 37381 28407
rect 36228 28376 37381 28404
rect 36228 28364 36234 28376
rect 37369 28373 37381 28376
rect 37415 28373 37427 28407
rect 37369 28367 37427 28373
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 3881 28203 3939 28209
rect 3881 28169 3893 28203
rect 3927 28200 3939 28203
rect 5258 28200 5264 28212
rect 3927 28172 5264 28200
rect 3927 28169 3939 28172
rect 3881 28163 3939 28169
rect 5258 28160 5264 28172
rect 5316 28160 5322 28212
rect 8478 28200 8484 28212
rect 8439 28172 8484 28200
rect 8478 28160 8484 28172
rect 8536 28160 8542 28212
rect 9309 28203 9367 28209
rect 9309 28169 9321 28203
rect 9355 28200 9367 28203
rect 9490 28200 9496 28212
rect 9355 28172 9496 28200
rect 9355 28169 9367 28172
rect 9309 28163 9367 28169
rect 9490 28160 9496 28172
rect 9548 28160 9554 28212
rect 11517 28203 11575 28209
rect 11517 28169 11529 28203
rect 11563 28200 11575 28203
rect 13078 28200 13084 28212
rect 11563 28172 13084 28200
rect 11563 28169 11575 28172
rect 11517 28163 11575 28169
rect 13078 28160 13084 28172
rect 13136 28160 13142 28212
rect 14737 28203 14795 28209
rect 14737 28200 14749 28203
rect 13924 28172 14749 28200
rect 2774 28141 2780 28144
rect 2768 28095 2780 28141
rect 2832 28132 2838 28144
rect 2832 28104 2868 28132
rect 2774 28092 2780 28095
rect 2832 28092 2838 28104
rect 6362 28092 6368 28144
rect 6420 28132 6426 28144
rect 7009 28135 7067 28141
rect 7009 28132 7021 28135
rect 6420 28104 7021 28132
rect 6420 28092 6426 28104
rect 7009 28101 7021 28104
rect 7055 28101 7067 28135
rect 7009 28095 7067 28101
rect 7837 28135 7895 28141
rect 7837 28101 7849 28135
rect 7883 28132 7895 28135
rect 8938 28132 8944 28144
rect 7883 28104 8524 28132
rect 8899 28104 8944 28132
rect 7883 28101 7895 28104
rect 7837 28095 7895 28101
rect 6638 28064 6644 28076
rect 6599 28036 6644 28064
rect 6638 28024 6644 28036
rect 6696 28024 6702 28076
rect 6730 28024 6736 28076
rect 6788 28064 6794 28076
rect 6914 28064 6920 28076
rect 6788 28036 6833 28064
rect 6875 28036 6920 28064
rect 6788 28024 6794 28036
rect 6914 28024 6920 28036
rect 6972 28024 6978 28076
rect 7147 28067 7205 28073
rect 7147 28033 7159 28067
rect 7193 28064 7205 28067
rect 7466 28064 7472 28076
rect 7193 28036 7472 28064
rect 7193 28033 7205 28036
rect 7147 28027 7205 28033
rect 7466 28024 7472 28036
rect 7524 28024 7530 28076
rect 8496 28073 8524 28104
rect 8938 28092 8944 28104
rect 8996 28092 9002 28144
rect 9125 28135 9183 28141
rect 9125 28101 9137 28135
rect 9171 28132 9183 28135
rect 9214 28132 9220 28144
rect 9171 28104 9220 28132
rect 9171 28101 9183 28104
rect 9125 28095 9183 28101
rect 9214 28092 9220 28104
rect 9272 28132 9278 28144
rect 9582 28132 9588 28144
rect 9272 28104 9588 28132
rect 9272 28092 9278 28104
rect 9582 28092 9588 28104
rect 9640 28092 9646 28144
rect 11974 28092 11980 28144
rect 12032 28132 12038 28144
rect 13924 28141 13952 28172
rect 14737 28169 14749 28172
rect 14783 28200 14795 28203
rect 15102 28200 15108 28212
rect 14783 28172 15108 28200
rect 14783 28169 14795 28172
rect 14737 28163 14795 28169
rect 15102 28160 15108 28172
rect 15160 28160 15166 28212
rect 16206 28160 16212 28212
rect 16264 28200 16270 28212
rect 23569 28203 23627 28209
rect 23569 28200 23581 28203
rect 16264 28172 23581 28200
rect 16264 28160 16270 28172
rect 23569 28169 23581 28172
rect 23615 28169 23627 28203
rect 23569 28163 23627 28169
rect 13909 28135 13967 28141
rect 12032 28104 13676 28132
rect 12032 28092 12038 28104
rect 8297 28067 8355 28073
rect 8297 28033 8309 28067
rect 8343 28033 8355 28067
rect 8297 28027 8355 28033
rect 8481 28067 8539 28073
rect 8481 28033 8493 28067
rect 8527 28064 8539 28067
rect 9398 28064 9404 28076
rect 8527 28036 9404 28064
rect 8527 28033 8539 28036
rect 8481 28027 8539 28033
rect 2406 27956 2412 28008
rect 2464 27996 2470 28008
rect 2501 27999 2559 28005
rect 2501 27996 2513 27999
rect 2464 27968 2513 27996
rect 2464 27956 2470 27968
rect 2501 27965 2513 27968
rect 2547 27965 2559 27999
rect 8312 27996 8340 28027
rect 9398 28024 9404 28036
rect 9456 28024 9462 28076
rect 11698 28064 11704 28076
rect 11659 28036 11704 28064
rect 11698 28024 11704 28036
rect 11756 28024 11762 28076
rect 12986 28024 12992 28076
rect 13044 28064 13050 28076
rect 13648 28073 13676 28104
rect 13909 28101 13921 28135
rect 13955 28101 13967 28135
rect 13909 28095 13967 28101
rect 14826 28092 14832 28144
rect 14884 28132 14890 28144
rect 22278 28132 22284 28144
rect 14884 28104 16160 28132
rect 14884 28092 14890 28104
rect 13541 28067 13599 28073
rect 13541 28064 13553 28067
rect 13044 28036 13553 28064
rect 13044 28024 13050 28036
rect 13541 28033 13553 28036
rect 13587 28033 13599 28067
rect 13541 28027 13599 28033
rect 13634 28067 13692 28073
rect 13634 28033 13646 28067
rect 13680 28033 13692 28067
rect 13634 28027 13692 28033
rect 13817 28067 13875 28073
rect 13817 28033 13829 28067
rect 13863 28033 13875 28067
rect 13817 28027 13875 28033
rect 9306 27996 9312 28008
rect 8312 27968 9312 27996
rect 2501 27959 2559 27965
rect 9306 27956 9312 27968
rect 9364 27996 9370 28008
rect 10689 27999 10747 28005
rect 10689 27996 10701 27999
rect 9364 27968 10701 27996
rect 9364 27956 9370 27968
rect 10689 27965 10701 27968
rect 10735 27965 10747 27999
rect 10689 27959 10747 27965
rect 10965 27999 11023 28005
rect 10965 27965 10977 27999
rect 11011 27996 11023 27999
rect 11146 27996 11152 28008
rect 11011 27968 11152 27996
rect 11011 27965 11023 27968
rect 10965 27959 11023 27965
rect 11146 27956 11152 27968
rect 11204 27956 11210 28008
rect 11885 27999 11943 28005
rect 11885 27965 11897 27999
rect 11931 27965 11943 27999
rect 11885 27959 11943 27965
rect 7285 27931 7343 27937
rect 7285 27897 7297 27931
rect 7331 27928 7343 27931
rect 11900 27928 11928 27959
rect 12342 27956 12348 28008
rect 12400 27996 12406 28008
rect 13832 27996 13860 28027
rect 13998 28024 14004 28076
rect 14056 28073 14062 28076
rect 14056 28064 14064 28073
rect 14056 28036 14101 28064
rect 14056 28027 14064 28036
rect 14056 28024 14062 28027
rect 15562 28024 15568 28076
rect 15620 28064 15626 28076
rect 16132 28073 16160 28104
rect 21468 28104 22284 28132
rect 21468 28076 21496 28104
rect 22278 28092 22284 28104
rect 22336 28092 22342 28144
rect 15850 28067 15908 28073
rect 15850 28064 15862 28067
rect 15620 28036 15862 28064
rect 15620 28024 15626 28036
rect 15850 28033 15862 28036
rect 15896 28033 15908 28067
rect 15850 28027 15908 28033
rect 16117 28067 16175 28073
rect 16117 28033 16129 28067
rect 16163 28033 16175 28067
rect 16117 28027 16175 28033
rect 18325 28067 18383 28073
rect 18325 28033 18337 28067
rect 18371 28064 18383 28067
rect 19334 28064 19340 28076
rect 18371 28036 19340 28064
rect 18371 28033 18383 28036
rect 18325 28027 18383 28033
rect 19334 28024 19340 28036
rect 19392 28024 19398 28076
rect 19705 28067 19763 28073
rect 19705 28033 19717 28067
rect 19751 28064 19763 28067
rect 20070 28064 20076 28076
rect 19751 28036 20076 28064
rect 19751 28033 19763 28036
rect 19705 28027 19763 28033
rect 20070 28024 20076 28036
rect 20128 28064 20134 28076
rect 21450 28064 21456 28076
rect 20128 28036 21456 28064
rect 20128 28024 20134 28036
rect 21450 28024 21456 28036
rect 21508 28024 21514 28076
rect 23584 28064 23612 28163
rect 23750 28160 23756 28212
rect 23808 28200 23814 28212
rect 24305 28203 24363 28209
rect 24305 28200 24317 28203
rect 23808 28172 24317 28200
rect 23808 28160 23814 28172
rect 24305 28169 24317 28172
rect 24351 28200 24363 28203
rect 33686 28200 33692 28212
rect 24351 28172 33692 28200
rect 24351 28169 24363 28172
rect 24305 28163 24363 28169
rect 33686 28160 33692 28172
rect 33744 28200 33750 28212
rect 35986 28200 35992 28212
rect 33744 28172 35992 28200
rect 33744 28160 33750 28172
rect 35986 28160 35992 28172
rect 36044 28160 36050 28212
rect 36354 28200 36360 28212
rect 36315 28172 36360 28200
rect 36354 28160 36360 28172
rect 36412 28160 36418 28212
rect 34241 28135 34299 28141
rect 34241 28101 34253 28135
rect 34287 28132 34299 28135
rect 36170 28132 36176 28144
rect 34287 28104 36176 28132
rect 34287 28101 34299 28104
rect 34241 28095 34299 28101
rect 36170 28092 36176 28104
rect 36228 28092 36234 28144
rect 24121 28067 24179 28073
rect 24121 28064 24133 28067
rect 23584 28036 24133 28064
rect 24121 28033 24133 28036
rect 24167 28064 24179 28067
rect 26878 28064 26884 28076
rect 24167 28036 26884 28064
rect 24167 28033 24179 28036
rect 24121 28027 24179 28033
rect 26878 28024 26884 28036
rect 26936 28024 26942 28076
rect 29730 28024 29736 28076
rect 29788 28064 29794 28076
rect 30009 28067 30067 28073
rect 30009 28064 30021 28067
rect 29788 28036 30021 28064
rect 29788 28024 29794 28036
rect 30009 28033 30021 28036
rect 30055 28033 30067 28067
rect 30009 28027 30067 28033
rect 30193 28067 30251 28073
rect 30193 28033 30205 28067
rect 30239 28064 30251 28067
rect 30742 28064 30748 28076
rect 30239 28036 30748 28064
rect 30239 28033 30251 28036
rect 30193 28027 30251 28033
rect 12400 27968 13860 27996
rect 14016 27968 15148 27996
rect 12400 27956 12406 27968
rect 12437 27931 12495 27937
rect 12437 27928 12449 27931
rect 7331 27900 9352 27928
rect 11900 27900 12449 27928
rect 7331 27897 7343 27900
rect 7285 27891 7343 27897
rect 9324 27872 9352 27900
rect 12437 27897 12449 27900
rect 12483 27928 12495 27931
rect 14016 27928 14044 27968
rect 14918 27928 14924 27940
rect 12483 27900 14044 27928
rect 14108 27900 14924 27928
rect 12483 27897 12495 27900
rect 12437 27891 12495 27897
rect 9306 27820 9312 27872
rect 9364 27820 9370 27872
rect 9858 27820 9864 27872
rect 9916 27860 9922 27872
rect 14108 27860 14136 27900
rect 14918 27888 14924 27900
rect 14976 27888 14982 27940
rect 15120 27928 15148 27968
rect 16666 27956 16672 28008
rect 16724 27996 16730 28008
rect 18049 27999 18107 28005
rect 18049 27996 18061 27999
rect 16724 27968 18061 27996
rect 16724 27956 16730 27968
rect 18049 27965 18061 27968
rect 18095 27965 18107 27999
rect 18049 27959 18107 27965
rect 19429 27999 19487 28005
rect 19429 27965 19441 27999
rect 19475 27965 19487 27999
rect 30208 27996 30236 28027
rect 30742 28024 30748 28036
rect 30800 28024 30806 28076
rect 31297 28067 31355 28073
rect 31297 28033 31309 28067
rect 31343 28064 31355 28067
rect 32766 28064 32772 28076
rect 31343 28036 32772 28064
rect 31343 28033 31355 28036
rect 31297 28027 31355 28033
rect 32766 28024 32772 28036
rect 32824 28024 32830 28076
rect 34146 28064 34152 28076
rect 34107 28036 34152 28064
rect 34146 28024 34152 28036
rect 34204 28024 34210 28076
rect 34333 28067 34391 28073
rect 34333 28033 34345 28067
rect 34379 28064 34391 28067
rect 34422 28064 34428 28076
rect 34379 28036 34428 28064
rect 34379 28033 34391 28036
rect 34333 28027 34391 28033
rect 34422 28024 34428 28036
rect 34480 28024 34486 28076
rect 34517 28067 34575 28073
rect 34517 28033 34529 28067
rect 34563 28064 34575 28067
rect 34698 28064 34704 28076
rect 34563 28036 34704 28064
rect 34563 28033 34575 28036
rect 34517 28027 34575 28033
rect 34698 28024 34704 28036
rect 34756 28024 34762 28076
rect 35342 28024 35348 28076
rect 35400 28064 35406 28076
rect 35989 28067 36047 28073
rect 35989 28064 36001 28067
rect 35400 28036 36001 28064
rect 35400 28024 35406 28036
rect 35989 28033 36001 28036
rect 36035 28033 36047 28067
rect 35989 28027 36047 28033
rect 31570 27996 31576 28008
rect 19429 27959 19487 27965
rect 29472 27968 30236 27996
rect 31531 27968 31576 27996
rect 17770 27928 17776 27940
rect 15120 27900 15240 27928
rect 9916 27832 14136 27860
rect 14185 27863 14243 27869
rect 9916 27820 9922 27832
rect 14185 27829 14197 27863
rect 14231 27860 14243 27863
rect 15010 27860 15016 27872
rect 14231 27832 15016 27860
rect 14231 27829 14243 27832
rect 14185 27823 14243 27829
rect 15010 27820 15016 27832
rect 15068 27820 15074 27872
rect 15212 27860 15240 27900
rect 16684 27900 17776 27928
rect 16684 27860 16712 27900
rect 17770 27888 17776 27900
rect 17828 27888 17834 27940
rect 19444 27928 19472 27959
rect 20070 27928 20076 27940
rect 19444 27900 20076 27928
rect 20070 27888 20076 27900
rect 20128 27888 20134 27940
rect 22465 27931 22523 27937
rect 22465 27897 22477 27931
rect 22511 27928 22523 27931
rect 22646 27928 22652 27940
rect 22511 27900 22652 27928
rect 22511 27897 22523 27900
rect 22465 27891 22523 27897
rect 22646 27888 22652 27900
rect 22704 27888 22710 27940
rect 27890 27928 27896 27940
rect 23492 27900 27896 27928
rect 16850 27860 16856 27872
rect 15212 27832 16712 27860
rect 16811 27832 16856 27860
rect 16850 27820 16856 27832
rect 16908 27820 16914 27872
rect 17954 27820 17960 27872
rect 18012 27860 18018 27872
rect 23492 27860 23520 27900
rect 27890 27888 27896 27900
rect 27948 27888 27954 27940
rect 29472 27872 29500 27968
rect 31570 27956 31576 27968
rect 31628 27996 31634 28008
rect 32125 27999 32183 28005
rect 32125 27996 32137 27999
rect 31628 27968 32137 27996
rect 31628 27956 31634 27968
rect 32125 27965 32137 27968
rect 32171 27965 32183 27999
rect 32125 27959 32183 27965
rect 58158 27928 58164 27940
rect 58119 27900 58164 27928
rect 58158 27888 58164 27900
rect 58216 27888 58222 27940
rect 18012 27832 23520 27860
rect 24949 27863 25007 27869
rect 18012 27820 18018 27832
rect 24949 27829 24961 27863
rect 24995 27860 25007 27863
rect 25038 27860 25044 27872
rect 24995 27832 25044 27860
rect 24995 27829 25007 27832
rect 24949 27823 25007 27829
rect 25038 27820 25044 27832
rect 25096 27820 25102 27872
rect 29454 27860 29460 27872
rect 29415 27832 29460 27860
rect 29454 27820 29460 27832
rect 29512 27820 29518 27872
rect 30006 27820 30012 27872
rect 30064 27860 30070 27872
rect 30101 27863 30159 27869
rect 30101 27860 30113 27863
rect 30064 27832 30113 27860
rect 30064 27820 30070 27832
rect 30101 27829 30113 27832
rect 30147 27860 30159 27863
rect 30282 27860 30288 27872
rect 30147 27832 30288 27860
rect 30147 27829 30159 27832
rect 30101 27823 30159 27829
rect 30282 27820 30288 27832
rect 30340 27820 30346 27872
rect 33502 27820 33508 27872
rect 33560 27860 33566 27872
rect 33965 27863 34023 27869
rect 33965 27860 33977 27863
rect 33560 27832 33977 27860
rect 33560 27820 33566 27832
rect 33965 27829 33977 27832
rect 34011 27829 34023 27863
rect 33965 27823 34023 27829
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 11517 27659 11575 27665
rect 11517 27625 11529 27659
rect 11563 27656 11575 27659
rect 11698 27656 11704 27668
rect 11563 27628 11704 27656
rect 11563 27625 11575 27628
rect 11517 27619 11575 27625
rect 11698 27616 11704 27628
rect 11756 27616 11762 27668
rect 13538 27656 13544 27668
rect 12176 27628 13124 27656
rect 13499 27628 13544 27656
rect 5629 27591 5687 27597
rect 5629 27557 5641 27591
rect 5675 27588 5687 27591
rect 7742 27588 7748 27600
rect 5675 27560 7748 27588
rect 5675 27557 5687 27560
rect 5629 27551 5687 27557
rect 7742 27548 7748 27560
rect 7800 27548 7806 27600
rect 10965 27591 11023 27597
rect 10965 27557 10977 27591
rect 11011 27588 11023 27591
rect 12176 27588 12204 27628
rect 11011 27560 12204 27588
rect 13096 27588 13124 27628
rect 13538 27616 13544 27628
rect 13596 27616 13602 27668
rect 16850 27616 16856 27668
rect 16908 27656 16914 27668
rect 29454 27656 29460 27668
rect 16908 27628 29460 27656
rect 16908 27616 16914 27628
rect 13998 27588 14004 27600
rect 13096 27560 14004 27588
rect 11011 27557 11023 27560
rect 10965 27551 11023 27557
rect 13998 27548 14004 27560
rect 14056 27548 14062 27600
rect 15565 27591 15623 27597
rect 15565 27557 15577 27591
rect 15611 27588 15623 27591
rect 16758 27588 16764 27600
rect 15611 27560 16764 27588
rect 15611 27557 15623 27560
rect 15565 27551 15623 27557
rect 16758 27548 16764 27560
rect 16816 27548 16822 27600
rect 7466 27520 7472 27532
rect 6656 27492 7472 27520
rect 4982 27452 4988 27464
rect 4943 27424 4988 27452
rect 4982 27412 4988 27424
rect 5040 27412 5046 27464
rect 5078 27455 5136 27461
rect 5078 27421 5090 27455
rect 5124 27421 5136 27455
rect 5350 27452 5356 27464
rect 5311 27424 5356 27452
rect 5078 27415 5136 27421
rect 3970 27344 3976 27396
rect 4028 27384 4034 27396
rect 5092 27384 5120 27415
rect 5350 27412 5356 27424
rect 5408 27412 5414 27464
rect 5442 27412 5448 27464
rect 5500 27461 5506 27464
rect 5500 27455 5549 27461
rect 5500 27421 5503 27455
rect 5537 27452 5549 27455
rect 6656 27452 6684 27492
rect 7466 27480 7472 27492
rect 7524 27480 7530 27532
rect 8294 27480 8300 27532
rect 8352 27520 8358 27532
rect 9033 27523 9091 27529
rect 9033 27520 9045 27523
rect 8352 27492 9045 27520
rect 8352 27480 8358 27492
rect 9033 27489 9045 27492
rect 9079 27520 9091 27523
rect 9861 27523 9919 27529
rect 9079 27492 9812 27520
rect 9079 27489 9091 27492
rect 9033 27483 9091 27489
rect 5537 27424 6684 27452
rect 5537 27421 5549 27424
rect 5500 27415 5549 27421
rect 5500 27412 5506 27415
rect 6730 27412 6736 27464
rect 6788 27452 6794 27464
rect 7561 27455 7619 27461
rect 7561 27452 7573 27455
rect 6788 27424 7573 27452
rect 6788 27412 6794 27424
rect 7561 27421 7573 27424
rect 7607 27421 7619 27455
rect 9490 27452 9496 27464
rect 9451 27424 9496 27452
rect 7561 27415 7619 27421
rect 9490 27412 9496 27424
rect 9548 27412 9554 27464
rect 9784 27461 9812 27492
rect 9861 27489 9873 27523
rect 9907 27520 9919 27523
rect 10226 27520 10232 27532
rect 9907 27492 10232 27520
rect 9907 27489 9919 27492
rect 9861 27483 9919 27489
rect 10226 27480 10232 27492
rect 10284 27480 10290 27532
rect 12158 27520 12164 27532
rect 12119 27492 12164 27520
rect 12158 27480 12164 27492
rect 12216 27480 12222 27532
rect 16868 27520 16896 27616
rect 18064 27597 18092 27628
rect 29454 27616 29460 27628
rect 29512 27616 29518 27668
rect 32766 27616 32772 27668
rect 32824 27656 32830 27668
rect 33778 27656 33784 27668
rect 32824 27628 33784 27656
rect 32824 27616 32830 27628
rect 33778 27616 33784 27628
rect 33836 27656 33842 27668
rect 34422 27656 34428 27668
rect 33836 27628 34428 27656
rect 33836 27616 33842 27628
rect 34422 27616 34428 27628
rect 34480 27616 34486 27668
rect 35986 27656 35992 27668
rect 35947 27628 35992 27656
rect 35986 27616 35992 27628
rect 36044 27616 36050 27668
rect 18049 27591 18107 27597
rect 18049 27557 18061 27591
rect 18095 27557 18107 27591
rect 20254 27588 20260 27600
rect 20215 27560 20260 27588
rect 18049 27551 18107 27557
rect 20254 27548 20260 27560
rect 20312 27548 20318 27600
rect 24026 27588 24032 27600
rect 20916 27560 24032 27588
rect 16500 27492 16896 27520
rect 9769 27455 9827 27461
rect 9769 27421 9781 27455
rect 9815 27452 9827 27455
rect 12428 27455 12486 27461
rect 9815 27424 11560 27452
rect 9815 27421 9827 27424
rect 9769 27415 9827 27421
rect 4028 27356 5120 27384
rect 4028 27344 4034 27356
rect 5166 27344 5172 27396
rect 5224 27384 5230 27396
rect 5261 27387 5319 27393
rect 5261 27384 5273 27387
rect 5224 27356 5273 27384
rect 5224 27344 5230 27356
rect 5261 27353 5273 27356
rect 5307 27384 5319 27387
rect 6914 27384 6920 27396
rect 5307 27356 6920 27384
rect 5307 27353 5319 27356
rect 5261 27347 5319 27353
rect 6914 27344 6920 27356
rect 6972 27344 6978 27396
rect 7374 27384 7380 27396
rect 7335 27356 7380 27384
rect 7374 27344 7380 27356
rect 7432 27344 7438 27396
rect 7466 27344 7472 27396
rect 7524 27384 7530 27396
rect 9508 27384 9536 27412
rect 7524 27356 9536 27384
rect 7524 27344 7530 27356
rect 10226 27344 10232 27396
rect 10284 27384 10290 27396
rect 10781 27387 10839 27393
rect 10781 27384 10793 27387
rect 10284 27356 10793 27384
rect 10284 27344 10290 27356
rect 10781 27353 10793 27356
rect 10827 27353 10839 27387
rect 10781 27347 10839 27353
rect 2498 27276 2504 27328
rect 2556 27316 2562 27328
rect 3145 27319 3203 27325
rect 3145 27316 3157 27319
rect 2556 27288 3157 27316
rect 2556 27276 2562 27288
rect 3145 27285 3157 27288
rect 3191 27316 3203 27319
rect 3326 27316 3332 27328
rect 3191 27288 3332 27316
rect 3191 27285 3203 27288
rect 3145 27279 3203 27285
rect 3326 27276 3332 27288
rect 3384 27276 3390 27328
rect 3881 27319 3939 27325
rect 3881 27285 3893 27319
rect 3927 27316 3939 27319
rect 5626 27316 5632 27328
rect 3927 27288 5632 27316
rect 3927 27285 3939 27288
rect 3881 27279 3939 27285
rect 5626 27276 5632 27288
rect 5684 27276 5690 27328
rect 7745 27319 7803 27325
rect 7745 27285 7757 27319
rect 7791 27316 7803 27319
rect 8662 27316 8668 27328
rect 7791 27288 8668 27316
rect 7791 27285 7803 27288
rect 7745 27279 7803 27285
rect 8662 27276 8668 27288
rect 8720 27276 8726 27328
rect 11532 27316 11560 27424
rect 12428 27421 12440 27455
rect 12474 27452 12486 27455
rect 13170 27452 13176 27464
rect 12474 27424 13176 27452
rect 12474 27421 12486 27424
rect 12428 27415 12486 27421
rect 13170 27412 13176 27424
rect 13228 27412 13234 27464
rect 16500 27461 16528 27492
rect 16485 27455 16543 27461
rect 16485 27452 16497 27455
rect 14752 27424 16497 27452
rect 11609 27387 11667 27393
rect 11609 27353 11621 27387
rect 11655 27384 11667 27387
rect 12894 27384 12900 27396
rect 11655 27356 12900 27384
rect 11655 27353 11667 27356
rect 11609 27347 11667 27353
rect 12894 27344 12900 27356
rect 12952 27344 12958 27396
rect 14752 27316 14780 27424
rect 16485 27421 16497 27424
rect 16531 27421 16543 27455
rect 16485 27415 16543 27421
rect 16669 27455 16727 27461
rect 16669 27421 16681 27455
rect 16715 27452 16727 27455
rect 17034 27452 17040 27464
rect 16715 27424 17040 27452
rect 16715 27421 16727 27424
rect 16669 27415 16727 27421
rect 17034 27412 17040 27424
rect 17092 27412 17098 27464
rect 17405 27455 17463 27461
rect 17405 27421 17417 27455
rect 17451 27452 17463 27455
rect 17770 27452 17776 27464
rect 17451 27424 17776 27452
rect 17451 27421 17463 27424
rect 17405 27415 17463 27421
rect 17770 27412 17776 27424
rect 17828 27452 17834 27464
rect 17865 27455 17923 27461
rect 17865 27452 17877 27455
rect 17828 27424 17877 27452
rect 17828 27412 17834 27424
rect 17865 27421 17877 27424
rect 17911 27421 17923 27455
rect 20272 27452 20300 27548
rect 20809 27455 20867 27461
rect 20809 27452 20821 27455
rect 20272 27424 20821 27452
rect 17865 27415 17923 27421
rect 20809 27421 20821 27424
rect 20855 27421 20867 27455
rect 20809 27415 20867 27421
rect 14829 27387 14887 27393
rect 14829 27353 14841 27387
rect 14875 27384 14887 27387
rect 15378 27384 15384 27396
rect 14875 27356 15384 27384
rect 14875 27353 14887 27356
rect 14829 27347 14887 27353
rect 15378 27344 15384 27356
rect 15436 27344 15442 27396
rect 15746 27344 15752 27396
rect 15804 27384 15810 27396
rect 16577 27387 16635 27393
rect 16577 27384 16589 27387
rect 15804 27356 16589 27384
rect 15804 27344 15810 27356
rect 16577 27353 16589 27356
rect 16623 27384 16635 27387
rect 16623 27356 17448 27384
rect 16623 27353 16635 27356
rect 16577 27347 16635 27353
rect 11532 27288 14780 27316
rect 17420 27316 17448 27356
rect 17494 27344 17500 27396
rect 17552 27384 17558 27396
rect 20916 27384 20944 27560
rect 24026 27548 24032 27560
rect 24084 27548 24090 27600
rect 33134 27588 33140 27600
rect 32600 27560 33140 27588
rect 24762 27480 24768 27532
rect 24820 27520 24826 27532
rect 24820 27492 25360 27520
rect 24820 27480 24826 27492
rect 24946 27452 24952 27464
rect 17552 27356 20944 27384
rect 21008 27424 24952 27452
rect 17552 27344 17558 27356
rect 21008 27316 21036 27424
rect 24946 27412 24952 27424
rect 25004 27412 25010 27464
rect 25038 27412 25044 27464
rect 25096 27452 25102 27464
rect 25222 27452 25228 27464
rect 25096 27424 25141 27452
rect 25183 27424 25228 27452
rect 25096 27412 25102 27424
rect 25222 27412 25228 27424
rect 25280 27412 25286 27464
rect 25332 27461 25360 27492
rect 29730 27480 29736 27532
rect 29788 27520 29794 27532
rect 30377 27523 30435 27529
rect 30377 27520 30389 27523
rect 29788 27492 30389 27520
rect 29788 27480 29794 27492
rect 30377 27489 30389 27492
rect 30423 27489 30435 27523
rect 30377 27483 30435 27489
rect 25317 27455 25375 27461
rect 25317 27421 25329 27455
rect 25363 27421 25375 27455
rect 25317 27415 25375 27421
rect 25409 27455 25467 27461
rect 25409 27421 25421 27455
rect 25455 27421 25467 27455
rect 25409 27415 25467 27421
rect 26513 27455 26571 27461
rect 26513 27421 26525 27455
rect 26559 27452 26571 27455
rect 27614 27452 27620 27464
rect 26559 27424 27620 27452
rect 26559 27421 26571 27424
rect 26513 27415 26571 27421
rect 21726 27344 21732 27396
rect 21784 27384 21790 27396
rect 22557 27387 22615 27393
rect 22557 27384 22569 27387
rect 21784 27356 22569 27384
rect 21784 27344 21790 27356
rect 22557 27353 22569 27356
rect 22603 27384 22615 27387
rect 24026 27384 24032 27396
rect 22603 27356 24032 27384
rect 22603 27353 22615 27356
rect 22557 27347 22615 27353
rect 24026 27344 24032 27356
rect 24084 27344 24090 27396
rect 25424 27384 25452 27415
rect 27614 27412 27620 27424
rect 27672 27412 27678 27464
rect 30653 27455 30711 27461
rect 30653 27452 30665 27455
rect 29012 27424 30665 27452
rect 24504 27356 25452 27384
rect 25685 27387 25743 27393
rect 24504 27328 24532 27356
rect 25685 27353 25697 27387
rect 25731 27384 25743 27387
rect 26758 27387 26816 27393
rect 26758 27384 26770 27387
rect 25731 27356 26770 27384
rect 25731 27353 25743 27356
rect 25685 27347 25743 27353
rect 26758 27353 26770 27356
rect 26804 27353 26816 27387
rect 26758 27347 26816 27353
rect 28442 27344 28448 27396
rect 28500 27384 28506 27396
rect 29012 27393 29040 27424
rect 30653 27421 30665 27424
rect 30699 27452 30711 27455
rect 30926 27452 30932 27464
rect 30699 27424 30932 27452
rect 30699 27421 30711 27424
rect 30653 27415 30711 27421
rect 30926 27412 30932 27424
rect 30984 27452 30990 27464
rect 32600 27461 32628 27560
rect 33134 27548 33140 27560
rect 33192 27588 33198 27600
rect 34146 27588 34152 27600
rect 33192 27560 34152 27588
rect 33192 27548 33198 27560
rect 34146 27548 34152 27560
rect 34204 27548 34210 27600
rect 31113 27455 31171 27461
rect 31113 27452 31125 27455
rect 30984 27424 31125 27452
rect 30984 27412 30990 27424
rect 31113 27421 31125 27424
rect 31159 27421 31171 27455
rect 31113 27415 31171 27421
rect 31389 27455 31447 27461
rect 31389 27421 31401 27455
rect 31435 27452 31447 27455
rect 32585 27455 32643 27461
rect 32585 27452 32597 27455
rect 31435 27424 32597 27452
rect 31435 27421 31447 27424
rect 31389 27415 31447 27421
rect 32585 27421 32597 27424
rect 32631 27421 32643 27455
rect 32585 27415 32643 27421
rect 32677 27455 32735 27461
rect 32677 27421 32689 27455
rect 32723 27452 32735 27455
rect 32723 27424 32904 27452
rect 32723 27421 32735 27424
rect 32677 27415 32735 27421
rect 28997 27387 29055 27393
rect 28997 27384 29009 27387
rect 28500 27356 29009 27384
rect 28500 27344 28506 27356
rect 28997 27353 29009 27356
rect 29043 27353 29055 27387
rect 32766 27384 32772 27396
rect 32727 27356 32772 27384
rect 28997 27347 29055 27353
rect 32766 27344 32772 27356
rect 32824 27344 32830 27396
rect 32876 27384 32904 27424
rect 32950 27412 32956 27464
rect 33008 27452 33014 27464
rect 33008 27424 33053 27452
rect 33008 27412 33014 27424
rect 33226 27412 33232 27464
rect 33284 27452 33290 27464
rect 33781 27455 33839 27461
rect 33781 27452 33793 27455
rect 33284 27424 33793 27452
rect 33284 27412 33290 27424
rect 33781 27421 33793 27424
rect 33827 27452 33839 27455
rect 34422 27452 34428 27464
rect 33827 27424 34428 27452
rect 33827 27421 33839 27424
rect 33781 27415 33839 27421
rect 34422 27412 34428 27424
rect 34480 27412 34486 27464
rect 33597 27387 33655 27393
rect 33597 27384 33609 27387
rect 32876 27356 33609 27384
rect 33597 27353 33609 27356
rect 33643 27384 33655 27387
rect 33686 27384 33692 27396
rect 33643 27356 33692 27384
rect 33643 27353 33655 27356
rect 33597 27347 33655 27353
rect 33686 27344 33692 27356
rect 33744 27344 33750 27396
rect 24486 27316 24492 27328
rect 17420 27288 21036 27316
rect 24447 27288 24492 27316
rect 24486 27276 24492 27288
rect 24544 27276 24550 27328
rect 27893 27319 27951 27325
rect 27893 27285 27905 27319
rect 27939 27316 27951 27319
rect 28534 27316 28540 27328
rect 27939 27288 28540 27316
rect 27939 27285 27951 27288
rect 27893 27279 27951 27285
rect 28534 27276 28540 27288
rect 28592 27276 28598 27328
rect 32398 27316 32404 27328
rect 32359 27288 32404 27316
rect 32398 27276 32404 27288
rect 32456 27276 32462 27328
rect 32582 27276 32588 27328
rect 32640 27316 32646 27328
rect 33413 27319 33471 27325
rect 33413 27316 33425 27319
rect 32640 27288 33425 27316
rect 32640 27276 32646 27288
rect 33413 27285 33425 27288
rect 33459 27285 33471 27319
rect 33413 27279 33471 27285
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 3142 27112 3148 27124
rect 2973 27084 3148 27112
rect 2973 26991 3001 27084
rect 3142 27072 3148 27084
rect 3200 27072 3206 27124
rect 5074 27072 5080 27124
rect 5132 27072 5138 27124
rect 6365 27115 6423 27121
rect 6365 27081 6377 27115
rect 6411 27112 6423 27115
rect 6730 27112 6736 27124
rect 6411 27084 6736 27112
rect 6411 27081 6423 27084
rect 6365 27075 6423 27081
rect 6730 27072 6736 27084
rect 6788 27072 6794 27124
rect 7926 27072 7932 27124
rect 7984 27112 7990 27124
rect 9490 27112 9496 27124
rect 7984 27084 8616 27112
rect 9451 27084 9496 27112
rect 7984 27072 7990 27084
rect 5092 27044 5120 27072
rect 5261 27047 5319 27053
rect 5261 27044 5273 27047
rect 3896 27016 5028 27044
rect 5092 27016 5273 27044
rect 2498 26936 2504 26988
rect 2556 26976 2562 26988
rect 2958 26985 3016 26991
rect 3896 26988 3924 27016
rect 2869 26979 2927 26985
rect 2869 26976 2881 26979
rect 2556 26948 2881 26976
rect 2556 26936 2562 26948
rect 2869 26945 2881 26948
rect 2915 26945 2927 26979
rect 2958 26951 2970 26985
rect 3004 26951 3016 26985
rect 2958 26945 3016 26951
rect 3058 26979 3116 26985
rect 3058 26945 3070 26979
rect 3104 26945 3116 26979
rect 3234 26976 3240 26988
rect 3195 26948 3240 26976
rect 2869 26939 2927 26945
rect 3058 26939 3116 26945
rect 3068 26908 3096 26939
rect 3234 26936 3240 26948
rect 3292 26936 3298 26988
rect 3878 26976 3884 26988
rect 3839 26948 3884 26976
rect 3878 26936 3884 26948
rect 3936 26936 3942 26988
rect 4062 26976 4068 26988
rect 4023 26948 4068 26976
rect 4062 26936 4068 26948
rect 4120 26936 4126 26988
rect 4890 26976 4896 26988
rect 4851 26948 4896 26976
rect 4890 26936 4896 26948
rect 4948 26936 4954 26988
rect 5000 26985 5028 27016
rect 5261 27013 5273 27016
rect 5307 27013 5319 27047
rect 5261 27007 5319 27013
rect 7500 27047 7558 27053
rect 7500 27013 7512 27047
rect 7546 27044 7558 27047
rect 8205 27047 8263 27053
rect 8205 27044 8217 27047
rect 7546 27016 8217 27044
rect 7546 27013 7558 27016
rect 7500 27007 7558 27013
rect 8205 27013 8217 27016
rect 8251 27013 8263 27047
rect 8205 27007 8263 27013
rect 4986 26979 5044 26985
rect 4986 26945 4998 26979
rect 5032 26945 5044 26979
rect 5166 26976 5172 26988
rect 5127 26948 5172 26976
rect 4986 26939 5044 26945
rect 5166 26936 5172 26948
rect 5224 26936 5230 26988
rect 5442 26985 5448 26988
rect 5399 26979 5448 26985
rect 5399 26945 5411 26979
rect 5445 26945 5448 26979
rect 5399 26939 5448 26945
rect 5442 26936 5448 26939
rect 5500 26936 5506 26988
rect 6730 26936 6736 26988
rect 6788 26976 6794 26988
rect 7190 26976 7196 26988
rect 6788 26948 7196 26976
rect 6788 26936 6794 26948
rect 7190 26936 7196 26948
rect 7248 26936 7254 26988
rect 7926 26936 7932 26988
rect 7984 26976 7990 26988
rect 8588 26985 8616 27084
rect 9490 27072 9496 27084
rect 9548 27072 9554 27124
rect 16206 27072 16212 27124
rect 16264 27112 16270 27124
rect 17218 27112 17224 27124
rect 16264 27084 17224 27112
rect 16264 27072 16270 27084
rect 17218 27072 17224 27084
rect 17276 27072 17282 27124
rect 17770 27072 17776 27124
rect 17828 27112 17834 27124
rect 20806 27112 20812 27124
rect 17828 27084 20812 27112
rect 17828 27072 17834 27084
rect 20806 27072 20812 27084
rect 20864 27072 20870 27124
rect 23750 27072 23756 27124
rect 23808 27112 23814 27124
rect 29362 27112 29368 27124
rect 23808 27084 29368 27112
rect 23808 27072 23814 27084
rect 29362 27072 29368 27084
rect 29420 27072 29426 27124
rect 30926 27112 30932 27124
rect 30887 27084 30932 27112
rect 30926 27072 30932 27084
rect 30984 27072 30990 27124
rect 36078 27112 36084 27124
rect 33980 27084 36084 27112
rect 9585 27047 9643 27053
rect 9585 27013 9597 27047
rect 9631 27044 9643 27047
rect 10226 27044 10232 27056
rect 9631 27016 10232 27044
rect 9631 27013 9643 27016
rect 9585 27007 9643 27013
rect 10226 27004 10232 27016
rect 10284 27004 10290 27056
rect 21726 27044 21732 27056
rect 17144 27016 21732 27044
rect 8481 26979 8539 26985
rect 8481 26976 8493 26979
rect 7984 26948 8493 26976
rect 7984 26936 7990 26948
rect 8481 26945 8493 26948
rect 8527 26945 8539 26979
rect 8481 26939 8539 26945
rect 8573 26979 8631 26985
rect 8573 26945 8585 26979
rect 8619 26945 8631 26979
rect 8573 26939 8631 26945
rect 8662 26936 8668 26988
rect 8720 26976 8726 26988
rect 8849 26979 8907 26985
rect 8720 26948 8765 26976
rect 8720 26936 8726 26948
rect 8849 26945 8861 26979
rect 8895 26976 8907 26979
rect 9030 26976 9036 26988
rect 8895 26948 9036 26976
rect 8895 26945 8907 26948
rect 8849 26939 8907 26945
rect 9030 26936 9036 26948
rect 9088 26936 9094 26988
rect 10137 26979 10195 26985
rect 10137 26945 10149 26979
rect 10183 26976 10195 26979
rect 10870 26976 10876 26988
rect 10183 26948 10876 26976
rect 10183 26945 10195 26948
rect 10137 26939 10195 26945
rect 10870 26936 10876 26948
rect 10928 26936 10934 26988
rect 11885 26979 11943 26985
rect 11885 26945 11897 26979
rect 11931 26976 11943 26979
rect 12526 26976 12532 26988
rect 11931 26948 12532 26976
rect 11931 26945 11943 26948
rect 11885 26939 11943 26945
rect 12526 26936 12532 26948
rect 12584 26936 12590 26988
rect 12802 26936 12808 26988
rect 12860 26976 12866 26988
rect 17144 26985 17172 27016
rect 13173 26979 13231 26985
rect 13173 26976 13185 26979
rect 12860 26948 13185 26976
rect 12860 26936 12866 26948
rect 13173 26945 13185 26948
rect 13219 26945 13231 26979
rect 13173 26939 13231 26945
rect 17129 26979 17187 26985
rect 17129 26945 17141 26979
rect 17175 26945 17187 26979
rect 17129 26939 17187 26945
rect 17396 26979 17454 26985
rect 17396 26945 17408 26979
rect 17442 26976 17454 26979
rect 17678 26976 17684 26988
rect 17442 26948 17684 26976
rect 17442 26945 17454 26948
rect 17396 26939 17454 26945
rect 17678 26936 17684 26948
rect 17736 26936 17742 26988
rect 18984 26985 19012 27016
rect 21726 27004 21732 27016
rect 21784 27004 21790 27056
rect 25406 27004 25412 27056
rect 25464 27044 25470 27056
rect 29546 27044 29552 27056
rect 25464 27016 29552 27044
rect 25464 27004 25470 27016
rect 29546 27004 29552 27016
rect 29604 27004 29610 27056
rect 29733 27047 29791 27053
rect 29733 27013 29745 27047
rect 29779 27044 29791 27047
rect 31754 27044 31760 27056
rect 29779 27016 31760 27044
rect 29779 27013 29791 27016
rect 29733 27007 29791 27013
rect 31754 27004 31760 27016
rect 31812 27044 31818 27056
rect 33980 27044 34008 27084
rect 36078 27072 36084 27084
rect 36136 27072 36142 27124
rect 35345 27047 35403 27053
rect 35345 27044 35357 27047
rect 31812 27016 34008 27044
rect 31812 27004 31818 27016
rect 19242 26985 19248 26988
rect 18969 26979 19027 26985
rect 18969 26945 18981 26979
rect 19015 26945 19027 26979
rect 18969 26939 19027 26945
rect 19236 26939 19248 26985
rect 19300 26976 19306 26988
rect 19300 26948 19336 26976
rect 19242 26936 19248 26939
rect 19300 26936 19306 26948
rect 20806 26936 20812 26988
rect 20864 26976 20870 26988
rect 20993 26979 21051 26985
rect 20993 26976 21005 26979
rect 20864 26948 21005 26976
rect 20864 26936 20870 26948
rect 20993 26945 21005 26948
rect 21039 26945 21051 26979
rect 20993 26939 21051 26945
rect 21821 26979 21879 26985
rect 21821 26945 21833 26979
rect 21867 26945 21879 26979
rect 21821 26939 21879 26945
rect 22005 26979 22063 26985
rect 22005 26945 22017 26979
rect 22051 26945 22063 26979
rect 22005 26939 22063 26945
rect 3697 26911 3755 26917
rect 3697 26908 3709 26911
rect 3068 26880 3709 26908
rect 3697 26877 3709 26880
rect 3743 26877 3755 26911
rect 3697 26871 3755 26877
rect 7745 26911 7803 26917
rect 7745 26877 7757 26911
rect 7791 26877 7803 26911
rect 7745 26871 7803 26877
rect 7760 26840 7788 26871
rect 9582 26868 9588 26920
rect 9640 26908 9646 26920
rect 10413 26911 10471 26917
rect 10413 26908 10425 26911
rect 9640 26880 10425 26908
rect 9640 26868 9646 26880
rect 10413 26877 10425 26880
rect 10459 26877 10471 26911
rect 10413 26871 10471 26877
rect 11146 26868 11152 26920
rect 11204 26908 11210 26920
rect 11609 26911 11667 26917
rect 11609 26908 11621 26911
rect 11204 26880 11621 26908
rect 11204 26868 11210 26880
rect 11609 26877 11621 26880
rect 11655 26877 11667 26911
rect 12894 26908 12900 26920
rect 12807 26880 12900 26908
rect 11609 26871 11667 26877
rect 12894 26868 12900 26880
rect 12952 26908 12958 26920
rect 13630 26908 13636 26920
rect 12952 26880 13636 26908
rect 12952 26868 12958 26880
rect 13630 26868 13636 26880
rect 13688 26868 13694 26920
rect 20162 26868 20168 26920
rect 20220 26908 20226 26920
rect 20438 26908 20444 26920
rect 20220 26880 20444 26908
rect 20220 26868 20226 26880
rect 20438 26868 20444 26880
rect 20496 26868 20502 26920
rect 20898 26868 20904 26920
rect 20956 26908 20962 26920
rect 21836 26908 21864 26939
rect 20956 26880 21864 26908
rect 22020 26908 22048 26939
rect 22462 26936 22468 26988
rect 22520 26976 22526 26988
rect 23762 26979 23820 26985
rect 23762 26976 23774 26979
rect 22520 26948 23774 26976
rect 22520 26936 22526 26948
rect 23762 26945 23774 26948
rect 23808 26945 23820 26979
rect 24026 26976 24032 26988
rect 23939 26948 24032 26976
rect 23762 26939 23820 26945
rect 24026 26936 24032 26948
rect 24084 26976 24090 26988
rect 25314 26985 25320 26988
rect 25041 26979 25099 26985
rect 25041 26976 25053 26979
rect 24084 26948 25053 26976
rect 24084 26936 24090 26948
rect 25041 26945 25053 26948
rect 25087 26945 25099 26979
rect 25041 26939 25099 26945
rect 25308 26939 25320 26985
rect 25372 26976 25378 26988
rect 25372 26948 25408 26976
rect 25314 26936 25320 26939
rect 25372 26936 25378 26948
rect 26418 26936 26424 26988
rect 26476 26976 26482 26988
rect 28149 26979 28207 26985
rect 28149 26976 28161 26979
rect 26476 26948 28161 26976
rect 26476 26936 26482 26948
rect 28149 26945 28161 26948
rect 28195 26945 28207 26979
rect 28149 26939 28207 26945
rect 29638 26936 29644 26988
rect 29696 26976 29702 26988
rect 32416 26985 32444 27016
rect 29917 26979 29975 26985
rect 29917 26976 29929 26979
rect 29696 26948 29929 26976
rect 29696 26936 29702 26948
rect 29917 26945 29929 26948
rect 29963 26945 29975 26979
rect 29917 26939 29975 26945
rect 32401 26979 32459 26985
rect 32401 26945 32413 26979
rect 32447 26945 32459 26979
rect 32582 26976 32588 26988
rect 32543 26948 32588 26976
rect 32401 26939 32459 26945
rect 32582 26936 32588 26948
rect 32640 26936 32646 26988
rect 32677 26979 32735 26985
rect 32677 26945 32689 26979
rect 32723 26945 32735 26979
rect 32677 26939 32735 26945
rect 22020 26880 22692 26908
rect 20956 26868 20962 26880
rect 12158 26840 12164 26852
rect 7760 26812 12164 26840
rect 12158 26800 12164 26812
rect 12216 26800 12222 26852
rect 20349 26843 20407 26849
rect 20349 26809 20361 26843
rect 20395 26840 20407 26843
rect 21910 26840 21916 26852
rect 20395 26812 21916 26840
rect 20395 26809 20407 26812
rect 20349 26803 20407 26809
rect 20456 26784 20484 26812
rect 21910 26800 21916 26812
rect 21968 26800 21974 26852
rect 2593 26775 2651 26781
rect 2593 26741 2605 26775
rect 2639 26772 2651 26775
rect 2774 26772 2780 26784
rect 2639 26744 2780 26772
rect 2639 26741 2651 26744
rect 2593 26735 2651 26741
rect 2774 26732 2780 26744
rect 2832 26732 2838 26784
rect 5537 26775 5595 26781
rect 5537 26741 5549 26775
rect 5583 26772 5595 26775
rect 6822 26772 6828 26784
rect 5583 26744 6828 26772
rect 5583 26741 5595 26744
rect 5537 26735 5595 26741
rect 6822 26732 6828 26744
rect 6880 26732 6886 26784
rect 18509 26775 18567 26781
rect 18509 26741 18521 26775
rect 18555 26772 18567 26775
rect 19334 26772 19340 26784
rect 18555 26744 19340 26772
rect 18555 26741 18567 26744
rect 18509 26735 18567 26741
rect 19334 26732 19340 26744
rect 19392 26732 19398 26784
rect 20438 26732 20444 26784
rect 20496 26732 20502 26784
rect 21174 26772 21180 26784
rect 21135 26744 21180 26772
rect 21174 26732 21180 26744
rect 21232 26732 21238 26784
rect 22002 26732 22008 26784
rect 22060 26772 22066 26784
rect 22664 26781 22692 26880
rect 27614 26868 27620 26920
rect 27672 26908 27678 26920
rect 27893 26911 27951 26917
rect 27893 26908 27905 26911
rect 27672 26880 27905 26908
rect 27672 26868 27678 26880
rect 27893 26877 27905 26880
rect 27939 26877 27951 26911
rect 27893 26871 27951 26877
rect 30282 26868 30288 26920
rect 30340 26908 30346 26920
rect 32692 26908 32720 26939
rect 32766 26936 32772 26988
rect 32824 26976 32830 26988
rect 33873 26979 33931 26985
rect 32824 26948 32869 26976
rect 32824 26936 32830 26948
rect 33873 26945 33885 26979
rect 33919 26976 33931 26979
rect 33980 26976 34008 27016
rect 34072 27016 35357 27044
rect 34072 26985 34100 27016
rect 35345 27013 35357 27016
rect 35391 27013 35403 27047
rect 35345 27007 35403 27013
rect 33919 26948 34008 26976
rect 34057 26979 34115 26985
rect 33919 26945 33931 26948
rect 33873 26939 33931 26945
rect 34057 26945 34069 26979
rect 34103 26945 34115 26979
rect 34057 26939 34115 26945
rect 34146 26936 34152 26988
rect 34204 26976 34210 26988
rect 34287 26979 34345 26985
rect 34204 26948 34249 26976
rect 34204 26936 34210 26948
rect 34287 26945 34299 26979
rect 34333 26976 34345 26979
rect 34422 26976 34428 26988
rect 34333 26948 34428 26976
rect 34333 26945 34345 26948
rect 34287 26939 34345 26945
rect 34422 26936 34428 26948
rect 34480 26936 34486 26988
rect 34514 26936 34520 26988
rect 34572 26976 34578 26988
rect 34977 26979 35035 26985
rect 34977 26976 34989 26979
rect 34572 26948 34989 26976
rect 34572 26936 34578 26948
rect 34977 26945 34989 26948
rect 35023 26945 35035 26979
rect 34977 26939 35035 26945
rect 35161 26979 35219 26985
rect 35161 26945 35173 26979
rect 35207 26976 35219 26979
rect 35434 26976 35440 26988
rect 35207 26948 35440 26976
rect 35207 26945 35219 26948
rect 35161 26939 35219 26945
rect 35434 26936 35440 26948
rect 35492 26936 35498 26988
rect 38657 26979 38715 26985
rect 38657 26945 38669 26979
rect 38703 26976 38715 26979
rect 39117 26979 39175 26985
rect 39117 26976 39129 26979
rect 38703 26948 39129 26976
rect 38703 26945 38715 26948
rect 38657 26939 38715 26945
rect 39117 26945 39129 26948
rect 39163 26945 39175 26979
rect 39117 26939 39175 26945
rect 30340 26880 32720 26908
rect 30340 26868 30346 26880
rect 32692 26840 32720 26880
rect 33962 26868 33968 26920
rect 34020 26908 34026 26920
rect 38672 26908 38700 26939
rect 34020 26880 38700 26908
rect 34020 26868 34026 26880
rect 34146 26840 34152 26852
rect 32692 26812 34152 26840
rect 34146 26800 34152 26812
rect 34204 26800 34210 26852
rect 22189 26775 22247 26781
rect 22189 26772 22201 26775
rect 22060 26744 22201 26772
rect 22060 26732 22066 26744
rect 22189 26741 22201 26744
rect 22235 26741 22247 26775
rect 22189 26735 22247 26741
rect 22649 26775 22707 26781
rect 22649 26741 22661 26775
rect 22695 26772 22707 26775
rect 23106 26772 23112 26784
rect 22695 26744 23112 26772
rect 22695 26741 22707 26744
rect 22649 26735 22707 26741
rect 23106 26732 23112 26744
rect 23164 26732 23170 26784
rect 26234 26732 26240 26784
rect 26292 26772 26298 26784
rect 26421 26775 26479 26781
rect 26421 26772 26433 26775
rect 26292 26744 26433 26772
rect 26292 26732 26298 26744
rect 26421 26741 26433 26744
rect 26467 26741 26479 26775
rect 29270 26772 29276 26784
rect 29231 26744 29276 26772
rect 26421 26735 26479 26741
rect 29270 26732 29276 26744
rect 29328 26732 29334 26784
rect 33045 26775 33103 26781
rect 33045 26741 33057 26775
rect 33091 26772 33103 26775
rect 33226 26772 33232 26784
rect 33091 26744 33232 26772
rect 33091 26741 33103 26744
rect 33045 26735 33103 26741
rect 33226 26732 33232 26744
rect 33284 26732 33290 26784
rect 34514 26772 34520 26784
rect 34475 26744 34520 26772
rect 34514 26732 34520 26744
rect 34572 26732 34578 26784
rect 39942 26732 39948 26784
rect 40000 26772 40006 26784
rect 40405 26775 40463 26781
rect 40405 26772 40417 26775
rect 40000 26744 40417 26772
rect 40000 26732 40006 26744
rect 40405 26741 40417 26744
rect 40451 26741 40463 26775
rect 58158 26772 58164 26784
rect 58119 26744 58164 26772
rect 40405 26735 40463 26741
rect 58158 26732 58164 26744
rect 58216 26732 58222 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 7374 26568 7380 26580
rect 6104 26540 7380 26568
rect 3970 26460 3976 26512
rect 4028 26460 4034 26512
rect 2133 26367 2191 26373
rect 2133 26333 2145 26367
rect 2179 26364 2191 26367
rect 2866 26364 2872 26376
rect 2179 26336 2872 26364
rect 2179 26333 2191 26336
rect 2133 26327 2191 26333
rect 2866 26324 2872 26336
rect 2924 26324 2930 26376
rect 2961 26364 3019 26370
rect 2961 26330 2973 26364
rect 3007 26330 3019 26364
rect 2961 26324 3019 26330
rect 3053 26367 3111 26373
rect 3053 26333 3065 26367
rect 3099 26333 3111 26367
rect 3053 26327 3111 26333
rect 2593 26299 2651 26305
rect 2593 26265 2605 26299
rect 2639 26296 2651 26299
rect 2639 26268 2774 26296
rect 2639 26265 2651 26268
rect 2593 26259 2651 26265
rect 2746 26228 2774 26268
rect 2866 26228 2872 26240
rect 2746 26200 2872 26228
rect 2866 26188 2872 26200
rect 2924 26188 2930 26240
rect 2976 26228 3004 26324
rect 3068 26296 3096 26327
rect 3234 26324 3240 26376
rect 3292 26364 3298 26376
rect 3988 26373 4016 26460
rect 3973 26367 4031 26373
rect 3292 26336 3924 26364
rect 3292 26324 3298 26336
rect 3789 26299 3847 26305
rect 3789 26296 3801 26299
rect 3068 26268 3801 26296
rect 3789 26265 3801 26268
rect 3835 26265 3847 26299
rect 3896 26296 3924 26336
rect 3973 26333 3985 26367
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 4062 26324 4068 26376
rect 4120 26364 4126 26376
rect 4157 26367 4215 26373
rect 4157 26364 4169 26367
rect 4120 26336 4169 26364
rect 4120 26324 4126 26336
rect 4157 26333 4169 26336
rect 4203 26364 4215 26367
rect 5997 26367 6055 26373
rect 5997 26364 6009 26367
rect 4203 26336 6009 26364
rect 4203 26333 4215 26336
rect 4157 26327 4215 26333
rect 5997 26333 6009 26336
rect 6043 26364 6055 26367
rect 6104 26364 6132 26540
rect 7374 26528 7380 26540
rect 7432 26528 7438 26580
rect 9493 26571 9551 26577
rect 9493 26537 9505 26571
rect 9539 26568 9551 26571
rect 9674 26568 9680 26580
rect 9539 26540 9680 26568
rect 9539 26537 9551 26540
rect 9493 26531 9551 26537
rect 9674 26528 9680 26540
rect 9732 26528 9738 26580
rect 11425 26571 11483 26577
rect 11425 26537 11437 26571
rect 11471 26568 11483 26571
rect 12342 26568 12348 26580
rect 11471 26540 12348 26568
rect 11471 26537 11483 26540
rect 11425 26531 11483 26537
rect 12342 26528 12348 26540
rect 12400 26528 12406 26580
rect 17221 26571 17279 26577
rect 17221 26537 17233 26571
rect 17267 26568 17279 26571
rect 17494 26568 17500 26580
rect 17267 26540 17500 26568
rect 17267 26537 17279 26540
rect 17221 26531 17279 26537
rect 17494 26528 17500 26540
rect 17552 26528 17558 26580
rect 18693 26571 18751 26577
rect 18693 26537 18705 26571
rect 18739 26568 18751 26571
rect 19242 26568 19248 26580
rect 18739 26540 19248 26568
rect 18739 26537 18751 26540
rect 18693 26531 18751 26537
rect 19242 26528 19248 26540
rect 19300 26528 19306 26580
rect 22462 26568 22468 26580
rect 21192 26540 22324 26568
rect 22423 26540 22468 26568
rect 6914 26460 6920 26512
rect 6972 26500 6978 26512
rect 7469 26503 7527 26509
rect 6972 26472 7328 26500
rect 6972 26460 6978 26472
rect 7300 26432 7328 26472
rect 7469 26469 7481 26503
rect 7515 26500 7527 26503
rect 7650 26500 7656 26512
rect 7515 26472 7656 26500
rect 7515 26469 7527 26472
rect 7469 26463 7527 26469
rect 7650 26460 7656 26472
rect 7708 26460 7714 26512
rect 10594 26460 10600 26512
rect 10652 26500 10658 26512
rect 21192 26500 21220 26540
rect 22296 26500 22324 26540
rect 22462 26528 22468 26540
rect 22520 26528 22526 26580
rect 24670 26528 24676 26580
rect 24728 26568 24734 26580
rect 25314 26568 25320 26580
rect 24728 26540 25176 26568
rect 25275 26540 25320 26568
rect 24728 26528 24734 26540
rect 24302 26500 24308 26512
rect 10652 26472 21220 26500
rect 21284 26472 22232 26500
rect 22296 26472 24308 26500
rect 10652 26460 10658 26472
rect 7208 26404 9628 26432
rect 6043 26336 6132 26364
rect 6043 26333 6055 26336
rect 5997 26327 6055 26333
rect 6730 26324 6736 26376
rect 6788 26364 6794 26376
rect 6988 26373 7052 26374
rect 6832 26367 6890 26373
rect 6832 26364 6844 26367
rect 6788 26336 6844 26364
rect 6788 26324 6794 26336
rect 6832 26333 6844 26336
rect 6878 26333 6890 26367
rect 6832 26327 6890 26333
rect 6973 26367 7052 26373
rect 6973 26333 6985 26367
rect 7019 26333 7052 26367
rect 6973 26327 7052 26333
rect 7101 26367 7159 26373
rect 7101 26333 7113 26367
rect 7147 26364 7159 26367
rect 7208 26364 7236 26404
rect 9600 26376 9628 26404
rect 9766 26392 9772 26444
rect 9824 26432 9830 26444
rect 10781 26435 10839 26441
rect 10781 26432 10793 26435
rect 9824 26404 10793 26432
rect 9824 26392 9830 26404
rect 10781 26401 10793 26404
rect 10827 26401 10839 26435
rect 12621 26435 12679 26441
rect 12621 26432 12633 26435
rect 10781 26395 10839 26401
rect 12406 26404 12633 26432
rect 7147 26336 7236 26364
rect 7331 26367 7389 26373
rect 7147 26333 7159 26336
rect 7101 26327 7159 26333
rect 7331 26333 7343 26367
rect 7377 26364 7389 26367
rect 7466 26364 7472 26376
rect 7377 26336 7472 26364
rect 7377 26333 7389 26336
rect 7331 26327 7389 26333
rect 4709 26299 4767 26305
rect 4709 26296 4721 26299
rect 3896 26268 4721 26296
rect 3789 26259 3847 26265
rect 4709 26265 4721 26268
rect 4755 26296 4767 26299
rect 5626 26296 5632 26308
rect 4755 26268 5632 26296
rect 4755 26265 4767 26268
rect 4709 26259 4767 26265
rect 5626 26256 5632 26268
rect 5684 26296 5690 26308
rect 5684 26268 6132 26296
rect 5684 26256 5690 26268
rect 3142 26228 3148 26240
rect 2976 26200 3148 26228
rect 3142 26188 3148 26200
rect 3200 26228 3206 26240
rect 3602 26228 3608 26240
rect 3200 26200 3608 26228
rect 3200 26188 3206 26200
rect 3602 26188 3608 26200
rect 3660 26188 3666 26240
rect 6104 26228 6132 26268
rect 6178 26256 6184 26308
rect 6236 26296 6242 26308
rect 7024 26296 7052 26327
rect 7466 26324 7472 26336
rect 7524 26324 7530 26376
rect 7926 26324 7932 26376
rect 7984 26364 7990 26376
rect 8021 26367 8079 26373
rect 8021 26364 8033 26367
rect 7984 26336 8033 26364
rect 7984 26324 7990 26336
rect 8021 26333 8033 26336
rect 8067 26333 8079 26367
rect 9398 26364 9404 26376
rect 9359 26336 9404 26364
rect 8021 26327 8079 26333
rect 9398 26324 9404 26336
rect 9456 26324 9462 26376
rect 9582 26364 9588 26376
rect 9543 26336 9588 26364
rect 9582 26324 9588 26336
rect 9640 26324 9646 26376
rect 6236 26268 7052 26296
rect 7193 26299 7251 26305
rect 6236 26256 6242 26268
rect 7193 26265 7205 26299
rect 7239 26296 7251 26299
rect 8110 26296 8116 26308
rect 7239 26268 8116 26296
rect 7239 26265 7251 26268
rect 7193 26259 7251 26265
rect 8110 26256 8116 26268
rect 8168 26256 8174 26308
rect 8202 26256 8208 26308
rect 8260 26296 8266 26308
rect 9784 26296 9812 26392
rect 10318 26324 10324 26376
rect 10376 26364 10382 26376
rect 10597 26367 10655 26373
rect 10597 26364 10609 26367
rect 10376 26336 10609 26364
rect 10376 26324 10382 26336
rect 10597 26333 10609 26336
rect 10643 26364 10655 26367
rect 12406 26364 12434 26404
rect 12621 26401 12633 26404
rect 12667 26401 12679 26435
rect 12621 26395 12679 26401
rect 16758 26392 16764 26444
rect 16816 26432 16822 26444
rect 21284 26441 21312 26472
rect 21269 26435 21327 26441
rect 21269 26432 21281 26435
rect 16816 26404 21281 26432
rect 16816 26392 16822 26404
rect 21269 26401 21281 26404
rect 21315 26401 21327 26435
rect 22204 26432 22232 26472
rect 24302 26460 24308 26472
rect 24360 26500 24366 26512
rect 25038 26500 25044 26512
rect 24360 26472 25044 26500
rect 24360 26460 24366 26472
rect 25038 26460 25044 26472
rect 25096 26460 25102 26512
rect 24486 26432 24492 26444
rect 22204 26404 24492 26432
rect 21269 26395 21327 26401
rect 10643 26336 12434 26364
rect 12897 26367 12955 26373
rect 10643 26333 10655 26336
rect 10597 26327 10655 26333
rect 12897 26333 12909 26367
rect 12943 26333 12955 26367
rect 12897 26327 12955 26333
rect 16393 26367 16451 26373
rect 16393 26333 16405 26367
rect 16439 26364 16451 26367
rect 16574 26364 16580 26376
rect 16439 26336 16580 26364
rect 16439 26333 16451 26336
rect 16393 26327 16451 26333
rect 8260 26268 9812 26296
rect 8260 26256 8266 26268
rect 10870 26256 10876 26308
rect 10928 26296 10934 26308
rect 11333 26299 11391 26305
rect 11333 26296 11345 26299
rect 10928 26268 11345 26296
rect 10928 26256 10934 26268
rect 11333 26265 11345 26268
rect 11379 26265 11391 26299
rect 12912 26296 12940 26327
rect 16574 26324 16580 26336
rect 16632 26364 16638 26376
rect 16853 26367 16911 26373
rect 16853 26364 16865 26367
rect 16632 26336 16865 26364
rect 16632 26324 16638 26336
rect 16853 26333 16865 26336
rect 16899 26333 16911 26367
rect 16853 26327 16911 26333
rect 13449 26299 13507 26305
rect 13449 26296 13461 26299
rect 12912 26268 13461 26296
rect 11333 26259 11391 26265
rect 13449 26265 13461 26268
rect 13495 26296 13507 26299
rect 14090 26296 14096 26308
rect 13495 26268 14096 26296
rect 13495 26265 13507 26268
rect 13449 26259 13507 26265
rect 14090 26256 14096 26268
rect 14148 26256 14154 26308
rect 16868 26296 16896 26327
rect 17034 26324 17040 26376
rect 17092 26364 17098 26376
rect 17770 26364 17776 26376
rect 17092 26336 17776 26364
rect 17092 26324 17098 26336
rect 17770 26324 17776 26336
rect 17828 26324 17834 26376
rect 18049 26367 18107 26373
rect 18049 26333 18061 26367
rect 18095 26333 18107 26367
rect 18230 26364 18236 26376
rect 18191 26336 18236 26364
rect 18049 26327 18107 26333
rect 17310 26296 17316 26308
rect 16868 26268 17316 26296
rect 17310 26256 17316 26268
rect 17368 26256 17374 26308
rect 18064 26296 18092 26327
rect 18230 26324 18236 26336
rect 18288 26324 18294 26376
rect 18325 26367 18383 26373
rect 18325 26333 18337 26367
rect 18371 26333 18383 26367
rect 18325 26327 18383 26333
rect 18417 26367 18475 26373
rect 18417 26333 18429 26367
rect 18463 26364 18475 26367
rect 18690 26364 18696 26376
rect 18463 26336 18696 26364
rect 18463 26333 18475 26336
rect 18417 26327 18475 26333
rect 18138 26296 18144 26308
rect 18064 26268 18144 26296
rect 18138 26256 18144 26268
rect 18196 26256 18202 26308
rect 6270 26228 6276 26240
rect 6104 26200 6276 26228
rect 6270 26188 6276 26200
rect 6328 26188 6334 26240
rect 6365 26231 6423 26237
rect 6365 26197 6377 26231
rect 6411 26228 6423 26231
rect 6546 26228 6552 26240
rect 6411 26200 6552 26228
rect 6411 26197 6423 26200
rect 6365 26191 6423 26197
rect 6546 26188 6552 26200
rect 6604 26188 6610 26240
rect 18046 26188 18052 26240
rect 18104 26228 18110 26240
rect 18340 26228 18368 26327
rect 18690 26324 18696 26336
rect 18748 26364 18754 26376
rect 19337 26367 19395 26373
rect 19337 26364 19349 26367
rect 18748 26336 19349 26364
rect 18748 26324 18754 26336
rect 19337 26333 19349 26336
rect 19383 26364 19395 26367
rect 21818 26364 21824 26376
rect 19383 26336 21726 26364
rect 21779 26336 21824 26364
rect 19383 26333 19395 26336
rect 19337 26327 19395 26333
rect 20806 26296 20812 26308
rect 20767 26268 20812 26296
rect 20806 26256 20812 26268
rect 20864 26256 20870 26308
rect 21698 26296 21726 26336
rect 21818 26324 21824 26336
rect 21876 26324 21882 26376
rect 21981 26364 21987 26376
rect 21942 26336 21987 26364
rect 21981 26324 21987 26336
rect 22039 26324 22045 26376
rect 22094 26324 22100 26376
rect 22152 26364 22158 26376
rect 22250 26373 22278 26404
rect 24486 26392 24492 26404
rect 24544 26392 24550 26444
rect 25148 26432 25176 26540
rect 25314 26528 25320 26540
rect 25372 26528 25378 26580
rect 26418 26568 26424 26580
rect 26379 26540 26424 26568
rect 26418 26528 26424 26540
rect 26476 26528 26482 26580
rect 29454 26528 29460 26580
rect 29512 26568 29518 26580
rect 29638 26568 29644 26580
rect 29512 26540 29644 26568
rect 29512 26528 29518 26540
rect 29638 26528 29644 26540
rect 29696 26528 29702 26580
rect 30098 26568 30104 26580
rect 30059 26540 30104 26568
rect 30098 26528 30104 26540
rect 30156 26568 30162 26580
rect 33962 26568 33968 26580
rect 30156 26540 33968 26568
rect 30156 26528 30162 26540
rect 33962 26528 33968 26540
rect 34020 26528 34026 26580
rect 35434 26568 35440 26580
rect 34716 26540 35440 26568
rect 32214 26500 32220 26512
rect 32175 26472 32220 26500
rect 32214 26460 32220 26472
rect 32272 26500 32278 26512
rect 32766 26500 32772 26512
rect 32272 26472 32772 26500
rect 32272 26460 32278 26472
rect 32766 26460 32772 26472
rect 32824 26460 32830 26512
rect 34716 26509 34744 26540
rect 35434 26528 35440 26540
rect 35492 26528 35498 26580
rect 37936 26540 40080 26568
rect 34701 26503 34759 26509
rect 34701 26500 34713 26503
rect 33060 26472 34713 26500
rect 25148 26404 25820 26432
rect 22235 26367 22293 26373
rect 22152 26336 22197 26364
rect 22152 26324 22158 26336
rect 22235 26333 22247 26367
rect 22281 26333 22293 26367
rect 24670 26364 24676 26376
rect 24631 26336 24676 26364
rect 22235 26327 22293 26333
rect 24670 26324 24676 26336
rect 24728 26324 24734 26376
rect 24854 26364 24860 26376
rect 24815 26336 24860 26364
rect 24854 26324 24860 26336
rect 24912 26324 24918 26376
rect 24952 26367 25010 26373
rect 24952 26364 24964 26367
rect 24951 26333 24964 26364
rect 24998 26333 25010 26367
rect 24951 26327 25010 26333
rect 25087 26367 25145 26373
rect 25087 26333 25099 26367
rect 25133 26364 25145 26367
rect 25682 26364 25688 26376
rect 25133 26336 25688 26364
rect 25133 26333 25145 26336
rect 25087 26327 25145 26333
rect 22462 26296 22468 26308
rect 21698 26268 22468 26296
rect 22462 26256 22468 26268
rect 22520 26256 22526 26308
rect 22094 26228 22100 26240
rect 18104 26200 22100 26228
rect 18104 26188 18110 26200
rect 22094 26188 22100 26200
rect 22152 26188 22158 26240
rect 24762 26188 24768 26240
rect 24820 26228 24826 26240
rect 24951 26228 24979 26327
rect 25682 26324 25688 26336
rect 25740 26324 25746 26376
rect 25792 26373 25820 26404
rect 25884 26404 27292 26432
rect 25777 26367 25835 26373
rect 25777 26333 25789 26367
rect 25823 26333 25835 26367
rect 25884 26364 25912 26404
rect 25940 26367 25998 26373
rect 25940 26364 25952 26367
rect 25884 26336 25952 26364
rect 25777 26327 25835 26333
rect 25940 26333 25952 26336
rect 25986 26333 25998 26367
rect 25940 26327 25998 26333
rect 26053 26367 26111 26373
rect 26053 26333 26065 26367
rect 26099 26333 26111 26367
rect 26053 26327 26111 26333
rect 26191 26367 26249 26373
rect 26191 26333 26203 26367
rect 26237 26364 26249 26367
rect 26970 26364 26976 26376
rect 26237 26336 26976 26364
rect 26237 26333 26249 26336
rect 26191 26327 26249 26333
rect 26068 26228 26096 26327
rect 26970 26324 26976 26336
rect 27028 26324 27034 26376
rect 27264 26373 27292 26404
rect 27249 26367 27307 26373
rect 27249 26333 27261 26367
rect 27295 26333 27307 26367
rect 32950 26364 32956 26376
rect 32911 26336 32956 26364
rect 27249 26327 27307 26333
rect 32950 26324 32956 26336
rect 33008 26324 33014 26376
rect 33060 26373 33088 26472
rect 34701 26469 34713 26472
rect 34747 26469 34759 26503
rect 34701 26463 34759 26469
rect 36906 26460 36912 26512
rect 36964 26500 36970 26512
rect 37936 26509 37964 26540
rect 37921 26503 37979 26509
rect 37921 26500 37933 26503
rect 36964 26472 37933 26500
rect 36964 26460 36970 26472
rect 37921 26469 37933 26472
rect 37967 26469 37979 26503
rect 37921 26463 37979 26469
rect 33778 26432 33784 26444
rect 33152 26404 33784 26432
rect 33152 26373 33180 26404
rect 33778 26392 33784 26404
rect 33836 26392 33842 26444
rect 33870 26392 33876 26444
rect 33928 26432 33934 26444
rect 34422 26432 34428 26444
rect 33928 26404 34428 26432
rect 33928 26392 33934 26404
rect 34422 26392 34428 26404
rect 34480 26392 34486 26444
rect 33045 26367 33103 26373
rect 33045 26333 33057 26367
rect 33091 26333 33103 26367
rect 33045 26327 33103 26333
rect 33137 26367 33195 26373
rect 33137 26333 33149 26367
rect 33183 26333 33195 26367
rect 33318 26364 33324 26376
rect 33279 26336 33324 26364
rect 33137 26327 33195 26333
rect 33318 26324 33324 26336
rect 33376 26324 33382 26376
rect 34514 26324 34520 26376
rect 34572 26364 34578 26376
rect 35814 26367 35872 26373
rect 35814 26364 35826 26367
rect 34572 26336 35826 26364
rect 34572 26324 34578 26336
rect 35814 26333 35826 26336
rect 35860 26333 35872 26367
rect 35814 26327 35872 26333
rect 36081 26367 36139 26373
rect 36081 26333 36093 26367
rect 36127 26364 36139 26367
rect 37090 26364 37096 26376
rect 36127 26336 37096 26364
rect 36127 26333 36139 26336
rect 36081 26327 36139 26333
rect 37090 26324 37096 26336
rect 37148 26364 37154 26376
rect 38746 26364 38752 26376
rect 37148 26336 38752 26364
rect 37148 26324 37154 26336
rect 38746 26324 38752 26336
rect 38804 26364 38810 26376
rect 39301 26367 39359 26373
rect 39301 26364 39313 26367
rect 38804 26336 39313 26364
rect 38804 26324 38810 26336
rect 39301 26333 39313 26336
rect 39347 26364 39359 26367
rect 39942 26364 39948 26376
rect 39347 26336 39948 26364
rect 39347 26333 39359 26336
rect 39301 26327 39359 26333
rect 39942 26324 39948 26336
rect 40000 26324 40006 26376
rect 40052 26373 40080 26540
rect 40037 26367 40095 26373
rect 40037 26333 40049 26367
rect 40083 26333 40095 26367
rect 40037 26327 40095 26333
rect 26326 26256 26332 26308
rect 26384 26296 26390 26308
rect 26881 26299 26939 26305
rect 26881 26296 26893 26299
rect 26384 26268 26893 26296
rect 26384 26256 26390 26268
rect 26881 26265 26893 26268
rect 26927 26265 26939 26299
rect 26881 26259 26939 26265
rect 27065 26299 27123 26305
rect 27065 26265 27077 26299
rect 27111 26296 27123 26299
rect 29270 26296 29276 26308
rect 27111 26268 29276 26296
rect 27111 26265 27123 26268
rect 27065 26259 27123 26265
rect 29270 26256 29276 26268
rect 29328 26256 29334 26308
rect 39056 26299 39114 26305
rect 39056 26265 39068 26299
rect 39102 26296 39114 26299
rect 39758 26296 39764 26308
rect 39102 26268 39764 26296
rect 39102 26265 39114 26268
rect 39056 26259 39114 26265
rect 39758 26256 39764 26268
rect 39816 26256 39822 26308
rect 39850 26256 39856 26308
rect 39908 26296 39914 26308
rect 39908 26268 39953 26296
rect 39908 26256 39914 26268
rect 32766 26228 32772 26240
rect 24820 26200 26096 26228
rect 32727 26200 32772 26228
rect 24820 26188 24826 26200
rect 32766 26188 32772 26200
rect 32824 26188 32830 26240
rect 40221 26231 40279 26237
rect 40221 26197 40233 26231
rect 40267 26228 40279 26231
rect 40402 26228 40408 26240
rect 40267 26200 40408 26228
rect 40267 26197 40279 26200
rect 40221 26191 40279 26197
rect 40402 26188 40408 26200
rect 40460 26188 40466 26240
rect 40770 26228 40776 26240
rect 40731 26200 40776 26228
rect 40770 26188 40776 26200
rect 40828 26188 40834 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 3970 26024 3976 26036
rect 3931 25996 3976 26024
rect 3970 25984 3976 25996
rect 4028 25984 4034 26036
rect 6362 25984 6368 26036
rect 6420 26024 6426 26036
rect 7561 26027 7619 26033
rect 7561 26024 7573 26027
rect 6420 25996 7573 26024
rect 6420 25984 6426 25996
rect 7561 25993 7573 25996
rect 7607 26024 7619 26027
rect 8202 26024 8208 26036
rect 7607 25996 8208 26024
rect 7607 25993 7619 25996
rect 7561 25987 7619 25993
rect 8202 25984 8208 25996
rect 8260 25984 8266 26036
rect 9030 26024 9036 26036
rect 8943 25996 9036 26024
rect 9030 25984 9036 25996
rect 9088 26024 9094 26036
rect 10594 26024 10600 26036
rect 9088 25996 10600 26024
rect 9088 25984 9094 25996
rect 10594 25984 10600 25996
rect 10652 25984 10658 26036
rect 13446 25984 13452 26036
rect 13504 26024 13510 26036
rect 13541 26027 13599 26033
rect 13541 26024 13553 26027
rect 13504 25996 13553 26024
rect 13504 25984 13510 25996
rect 13541 25993 13553 25996
rect 13587 25993 13599 26027
rect 17678 26024 17684 26036
rect 17639 25996 17684 26024
rect 13541 25987 13599 25993
rect 17678 25984 17684 25996
rect 17736 25984 17742 26036
rect 18230 25984 18236 26036
rect 18288 26024 18294 26036
rect 18785 26027 18843 26033
rect 18785 26024 18797 26027
rect 18288 25996 18797 26024
rect 18288 25984 18294 25996
rect 18785 25993 18797 25996
rect 18831 25993 18843 26027
rect 21818 26024 21824 26036
rect 18785 25987 18843 25993
rect 18892 25996 21824 26024
rect 2866 25965 2872 25968
rect 2860 25919 2872 25965
rect 2924 25956 2930 25968
rect 2924 25928 2960 25956
rect 2866 25916 2872 25919
rect 2924 25916 2930 25928
rect 6086 25916 6092 25968
rect 6144 25956 6150 25968
rect 8021 25959 8079 25965
rect 8021 25956 8033 25959
rect 6144 25928 8033 25956
rect 6144 25916 6150 25928
rect 6748 25900 6776 25928
rect 8021 25925 8033 25928
rect 8067 25925 8079 25959
rect 8021 25919 8079 25925
rect 10318 25916 10324 25968
rect 10376 25956 10382 25968
rect 10689 25959 10747 25965
rect 10689 25956 10701 25959
rect 10376 25928 10701 25956
rect 10376 25916 10382 25928
rect 10689 25925 10701 25928
rect 10735 25925 10747 25959
rect 18414 25956 18420 25968
rect 10689 25919 10747 25925
rect 17926 25928 18420 25956
rect 6362 25888 6368 25900
rect 6323 25860 6368 25888
rect 6362 25848 6368 25860
rect 6420 25848 6426 25900
rect 6546 25888 6552 25900
rect 6507 25860 6552 25888
rect 6546 25848 6552 25860
rect 6604 25848 6610 25900
rect 6641 25891 6699 25897
rect 6641 25857 6653 25891
rect 6687 25857 6699 25891
rect 6641 25851 6699 25857
rect 2406 25780 2412 25832
rect 2464 25820 2470 25832
rect 2593 25823 2651 25829
rect 2593 25820 2605 25823
rect 2464 25792 2605 25820
rect 2464 25780 2470 25792
rect 2593 25789 2605 25792
rect 2639 25789 2651 25823
rect 2593 25783 2651 25789
rect 3602 25780 3608 25832
rect 3660 25820 3666 25832
rect 6656 25820 6684 25851
rect 6730 25848 6736 25900
rect 6788 25888 6794 25900
rect 6788 25860 6881 25888
rect 6788 25848 6794 25860
rect 12802 25848 12808 25900
rect 12860 25888 12866 25900
rect 13633 25891 13691 25897
rect 13633 25888 13645 25891
rect 12860 25860 13645 25888
rect 12860 25848 12866 25860
rect 13633 25857 13645 25860
rect 13679 25857 13691 25891
rect 13633 25851 13691 25857
rect 14090 25848 14096 25900
rect 14148 25888 14154 25900
rect 14277 25891 14335 25897
rect 14277 25888 14289 25891
rect 14148 25860 14289 25888
rect 14148 25848 14154 25860
rect 14277 25857 14289 25860
rect 14323 25857 14335 25891
rect 15746 25888 15752 25900
rect 15707 25860 15752 25888
rect 14277 25851 14335 25857
rect 15746 25848 15752 25860
rect 15804 25848 15810 25900
rect 16853 25891 16911 25897
rect 16853 25857 16865 25891
rect 16899 25888 16911 25891
rect 17494 25888 17500 25900
rect 16899 25860 17500 25888
rect 16899 25857 16911 25860
rect 16853 25851 16911 25857
rect 17494 25848 17500 25860
rect 17552 25848 17558 25900
rect 17926 25897 17954 25928
rect 18414 25916 18420 25928
rect 18472 25956 18478 25968
rect 18598 25956 18604 25968
rect 18472 25928 18604 25956
rect 18472 25916 18478 25928
rect 18598 25916 18604 25928
rect 18656 25916 18662 25968
rect 17911 25891 17969 25897
rect 17911 25857 17923 25891
rect 17957 25857 17969 25891
rect 18046 25888 18052 25900
rect 18007 25860 18052 25888
rect 17911 25851 17969 25857
rect 18046 25848 18052 25860
rect 18104 25848 18110 25900
rect 18162 25891 18220 25897
rect 18162 25857 18174 25891
rect 18208 25888 18220 25891
rect 18325 25891 18383 25897
rect 18208 25860 18276 25888
rect 18208 25857 18220 25860
rect 18162 25851 18220 25857
rect 7834 25820 7840 25832
rect 3660 25792 7840 25820
rect 3660 25780 3666 25792
rect 7834 25780 7840 25792
rect 7892 25780 7898 25832
rect 9398 25780 9404 25832
rect 9456 25820 9462 25832
rect 9769 25823 9827 25829
rect 9769 25820 9781 25823
rect 9456 25792 9781 25820
rect 9456 25780 9462 25792
rect 9769 25789 9781 25792
rect 9815 25820 9827 25823
rect 13814 25820 13820 25832
rect 9815 25792 13820 25820
rect 9815 25789 9827 25792
rect 9769 25783 9827 25789
rect 13814 25780 13820 25792
rect 13872 25780 13878 25832
rect 13906 25780 13912 25832
rect 13964 25820 13970 25832
rect 15473 25823 15531 25829
rect 15473 25820 15485 25823
rect 13964 25792 15485 25820
rect 13964 25780 13970 25792
rect 15473 25789 15485 25792
rect 15519 25789 15531 25823
rect 18248 25820 18276 25860
rect 18325 25857 18337 25891
rect 18371 25888 18383 25891
rect 18892 25888 18920 25996
rect 21818 25984 21824 25996
rect 21876 25984 21882 26036
rect 25222 25984 25228 26036
rect 25280 26024 25286 26036
rect 25777 26027 25835 26033
rect 25777 26024 25789 26027
rect 25280 25996 25789 26024
rect 25280 25984 25286 25996
rect 25777 25993 25789 25996
rect 25823 25993 25835 26027
rect 26970 26024 26976 26036
rect 25777 25987 25835 25993
rect 25875 25996 26976 26024
rect 18969 25959 19027 25965
rect 18969 25925 18981 25959
rect 19015 25956 19027 25959
rect 20438 25956 20444 25968
rect 19015 25928 20444 25956
rect 19015 25925 19027 25928
rect 18969 25919 19027 25925
rect 20438 25916 20444 25928
rect 20496 25916 20502 25968
rect 21269 25959 21327 25965
rect 21269 25925 21281 25959
rect 21315 25956 21327 25959
rect 21315 25928 21956 25956
rect 21315 25925 21327 25928
rect 21269 25919 21327 25925
rect 18371 25860 18920 25888
rect 19153 25891 19211 25897
rect 18371 25857 18383 25860
rect 18325 25851 18383 25857
rect 19153 25857 19165 25891
rect 19199 25888 19211 25891
rect 19242 25888 19248 25900
rect 19199 25860 19248 25888
rect 19199 25857 19211 25860
rect 19153 25851 19211 25857
rect 19242 25848 19248 25860
rect 19300 25848 19306 25900
rect 19426 25848 19432 25900
rect 19484 25888 19490 25900
rect 19797 25891 19855 25897
rect 19797 25888 19809 25891
rect 19484 25860 19809 25888
rect 19484 25848 19490 25860
rect 19797 25857 19809 25860
rect 19843 25857 19855 25891
rect 19981 25891 20039 25897
rect 19981 25888 19993 25891
rect 19797 25851 19855 25857
rect 19904 25860 19993 25888
rect 19613 25823 19671 25829
rect 19613 25820 19625 25823
rect 18248 25792 19625 25820
rect 15473 25783 15531 25789
rect 19613 25789 19625 25792
rect 19659 25789 19671 25823
rect 19613 25783 19671 25789
rect 11330 25712 11336 25764
rect 11388 25752 11394 25764
rect 14461 25755 14519 25761
rect 14461 25752 14473 25755
rect 11388 25724 14473 25752
rect 11388 25712 11394 25724
rect 14461 25721 14473 25724
rect 14507 25752 14519 25755
rect 16022 25752 16028 25764
rect 14507 25724 16028 25752
rect 14507 25721 14519 25724
rect 14461 25715 14519 25721
rect 16022 25712 16028 25724
rect 16080 25712 16086 25764
rect 19242 25712 19248 25764
rect 19300 25752 19306 25764
rect 19904 25752 19932 25860
rect 19981 25857 19993 25860
rect 20027 25888 20039 25891
rect 20898 25888 20904 25900
rect 20027 25860 20904 25888
rect 20027 25857 20039 25860
rect 19981 25851 20039 25857
rect 20898 25848 20904 25860
rect 20956 25848 20962 25900
rect 21085 25891 21143 25897
rect 21085 25857 21097 25891
rect 21131 25888 21143 25891
rect 21634 25888 21640 25900
rect 21131 25860 21640 25888
rect 21131 25857 21143 25860
rect 21085 25851 21143 25857
rect 21634 25848 21640 25860
rect 21692 25848 21698 25900
rect 21818 25888 21824 25900
rect 21779 25860 21824 25888
rect 21818 25848 21824 25860
rect 21876 25848 21882 25900
rect 21928 25888 21956 25928
rect 22462 25916 22468 25968
rect 22520 25956 22526 25968
rect 25317 25959 25375 25965
rect 25317 25956 25329 25959
rect 22520 25928 25329 25956
rect 22520 25916 22526 25928
rect 25317 25925 25329 25928
rect 25363 25956 25375 25959
rect 25682 25956 25688 25968
rect 25363 25928 25688 25956
rect 25363 25925 25375 25928
rect 25317 25919 25375 25925
rect 25682 25916 25688 25928
rect 25740 25916 25746 25968
rect 21984 25891 22042 25897
rect 21984 25888 21996 25891
rect 21928 25860 21996 25888
rect 21984 25857 21996 25860
rect 22030 25857 22042 25891
rect 21984 25851 22042 25857
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 22235 25891 22293 25897
rect 22152 25860 22197 25888
rect 22152 25848 22158 25860
rect 22235 25857 22247 25891
rect 22281 25888 22293 25891
rect 23017 25891 23075 25897
rect 23017 25888 23029 25891
rect 22281 25860 23029 25888
rect 22281 25857 22293 25860
rect 22235 25851 22293 25857
rect 23017 25857 23029 25860
rect 23063 25888 23075 25891
rect 25875 25888 25903 25996
rect 26970 25984 26976 25996
rect 27028 25984 27034 26036
rect 30098 25984 30104 26036
rect 30156 25984 30162 26036
rect 31570 25984 31576 26036
rect 31628 26024 31634 26036
rect 32766 26024 32772 26036
rect 31628 25996 32772 26024
rect 31628 25984 31634 25996
rect 32766 25984 32772 25996
rect 32824 25984 32830 26036
rect 33686 25984 33692 26036
rect 33744 26024 33750 26036
rect 34333 26027 34391 26033
rect 34333 26024 34345 26027
rect 33744 25996 34345 26024
rect 33744 25984 33750 25996
rect 34333 25993 34345 25996
rect 34379 25993 34391 26027
rect 34333 25987 34391 25993
rect 26145 25959 26203 25965
rect 26145 25925 26157 25959
rect 26191 25956 26203 25959
rect 26326 25956 26332 25968
rect 26191 25928 26332 25956
rect 26191 25925 26203 25928
rect 26145 25919 26203 25925
rect 26326 25916 26332 25928
rect 26384 25916 26390 25968
rect 27709 25959 27767 25965
rect 27709 25925 27721 25959
rect 27755 25956 27767 25959
rect 30116 25956 30144 25984
rect 33226 25965 33232 25968
rect 33220 25956 33232 25965
rect 27755 25928 30144 25956
rect 33187 25928 33232 25956
rect 27755 25925 27767 25928
rect 27709 25919 27767 25925
rect 33220 25919 33232 25928
rect 33226 25916 33232 25919
rect 33284 25916 33290 25968
rect 39700 25959 39758 25965
rect 39700 25925 39712 25959
rect 39746 25956 39758 25959
rect 41049 25959 41107 25965
rect 41049 25956 41061 25959
rect 39746 25928 41061 25956
rect 39746 25925 39758 25928
rect 39700 25919 39758 25925
rect 41049 25925 41061 25928
rect 41095 25925 41107 25959
rect 41049 25919 41107 25925
rect 23063 25860 25903 25888
rect 25961 25891 26019 25897
rect 23063 25857 23075 25860
rect 23017 25851 23075 25857
rect 25961 25857 25973 25891
rect 26007 25888 26019 25891
rect 28534 25888 28540 25900
rect 26007 25860 28540 25888
rect 26007 25857 26019 25860
rect 25961 25851 26019 25857
rect 28534 25848 28540 25860
rect 28592 25848 28598 25900
rect 28626 25848 28632 25900
rect 28684 25888 28690 25900
rect 29917 25891 29975 25897
rect 29917 25888 29929 25891
rect 28684 25860 29929 25888
rect 28684 25848 28690 25860
rect 29917 25857 29929 25860
rect 29963 25857 29975 25891
rect 29917 25851 29975 25857
rect 30101 25891 30159 25897
rect 30101 25857 30113 25891
rect 30147 25857 30159 25891
rect 30101 25851 30159 25857
rect 40405 25891 40463 25897
rect 40405 25857 40417 25891
rect 40451 25857 40463 25891
rect 40586 25888 40592 25900
rect 40547 25860 40592 25888
rect 40405 25851 40463 25857
rect 24118 25780 24124 25832
rect 24176 25820 24182 25832
rect 30116 25820 30144 25851
rect 31294 25820 31300 25832
rect 24176 25792 31300 25820
rect 24176 25780 24182 25792
rect 31294 25780 31300 25792
rect 31352 25780 31358 25832
rect 32953 25823 33011 25829
rect 32953 25789 32965 25823
rect 32999 25789 33011 25823
rect 39942 25820 39948 25832
rect 39903 25792 39948 25820
rect 32953 25783 33011 25789
rect 19300 25724 19932 25752
rect 19300 25712 19306 25724
rect 25498 25712 25504 25764
rect 25556 25752 25562 25764
rect 31202 25752 31208 25764
rect 25556 25724 31208 25752
rect 25556 25712 25562 25724
rect 31202 25712 31208 25724
rect 31260 25712 31266 25764
rect 7006 25684 7012 25696
rect 6967 25656 7012 25684
rect 7006 25644 7012 25656
rect 7064 25644 7070 25696
rect 12802 25644 12808 25696
rect 12860 25684 12866 25696
rect 12897 25687 12955 25693
rect 12897 25684 12909 25687
rect 12860 25656 12909 25684
rect 12860 25644 12866 25656
rect 12897 25653 12909 25656
rect 12943 25653 12955 25687
rect 12897 25647 12955 25653
rect 15562 25644 15568 25696
rect 15620 25684 15626 25696
rect 16669 25687 16727 25693
rect 16669 25684 16681 25687
rect 15620 25656 16681 25684
rect 15620 25644 15626 25656
rect 16669 25653 16681 25656
rect 16715 25653 16727 25687
rect 22462 25684 22468 25696
rect 22423 25656 22468 25684
rect 16669 25647 16727 25653
rect 22462 25644 22468 25656
rect 22520 25644 22526 25696
rect 27614 25644 27620 25696
rect 27672 25684 27678 25696
rect 28997 25687 29055 25693
rect 28997 25684 29009 25687
rect 27672 25656 29009 25684
rect 27672 25644 27678 25656
rect 28997 25653 29009 25656
rect 29043 25653 29055 25687
rect 28997 25647 29055 25653
rect 30285 25687 30343 25693
rect 30285 25653 30297 25687
rect 30331 25684 30343 25687
rect 30742 25684 30748 25696
rect 30331 25656 30748 25684
rect 30331 25653 30343 25656
rect 30285 25647 30343 25653
rect 30742 25644 30748 25656
rect 30800 25644 30806 25696
rect 32968 25684 32996 25783
rect 39942 25780 39948 25792
rect 40000 25780 40006 25832
rect 40420 25820 40448 25851
rect 40586 25848 40592 25860
rect 40644 25848 40650 25900
rect 40681 25891 40739 25897
rect 40681 25857 40693 25891
rect 40727 25857 40739 25891
rect 40681 25851 40739 25857
rect 40494 25820 40500 25832
rect 40420 25792 40500 25820
rect 40494 25780 40500 25792
rect 40552 25780 40558 25832
rect 37274 25712 37280 25764
rect 37332 25752 37338 25764
rect 38562 25752 38568 25764
rect 37332 25724 38568 25752
rect 37332 25712 37338 25724
rect 38562 25712 38568 25724
rect 38620 25712 38626 25764
rect 40218 25712 40224 25764
rect 40276 25752 40282 25764
rect 40696 25752 40724 25851
rect 40770 25848 40776 25900
rect 40828 25888 40834 25900
rect 40828 25860 40873 25888
rect 40828 25848 40834 25860
rect 40276 25724 40724 25752
rect 40276 25712 40282 25724
rect 33134 25684 33140 25696
rect 32968 25656 33140 25684
rect 33134 25644 33140 25656
rect 33192 25644 33198 25696
rect 36354 25644 36360 25696
rect 36412 25684 36418 25696
rect 37366 25684 37372 25696
rect 36412 25656 37372 25684
rect 36412 25644 36418 25656
rect 37366 25644 37372 25656
rect 37424 25644 37430 25696
rect 39298 25644 39304 25696
rect 39356 25684 39362 25696
rect 40586 25684 40592 25696
rect 39356 25656 40592 25684
rect 39356 25644 39362 25656
rect 40586 25644 40592 25656
rect 40644 25644 40650 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 6178 25440 6184 25492
rect 6236 25480 6242 25492
rect 7745 25483 7803 25489
rect 7745 25480 7757 25483
rect 6236 25452 7757 25480
rect 6236 25440 6242 25452
rect 7745 25449 7757 25452
rect 7791 25449 7803 25483
rect 7745 25443 7803 25449
rect 8389 25483 8447 25489
rect 8389 25449 8401 25483
rect 8435 25480 8447 25483
rect 8570 25480 8576 25492
rect 8435 25452 8576 25480
rect 8435 25449 8447 25452
rect 8389 25443 8447 25449
rect 8570 25440 8576 25452
rect 8628 25440 8634 25492
rect 18046 25440 18052 25492
rect 18104 25480 18110 25492
rect 18104 25452 18368 25480
rect 18104 25440 18110 25452
rect 17954 25412 17960 25424
rect 9508 25384 17960 25412
rect 2406 25236 2412 25288
rect 2464 25276 2470 25288
rect 4341 25279 4399 25285
rect 4341 25276 4353 25279
rect 2464 25248 4353 25276
rect 2464 25236 2470 25248
rect 4341 25245 4353 25248
rect 4387 25276 4399 25279
rect 6362 25276 6368 25288
rect 4387 25248 6368 25276
rect 4387 25245 4399 25248
rect 4341 25239 4399 25245
rect 6362 25236 6368 25248
rect 6420 25236 6426 25288
rect 6632 25279 6690 25285
rect 6632 25245 6644 25279
rect 6678 25276 6690 25279
rect 7006 25276 7012 25288
rect 6678 25248 7012 25276
rect 6678 25245 6690 25248
rect 6632 25239 6690 25245
rect 7006 25236 7012 25248
rect 7064 25236 7070 25288
rect 8570 25236 8576 25288
rect 8628 25276 8634 25288
rect 9508 25285 9536 25384
rect 17954 25372 17960 25384
rect 18012 25372 18018 25424
rect 18230 25372 18236 25424
rect 18288 25372 18294 25424
rect 9950 25344 9956 25356
rect 9600 25316 9956 25344
rect 9600 25285 9628 25316
rect 9950 25304 9956 25316
rect 10008 25304 10014 25356
rect 10318 25304 10324 25356
rect 10376 25304 10382 25356
rect 11054 25304 11060 25356
rect 11112 25344 11118 25356
rect 12069 25347 12127 25353
rect 12069 25344 12081 25347
rect 11112 25316 12081 25344
rect 11112 25304 11118 25316
rect 12069 25313 12081 25316
rect 12115 25344 12127 25347
rect 12158 25344 12164 25356
rect 12115 25316 12164 25344
rect 12115 25313 12127 25316
rect 12069 25307 12127 25313
rect 12158 25304 12164 25316
rect 12216 25304 12222 25356
rect 9493 25279 9551 25285
rect 9493 25276 9505 25279
rect 8628 25248 9505 25276
rect 8628 25236 8634 25248
rect 9493 25245 9505 25248
rect 9539 25245 9551 25279
rect 9493 25239 9551 25245
rect 9585 25279 9643 25285
rect 9585 25245 9597 25279
rect 9631 25245 9643 25279
rect 9585 25239 9643 25245
rect 9677 25279 9735 25285
rect 9677 25245 9689 25279
rect 9723 25276 9735 25279
rect 9766 25276 9772 25288
rect 9723 25248 9772 25276
rect 9723 25245 9735 25248
rect 9677 25239 9735 25245
rect 9766 25236 9772 25248
rect 9824 25236 9830 25288
rect 9858 25236 9864 25288
rect 9916 25276 9922 25288
rect 10336 25276 10364 25304
rect 12529 25279 12587 25285
rect 12529 25276 12541 25279
rect 9916 25248 10364 25276
rect 12406 25248 12541 25276
rect 9916 25236 9922 25248
rect 5902 25208 5908 25220
rect 5863 25180 5908 25208
rect 5902 25168 5908 25180
rect 5960 25168 5966 25220
rect 7282 25168 7288 25220
rect 7340 25208 7346 25220
rect 10321 25211 10379 25217
rect 10321 25208 10333 25211
rect 7340 25180 10333 25208
rect 7340 25168 7346 25180
rect 10321 25177 10333 25180
rect 10367 25208 10379 25211
rect 12406 25208 12434 25248
rect 12529 25245 12541 25248
rect 12575 25245 12587 25279
rect 12529 25239 12587 25245
rect 13354 25236 13360 25288
rect 13412 25276 13418 25288
rect 13541 25279 13599 25285
rect 13541 25276 13553 25279
rect 13412 25248 13553 25276
rect 13412 25236 13418 25248
rect 13541 25245 13553 25248
rect 13587 25276 13599 25279
rect 15930 25276 15936 25288
rect 13587 25248 15936 25276
rect 13587 25245 13599 25248
rect 13541 25239 13599 25245
rect 15930 25236 15936 25248
rect 15988 25236 15994 25288
rect 18049 25279 18107 25285
rect 16776 25248 18000 25276
rect 10367 25180 12434 25208
rect 15105 25211 15163 25217
rect 10367 25177 10379 25180
rect 10321 25171 10379 25177
rect 15105 25177 15117 25211
rect 15151 25177 15163 25211
rect 15105 25171 15163 25177
rect 15289 25211 15347 25217
rect 15289 25177 15301 25211
rect 15335 25208 15347 25211
rect 15562 25208 15568 25220
rect 15335 25180 15568 25208
rect 15335 25177 15347 25180
rect 15289 25171 15347 25177
rect 8570 25100 8576 25152
rect 8628 25140 8634 25152
rect 9217 25143 9275 25149
rect 9217 25140 9229 25143
rect 8628 25112 9229 25140
rect 8628 25100 8634 25112
rect 9217 25109 9229 25112
rect 9263 25109 9275 25143
rect 14090 25140 14096 25152
rect 14051 25112 14096 25140
rect 9217 25103 9275 25109
rect 14090 25100 14096 25112
rect 14148 25100 14154 25152
rect 14826 25100 14832 25152
rect 14884 25140 14890 25152
rect 14921 25143 14979 25149
rect 14921 25140 14933 25143
rect 14884 25112 14933 25140
rect 14884 25100 14890 25112
rect 14921 25109 14933 25112
rect 14967 25109 14979 25143
rect 15120 25140 15148 25171
rect 15562 25168 15568 25180
rect 15620 25168 15626 25220
rect 16022 25168 16028 25220
rect 16080 25208 16086 25220
rect 16776 25217 16804 25248
rect 16209 25211 16267 25217
rect 16209 25208 16221 25211
rect 16080 25180 16221 25208
rect 16080 25168 16086 25180
rect 16209 25177 16221 25180
rect 16255 25208 16267 25211
rect 16761 25211 16819 25217
rect 16761 25208 16773 25211
rect 16255 25180 16773 25208
rect 16255 25177 16267 25180
rect 16209 25171 16267 25177
rect 16761 25177 16773 25180
rect 16807 25177 16819 25211
rect 16942 25208 16948 25220
rect 16903 25180 16948 25208
rect 16761 25171 16819 25177
rect 16942 25168 16948 25180
rect 17000 25168 17006 25220
rect 17972 25208 18000 25248
rect 18049 25245 18061 25279
rect 18095 25276 18107 25279
rect 18138 25276 18144 25288
rect 18095 25248 18144 25276
rect 18095 25245 18107 25248
rect 18049 25239 18107 25245
rect 18138 25236 18144 25248
rect 18196 25236 18202 25288
rect 18248 25285 18276 25372
rect 18340 25285 18368 25452
rect 24854 25440 24860 25492
rect 24912 25480 24918 25492
rect 25593 25483 25651 25489
rect 25593 25480 25605 25483
rect 24912 25452 25605 25480
rect 24912 25440 24918 25452
rect 25593 25449 25605 25452
rect 25639 25449 25651 25483
rect 31294 25480 31300 25492
rect 31255 25452 31300 25480
rect 25593 25443 25651 25449
rect 31294 25440 31300 25452
rect 31352 25440 31358 25492
rect 39298 25480 39304 25492
rect 39259 25452 39304 25480
rect 39298 25440 39304 25452
rect 39356 25440 39362 25492
rect 39758 25440 39764 25492
rect 39816 25480 39822 25492
rect 39853 25483 39911 25489
rect 39853 25480 39865 25483
rect 39816 25452 39865 25480
rect 39816 25440 39822 25452
rect 39853 25449 39865 25452
rect 39899 25449 39911 25483
rect 40218 25480 40224 25492
rect 39853 25443 39911 25449
rect 39960 25452 40224 25480
rect 29822 25372 29828 25424
rect 29880 25412 29886 25424
rect 30374 25412 30380 25424
rect 29880 25384 30380 25412
rect 29880 25372 29886 25384
rect 30374 25372 30380 25384
rect 30432 25412 30438 25424
rect 30432 25384 30788 25412
rect 30432 25372 30438 25384
rect 18233 25279 18291 25285
rect 18233 25245 18245 25279
rect 18279 25245 18291 25279
rect 18233 25239 18291 25245
rect 18325 25279 18383 25285
rect 18325 25245 18337 25279
rect 18371 25245 18383 25279
rect 18325 25239 18383 25245
rect 18463 25279 18521 25285
rect 18463 25245 18475 25279
rect 18509 25276 18521 25279
rect 19334 25276 19340 25288
rect 18509 25248 19340 25276
rect 18509 25245 18521 25248
rect 18463 25239 18521 25245
rect 19334 25236 19340 25248
rect 19392 25236 19398 25288
rect 21726 25236 21732 25288
rect 21784 25276 21790 25288
rect 23017 25279 23075 25285
rect 23017 25276 23029 25279
rect 21784 25248 23029 25276
rect 21784 25236 21790 25248
rect 23017 25245 23029 25248
rect 23063 25245 23075 25279
rect 23017 25239 23075 25245
rect 24946 25236 24952 25288
rect 25004 25276 25010 25288
rect 25961 25279 26019 25285
rect 25961 25276 25973 25279
rect 25004 25248 25973 25276
rect 25004 25236 25010 25248
rect 25961 25245 25973 25248
rect 26007 25276 26019 25279
rect 26326 25276 26332 25288
rect 26007 25248 26332 25276
rect 26007 25245 26019 25248
rect 25961 25239 26019 25245
rect 26326 25236 26332 25248
rect 26384 25236 26390 25288
rect 29822 25276 29828 25288
rect 29783 25248 29828 25276
rect 29822 25236 29828 25248
rect 29880 25236 29886 25288
rect 29914 25276 29972 25282
rect 30193 25279 30251 25285
rect 29914 25242 29926 25276
rect 29960 25242 29972 25276
rect 29914 25236 29972 25242
rect 30009 25273 30067 25279
rect 30009 25239 30021 25273
rect 30055 25239 30067 25273
rect 30193 25245 30205 25279
rect 30239 25276 30251 25279
rect 30650 25276 30656 25288
rect 30239 25248 30656 25276
rect 30239 25245 30251 25248
rect 30193 25239 30251 25245
rect 20162 25208 20168 25220
rect 17972 25180 20168 25208
rect 20162 25168 20168 25180
rect 20220 25168 20226 25220
rect 22462 25168 22468 25220
rect 22520 25208 22526 25220
rect 22750 25211 22808 25217
rect 22750 25208 22762 25211
rect 22520 25180 22762 25208
rect 22520 25168 22526 25180
rect 22750 25177 22762 25180
rect 22796 25177 22808 25211
rect 22750 25171 22808 25177
rect 25777 25211 25835 25217
rect 25777 25177 25789 25211
rect 25823 25208 25835 25211
rect 26234 25208 26240 25220
rect 25823 25180 26240 25208
rect 25823 25177 25835 25180
rect 25777 25171 25835 25177
rect 26234 25168 26240 25180
rect 26292 25168 26298 25220
rect 29730 25168 29736 25220
rect 29788 25208 29794 25220
rect 29929 25208 29957 25236
rect 30009 25233 30067 25239
rect 30650 25236 30656 25248
rect 30708 25236 30714 25288
rect 29788 25180 29957 25208
rect 29788 25168 29794 25180
rect 30024 25152 30052 25233
rect 15838 25140 15844 25152
rect 15120 25112 15844 25140
rect 14921 25103 14979 25109
rect 15838 25100 15844 25112
rect 15896 25100 15902 25152
rect 17589 25143 17647 25149
rect 17589 25109 17601 25143
rect 17635 25140 17647 25143
rect 18598 25140 18604 25152
rect 17635 25112 18604 25140
rect 17635 25109 17647 25112
rect 17589 25103 17647 25109
rect 18598 25100 18604 25112
rect 18656 25100 18662 25152
rect 18693 25143 18751 25149
rect 18693 25109 18705 25143
rect 18739 25140 18751 25143
rect 19150 25140 19156 25152
rect 18739 25112 19156 25140
rect 18739 25109 18751 25112
rect 18693 25103 18751 25109
rect 19150 25100 19156 25112
rect 19208 25100 19214 25152
rect 19334 25100 19340 25152
rect 19392 25140 19398 25152
rect 20438 25140 20444 25152
rect 19392 25112 20444 25140
rect 19392 25100 19398 25112
rect 20438 25100 20444 25112
rect 20496 25100 20502 25152
rect 21634 25140 21640 25152
rect 21547 25112 21640 25140
rect 21634 25100 21640 25112
rect 21692 25140 21698 25152
rect 22830 25140 22836 25152
rect 21692 25112 22836 25140
rect 21692 25100 21698 25112
rect 22830 25100 22836 25112
rect 22888 25100 22894 25152
rect 28258 25100 28264 25152
rect 28316 25140 28322 25152
rect 28905 25143 28963 25149
rect 28905 25140 28917 25143
rect 28316 25112 28917 25140
rect 28316 25100 28322 25112
rect 28905 25109 28917 25112
rect 28951 25109 28963 25143
rect 28905 25103 28963 25109
rect 29549 25143 29607 25149
rect 29549 25109 29561 25143
rect 29595 25140 29607 25143
rect 29638 25140 29644 25152
rect 29595 25112 29644 25140
rect 29595 25109 29607 25112
rect 29549 25103 29607 25109
rect 29638 25100 29644 25112
rect 29696 25100 29702 25152
rect 30006 25100 30012 25152
rect 30064 25100 30070 25152
rect 30760 25149 30788 25384
rect 37090 25344 37096 25356
rect 37051 25316 37096 25344
rect 37090 25304 37096 25316
rect 37148 25304 37154 25356
rect 39960 25344 39988 25452
rect 40218 25440 40224 25452
rect 40276 25440 40282 25492
rect 37936 25316 39988 25344
rect 32677 25279 32735 25285
rect 32677 25245 32689 25279
rect 32723 25276 32735 25279
rect 33134 25276 33140 25288
rect 32723 25248 33140 25276
rect 32723 25245 32735 25248
rect 32677 25239 32735 25245
rect 33134 25236 33140 25248
rect 33192 25276 33198 25288
rect 34054 25276 34060 25288
rect 33192 25248 34060 25276
rect 33192 25236 33198 25248
rect 34054 25236 34060 25248
rect 34112 25236 34118 25288
rect 37366 25236 37372 25288
rect 37424 25276 37430 25288
rect 37936 25285 37964 25316
rect 37783 25279 37841 25285
rect 37783 25276 37795 25279
rect 37424 25248 37795 25276
rect 37424 25236 37430 25248
rect 37783 25245 37795 25248
rect 37829 25245 37841 25279
rect 37783 25239 37841 25245
rect 37934 25279 37992 25285
rect 37934 25245 37946 25279
rect 37980 25245 37992 25279
rect 38034 25279 38092 25285
rect 38034 25276 38046 25279
rect 37934 25239 37992 25245
rect 38028 25245 38046 25276
rect 38080 25245 38092 25279
rect 38028 25239 38092 25245
rect 38197 25279 38255 25285
rect 38197 25245 38209 25279
rect 38243 25276 38255 25279
rect 38930 25276 38936 25288
rect 38243 25248 38424 25276
rect 38843 25248 38936 25276
rect 38243 25245 38255 25248
rect 38197 25239 38255 25245
rect 32030 25168 32036 25220
rect 32088 25208 32094 25220
rect 32410 25211 32468 25217
rect 32410 25208 32422 25211
rect 32088 25180 32422 25208
rect 32088 25168 32094 25180
rect 32410 25177 32422 25180
rect 32456 25177 32468 25211
rect 32410 25171 32468 25177
rect 36848 25211 36906 25217
rect 36848 25177 36860 25211
rect 36894 25208 36906 25211
rect 37553 25211 37611 25217
rect 37553 25208 37565 25211
rect 36894 25180 37565 25208
rect 36894 25177 36906 25180
rect 36848 25171 36906 25177
rect 37553 25177 37565 25180
rect 37599 25177 37611 25211
rect 37553 25171 37611 25177
rect 37642 25168 37648 25220
rect 37700 25208 37706 25220
rect 38028 25208 38056 25239
rect 37700 25180 38056 25208
rect 37700 25168 37706 25180
rect 30745 25143 30803 25149
rect 30745 25109 30757 25143
rect 30791 25140 30803 25143
rect 32490 25140 32496 25152
rect 30791 25112 32496 25140
rect 30791 25109 30803 25112
rect 30745 25103 30803 25109
rect 32490 25100 32496 25112
rect 32548 25100 32554 25152
rect 35618 25100 35624 25152
rect 35676 25140 35682 25152
rect 35713 25143 35771 25149
rect 35713 25140 35725 25143
rect 35676 25112 35725 25140
rect 35676 25100 35682 25112
rect 35713 25109 35725 25112
rect 35759 25109 35771 25143
rect 38396 25140 38424 25248
rect 38930 25236 38936 25248
rect 38988 25276 38994 25288
rect 39850 25276 39856 25288
rect 38988 25248 39856 25276
rect 38988 25236 38994 25248
rect 39850 25236 39856 25248
rect 39908 25236 39914 25288
rect 40126 25276 40132 25288
rect 40087 25248 40132 25276
rect 40126 25236 40132 25248
rect 40184 25236 40190 25288
rect 40236 25285 40264 25440
rect 40218 25279 40276 25285
rect 40218 25245 40230 25279
rect 40264 25245 40276 25279
rect 40218 25239 40276 25245
rect 40313 25279 40371 25285
rect 40313 25245 40325 25279
rect 40359 25276 40371 25279
rect 40509 25279 40567 25285
rect 40359 25248 40448 25276
rect 40359 25245 40371 25248
rect 40313 25239 40371 25245
rect 40420 25220 40448 25248
rect 40509 25245 40521 25279
rect 40555 25276 40567 25279
rect 58158 25276 58164 25288
rect 40555 25248 40632 25276
rect 58119 25248 58164 25276
rect 40555 25245 40567 25248
rect 40509 25239 40567 25245
rect 38562 25168 38568 25220
rect 38620 25208 38626 25220
rect 39117 25211 39175 25217
rect 39117 25208 39129 25211
rect 38620 25180 39129 25208
rect 38620 25168 38626 25180
rect 39117 25177 39129 25180
rect 39163 25177 39175 25211
rect 39117 25171 39175 25177
rect 40402 25168 40408 25220
rect 40460 25168 40466 25220
rect 40604 25208 40632 25248
rect 58158 25236 58164 25248
rect 58216 25236 58222 25288
rect 40512 25180 40632 25208
rect 40512 25152 40540 25180
rect 40494 25140 40500 25152
rect 38396 25112 40500 25140
rect 35713 25103 35771 25109
rect 40494 25100 40500 25112
rect 40552 25100 40558 25152
rect 40862 25100 40868 25152
rect 40920 25140 40926 25152
rect 40957 25143 41015 25149
rect 40957 25140 40969 25143
rect 40920 25112 40969 25140
rect 40920 25100 40926 25112
rect 40957 25109 40969 25112
rect 41003 25109 41015 25143
rect 40957 25103 41015 25109
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 3878 24936 3884 24948
rect 3839 24908 3884 24936
rect 3878 24896 3884 24908
rect 3936 24896 3942 24948
rect 5902 24896 5908 24948
rect 5960 24936 5966 24948
rect 6457 24939 6515 24945
rect 6457 24936 6469 24939
rect 5960 24908 6469 24936
rect 5960 24896 5966 24908
rect 6457 24905 6469 24908
rect 6503 24936 6515 24939
rect 7282 24936 7288 24948
rect 6503 24908 7288 24936
rect 6503 24905 6515 24908
rect 6457 24899 6515 24905
rect 7282 24896 7288 24908
rect 7340 24896 7346 24948
rect 8849 24939 8907 24945
rect 8849 24905 8861 24939
rect 8895 24936 8907 24939
rect 8895 24908 10180 24936
rect 8895 24905 8907 24908
rect 8849 24899 8907 24905
rect 2774 24809 2780 24812
rect 2768 24763 2780 24809
rect 2832 24800 2838 24812
rect 2832 24772 2868 24800
rect 2774 24760 2780 24763
rect 2832 24760 2838 24772
rect 5718 24760 5724 24812
rect 5776 24800 5782 24812
rect 7190 24800 7196 24812
rect 5776 24772 7196 24800
rect 5776 24760 5782 24772
rect 7190 24760 7196 24772
rect 7248 24760 7254 24812
rect 9030 24800 9036 24812
rect 8991 24772 9036 24800
rect 9030 24760 9036 24772
rect 9088 24760 9094 24812
rect 9217 24803 9275 24809
rect 9217 24769 9229 24803
rect 9263 24800 9275 24803
rect 9582 24800 9588 24812
rect 9263 24772 9588 24800
rect 9263 24769 9275 24772
rect 9217 24763 9275 24769
rect 9582 24760 9588 24772
rect 9640 24760 9646 24812
rect 10152 24809 10180 24908
rect 22664 24908 27476 24936
rect 22664 24877 22692 24908
rect 22649 24871 22707 24877
rect 18984 24840 19288 24868
rect 9907 24803 9965 24809
rect 9907 24800 9919 24803
rect 9784 24772 9919 24800
rect 2406 24692 2412 24744
rect 2464 24732 2470 24744
rect 2501 24735 2559 24741
rect 2501 24732 2513 24735
rect 2464 24704 2513 24732
rect 2464 24692 2470 24704
rect 2501 24701 2513 24704
rect 2547 24701 2559 24735
rect 9784 24732 9812 24772
rect 9907 24769 9919 24772
rect 9953 24769 9965 24803
rect 9907 24763 9965 24769
rect 10045 24803 10103 24809
rect 10045 24769 10057 24803
rect 10091 24769 10103 24803
rect 10045 24763 10103 24769
rect 10137 24803 10195 24809
rect 10137 24769 10149 24803
rect 10183 24769 10195 24803
rect 10318 24800 10324 24812
rect 10279 24772 10324 24800
rect 10137 24763 10195 24769
rect 2501 24695 2559 24701
rect 8266 24704 9812 24732
rect 7190 24624 7196 24676
rect 7248 24664 7254 24676
rect 8266 24664 8294 24704
rect 7248 24636 8294 24664
rect 7248 24624 7254 24636
rect 9674 24596 9680 24608
rect 9635 24568 9680 24596
rect 9674 24556 9680 24568
rect 9732 24556 9738 24608
rect 9784 24596 9812 24704
rect 9950 24624 9956 24676
rect 10008 24664 10014 24676
rect 10060 24664 10088 24763
rect 10318 24760 10324 24772
rect 10376 24760 10382 24812
rect 13541 24803 13599 24809
rect 13541 24769 13553 24803
rect 13587 24769 13599 24803
rect 13722 24800 13728 24812
rect 13683 24772 13728 24800
rect 13541 24763 13599 24769
rect 12434 24692 12440 24744
rect 12492 24732 12498 24744
rect 12529 24735 12587 24741
rect 12529 24732 12541 24735
rect 12492 24704 12541 24732
rect 12492 24692 12498 24704
rect 12529 24701 12541 24704
rect 12575 24701 12587 24735
rect 13556 24732 13584 24763
rect 13722 24760 13728 24772
rect 13780 24760 13786 24812
rect 14366 24760 14372 24812
rect 14424 24800 14430 24812
rect 14717 24803 14775 24809
rect 14717 24800 14729 24803
rect 14424 24772 14729 24800
rect 14424 24760 14430 24772
rect 14717 24769 14729 24772
rect 14763 24769 14775 24803
rect 14717 24763 14775 24769
rect 16574 24760 16580 24812
rect 16632 24800 16638 24812
rect 16945 24803 17003 24809
rect 16945 24800 16957 24803
rect 16632 24772 16957 24800
rect 16632 24760 16638 24772
rect 16945 24769 16957 24772
rect 16991 24769 17003 24803
rect 16945 24763 17003 24769
rect 18877 24803 18935 24809
rect 18877 24769 18889 24803
rect 18923 24800 18935 24803
rect 18984 24800 19012 24840
rect 19150 24809 19156 24812
rect 19144 24800 19156 24809
rect 18923 24772 19012 24800
rect 19111 24772 19156 24800
rect 18923 24769 18935 24772
rect 18877 24763 18935 24769
rect 19144 24763 19156 24772
rect 19150 24760 19156 24763
rect 19208 24760 19214 24812
rect 19260 24800 19288 24840
rect 22649 24837 22661 24871
rect 22695 24837 22707 24871
rect 27448 24868 27476 24908
rect 27522 24896 27528 24948
rect 27580 24936 27586 24948
rect 32398 24936 32404 24948
rect 27580 24908 32404 24936
rect 27580 24896 27586 24908
rect 32398 24896 32404 24908
rect 32456 24896 32462 24948
rect 32490 24896 32496 24948
rect 32548 24936 32554 24948
rect 40126 24936 40132 24948
rect 32548 24908 40132 24936
rect 32548 24896 32554 24908
rect 40126 24896 40132 24908
rect 40184 24936 40190 24948
rect 40862 24936 40868 24948
rect 40184 24908 40868 24936
rect 40184 24896 40190 24908
rect 40862 24896 40868 24908
rect 40920 24896 40926 24948
rect 27982 24868 27988 24880
rect 22649 24831 22707 24837
rect 25240 24840 25360 24868
rect 27448 24840 27988 24868
rect 21726 24800 21732 24812
rect 19260 24772 21732 24800
rect 21726 24760 21732 24772
rect 21784 24760 21790 24812
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 22511 24803 22569 24809
rect 22511 24800 22523 24803
rect 22152 24772 22523 24800
rect 22152 24760 22158 24772
rect 22511 24769 22523 24772
rect 22557 24769 22569 24803
rect 22738 24800 22744 24812
rect 22699 24772 22744 24800
rect 22511 24763 22569 24769
rect 22738 24760 22744 24772
rect 22796 24760 22802 24812
rect 22830 24760 22836 24812
rect 22888 24809 22894 24812
rect 22888 24803 22927 24809
rect 22915 24769 22927 24803
rect 22888 24763 22927 24769
rect 22888 24760 22894 24763
rect 23014 24760 23020 24812
rect 23072 24800 23078 24812
rect 24670 24800 24676 24812
rect 23072 24772 23117 24800
rect 23317 24772 24676 24800
rect 23072 24760 23078 24772
rect 14182 24732 14188 24744
rect 13556 24704 14188 24732
rect 12529 24695 12587 24701
rect 14182 24692 14188 24704
rect 14240 24692 14246 24744
rect 14461 24735 14519 24741
rect 14461 24701 14473 24735
rect 14507 24701 14519 24735
rect 14461 24695 14519 24701
rect 10008 24636 10088 24664
rect 10008 24624 10014 24636
rect 10134 24624 10140 24676
rect 10192 24664 10198 24676
rect 12618 24664 12624 24676
rect 10192 24636 12624 24664
rect 10192 24624 10198 24636
rect 12618 24624 12624 24636
rect 12676 24624 12682 24676
rect 10781 24599 10839 24605
rect 10781 24596 10793 24599
rect 9784 24568 10793 24596
rect 10781 24565 10793 24568
rect 10827 24565 10839 24599
rect 10781 24559 10839 24565
rect 12069 24599 12127 24605
rect 12069 24565 12081 24599
rect 12115 24596 12127 24599
rect 12250 24596 12256 24608
rect 12115 24568 12256 24596
rect 12115 24565 12127 24568
rect 12069 24559 12127 24565
rect 12250 24556 12256 24568
rect 12308 24556 12314 24608
rect 13170 24556 13176 24608
rect 13228 24596 13234 24608
rect 13357 24599 13415 24605
rect 13357 24596 13369 24599
rect 13228 24568 13369 24596
rect 13228 24556 13234 24568
rect 13357 24565 13369 24568
rect 13403 24565 13415 24599
rect 14476 24596 14504 24695
rect 17770 24692 17776 24744
rect 17828 24732 17834 24744
rect 18141 24735 18199 24741
rect 18141 24732 18153 24735
rect 17828 24704 18153 24732
rect 17828 24692 17834 24704
rect 18141 24701 18153 24704
rect 18187 24701 18199 24735
rect 18141 24695 18199 24701
rect 18417 24735 18475 24741
rect 18417 24701 18429 24735
rect 18463 24701 18475 24735
rect 18417 24695 18475 24701
rect 16482 24664 16488 24676
rect 15396 24636 16488 24664
rect 15194 24596 15200 24608
rect 14476 24568 15200 24596
rect 13357 24559 13415 24565
rect 15194 24556 15200 24568
rect 15252 24596 15258 24608
rect 15396 24596 15424 24636
rect 16482 24624 16488 24636
rect 16540 24624 16546 24676
rect 15838 24596 15844 24608
rect 15252 24568 15424 24596
rect 15799 24568 15844 24596
rect 15252 24556 15258 24568
rect 15838 24556 15844 24568
rect 15896 24556 15902 24608
rect 16298 24556 16304 24608
rect 16356 24596 16362 24608
rect 16761 24599 16819 24605
rect 16761 24596 16773 24599
rect 16356 24568 16773 24596
rect 16356 24556 16362 24568
rect 16761 24565 16773 24568
rect 16807 24565 16819 24599
rect 18432 24596 18460 24695
rect 20898 24692 20904 24744
rect 20956 24732 20962 24744
rect 23317 24732 23345 24772
rect 24670 24760 24676 24772
rect 24728 24800 24734 24812
rect 24857 24803 24915 24809
rect 24857 24800 24869 24803
rect 24728 24772 24869 24800
rect 24728 24760 24734 24772
rect 24857 24769 24869 24772
rect 24903 24769 24915 24803
rect 25038 24800 25044 24812
rect 24999 24772 25044 24800
rect 24857 24763 24915 24769
rect 25038 24760 25044 24772
rect 25096 24760 25102 24812
rect 25240 24809 25268 24840
rect 25133 24803 25191 24809
rect 25133 24769 25145 24803
rect 25179 24769 25191 24803
rect 25133 24763 25191 24769
rect 25225 24803 25283 24809
rect 25225 24769 25237 24803
rect 25271 24769 25283 24803
rect 25225 24763 25283 24769
rect 20956 24704 23345 24732
rect 20956 24692 20962 24704
rect 24762 24692 24768 24744
rect 24820 24732 24826 24744
rect 25148 24732 25176 24763
rect 24820 24704 25176 24732
rect 24820 24692 24826 24704
rect 19886 24624 19892 24676
rect 19944 24664 19950 24676
rect 19944 24636 20300 24664
rect 19944 24624 19950 24636
rect 18506 24596 18512 24608
rect 18419 24568 18512 24596
rect 16761 24559 16819 24565
rect 18506 24556 18512 24568
rect 18564 24596 18570 24608
rect 20070 24596 20076 24608
rect 18564 24568 20076 24596
rect 18564 24556 18570 24568
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 20272 24605 20300 24636
rect 20438 24624 20444 24676
rect 20496 24664 20502 24676
rect 21634 24664 21640 24676
rect 20496 24636 21640 24664
rect 20496 24624 20502 24636
rect 21634 24624 21640 24636
rect 21692 24664 21698 24676
rect 24397 24667 24455 24673
rect 24397 24664 24409 24667
rect 21692 24636 24409 24664
rect 21692 24624 21698 24636
rect 24397 24633 24409 24636
rect 24443 24664 24455 24667
rect 25332 24664 25360 24840
rect 27982 24828 27988 24840
rect 28040 24828 28046 24880
rect 28994 24828 29000 24880
rect 29052 24868 29058 24880
rect 29730 24868 29736 24880
rect 29052 24840 29736 24868
rect 29052 24828 29058 24840
rect 29730 24828 29736 24840
rect 29788 24868 29794 24880
rect 29788 24840 30972 24868
rect 29788 24828 29794 24840
rect 29937 24803 29995 24809
rect 29937 24769 29949 24803
rect 29983 24800 29995 24803
rect 30098 24800 30104 24812
rect 29983 24772 30104 24800
rect 29983 24769 29995 24772
rect 29937 24763 29995 24769
rect 30098 24760 30104 24772
rect 30156 24760 30162 24812
rect 30650 24800 30656 24812
rect 30611 24772 30656 24800
rect 30650 24760 30656 24772
rect 30708 24760 30714 24812
rect 30742 24760 30748 24812
rect 30800 24800 30806 24812
rect 30837 24806 30895 24812
rect 30944 24809 30972 24840
rect 37384 24840 37596 24868
rect 30837 24800 30849 24806
rect 30800 24772 30849 24800
rect 30883 24772 30895 24806
rect 30800 24760 30806 24772
rect 30837 24766 30895 24772
rect 30929 24803 30987 24809
rect 30929 24769 30941 24803
rect 30975 24769 30987 24803
rect 30929 24763 30987 24769
rect 31021 24803 31079 24809
rect 32125 24803 32183 24809
rect 31021 24769 31033 24803
rect 31067 24800 31156 24803
rect 32125 24800 32137 24803
rect 31067 24775 32137 24800
rect 31067 24769 31079 24775
rect 31128 24772 32137 24775
rect 31021 24763 31079 24769
rect 32125 24769 32137 24772
rect 32171 24800 32183 24803
rect 33505 24803 33563 24809
rect 32171 24772 33134 24800
rect 32171 24769 32183 24772
rect 32125 24763 32183 24769
rect 30193 24735 30251 24741
rect 30193 24701 30205 24735
rect 30239 24701 30251 24735
rect 30193 24695 30251 24701
rect 31297 24735 31355 24741
rect 31297 24701 31309 24735
rect 31343 24732 31355 24735
rect 32030 24732 32036 24744
rect 31343 24704 32036 24732
rect 31343 24701 31355 24704
rect 31297 24695 31355 24701
rect 24443 24636 25360 24664
rect 24443 24633 24455 24636
rect 24397 24627 24455 24633
rect 20257 24599 20315 24605
rect 20257 24565 20269 24599
rect 20303 24596 20315 24599
rect 21542 24596 21548 24608
rect 20303 24568 21548 24596
rect 20303 24565 20315 24568
rect 20257 24559 20315 24565
rect 21542 24556 21548 24568
rect 21600 24556 21606 24608
rect 22186 24556 22192 24608
rect 22244 24596 22250 24608
rect 22373 24599 22431 24605
rect 22373 24596 22385 24599
rect 22244 24568 22385 24596
rect 22244 24556 22250 24568
rect 22373 24565 22385 24568
rect 22419 24565 22431 24599
rect 25498 24596 25504 24608
rect 25459 24568 25504 24596
rect 22373 24559 22431 24565
rect 25498 24556 25504 24568
rect 25556 24556 25562 24608
rect 28258 24596 28264 24608
rect 28219 24568 28264 24596
rect 28258 24556 28264 24568
rect 28316 24556 28322 24608
rect 28810 24596 28816 24608
rect 28771 24568 28816 24596
rect 28810 24556 28816 24568
rect 28868 24556 28874 24608
rect 28902 24556 28908 24608
rect 28960 24596 28966 24608
rect 30208 24596 30236 24695
rect 32030 24692 32036 24704
rect 32088 24692 32094 24744
rect 28960 24568 30236 24596
rect 33106 24596 33134 24772
rect 33505 24769 33517 24803
rect 33551 24800 33563 24803
rect 33962 24800 33968 24812
rect 33551 24772 33968 24800
rect 33551 24769 33563 24772
rect 33505 24763 33563 24769
rect 33962 24760 33968 24772
rect 34020 24760 34026 24812
rect 37277 24803 37335 24809
rect 37277 24769 37289 24803
rect 37323 24800 37335 24803
rect 37384 24800 37412 24840
rect 37323 24772 37412 24800
rect 37461 24803 37519 24809
rect 37323 24769 37335 24772
rect 37277 24763 37335 24769
rect 37461 24769 37473 24803
rect 37507 24769 37519 24803
rect 37568 24800 37596 24840
rect 38930 24800 38936 24812
rect 37568 24772 38936 24800
rect 37461 24763 37519 24769
rect 35710 24732 35716 24744
rect 35671 24704 35716 24732
rect 35710 24692 35716 24704
rect 35768 24692 35774 24744
rect 35618 24624 35624 24676
rect 35676 24664 35682 24676
rect 37476 24664 37504 24763
rect 38930 24760 38936 24772
rect 38988 24760 38994 24812
rect 39758 24800 39764 24812
rect 39816 24809 39822 24812
rect 39728 24772 39764 24800
rect 39758 24760 39764 24772
rect 39816 24763 39828 24809
rect 39816 24760 39822 24763
rect 39942 24760 39948 24812
rect 40000 24800 40006 24812
rect 40037 24803 40095 24809
rect 40037 24800 40049 24803
rect 40000 24772 40049 24800
rect 40000 24760 40006 24772
rect 40037 24769 40049 24772
rect 40083 24769 40095 24803
rect 40037 24763 40095 24769
rect 37642 24732 37648 24744
rect 37603 24704 37648 24732
rect 37642 24692 37648 24704
rect 37700 24692 37706 24744
rect 35676 24636 37504 24664
rect 35676 24624 35682 24636
rect 33870 24596 33876 24608
rect 33106 24568 33876 24596
rect 28960 24556 28966 24568
rect 33870 24556 33876 24568
rect 33928 24556 33934 24608
rect 36078 24556 36084 24608
rect 36136 24596 36142 24608
rect 38654 24596 38660 24608
rect 36136 24568 38660 24596
rect 36136 24556 36142 24568
rect 38654 24556 38660 24568
rect 38712 24556 38718 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 9950 24352 9956 24404
rect 10008 24392 10014 24404
rect 10008 24364 10364 24392
rect 10008 24352 10014 24364
rect 10336 24324 10364 24364
rect 11882 24352 11888 24404
rect 11940 24392 11946 24404
rect 14366 24392 14372 24404
rect 11940 24364 12434 24392
rect 14327 24364 14372 24392
rect 11940 24352 11946 24364
rect 12406 24324 12434 24364
rect 14366 24352 14372 24364
rect 14424 24352 14430 24404
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 15930 24392 15936 24404
rect 15519 24364 15936 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 13538 24324 13544 24336
rect 10336 24296 12020 24324
rect 12406 24296 13544 24324
rect 10321 24259 10379 24265
rect 10321 24225 10333 24259
rect 10367 24256 10379 24259
rect 11054 24256 11060 24268
rect 10367 24228 11060 24256
rect 10367 24225 10379 24228
rect 10321 24219 10379 24225
rect 11054 24216 11060 24228
rect 11112 24216 11118 24268
rect 11992 24256 12020 24296
rect 13538 24284 13544 24296
rect 13596 24284 13602 24336
rect 13722 24284 13728 24336
rect 13780 24324 13786 24336
rect 15562 24324 15568 24336
rect 13780 24296 15568 24324
rect 13780 24284 13786 24296
rect 15562 24284 15568 24296
rect 15620 24284 15626 24336
rect 13906 24256 13912 24268
rect 11992 24228 13912 24256
rect 9674 24148 9680 24200
rect 9732 24188 9738 24200
rect 10054 24191 10112 24197
rect 10054 24188 10066 24191
rect 9732 24160 10066 24188
rect 9732 24148 9738 24160
rect 10054 24157 10066 24160
rect 10100 24157 10112 24191
rect 10054 24151 10112 24157
rect 11238 24148 11244 24200
rect 11296 24188 11302 24200
rect 11882 24188 11888 24200
rect 11296 24160 11888 24188
rect 11296 24148 11302 24160
rect 11882 24148 11888 24160
rect 11940 24148 11946 24200
rect 11992 24197 12020 24228
rect 11977 24191 12035 24197
rect 11977 24157 11989 24191
rect 12023 24157 12035 24191
rect 11977 24151 12035 24157
rect 12066 24148 12072 24200
rect 12124 24188 12130 24200
rect 12124 24160 12169 24188
rect 12124 24148 12130 24160
rect 12250 24148 12256 24200
rect 12308 24188 12314 24200
rect 12308 24160 12401 24188
rect 12308 24148 12314 24160
rect 12434 24148 12440 24200
rect 12492 24188 12498 24200
rect 13096 24197 13124 24228
rect 13906 24216 13912 24228
rect 13964 24216 13970 24268
rect 12989 24191 13047 24197
rect 12989 24188 13001 24191
rect 12492 24160 13001 24188
rect 12492 24148 12498 24160
rect 12989 24157 13001 24160
rect 13035 24157 13047 24191
rect 12989 24151 13047 24157
rect 13081 24191 13139 24197
rect 13081 24157 13093 24191
rect 13127 24157 13139 24191
rect 13081 24151 13139 24157
rect 13170 24148 13176 24200
rect 13228 24188 13234 24200
rect 13228 24160 13273 24188
rect 13228 24148 13234 24160
rect 13354 24148 13360 24200
rect 13412 24188 13418 24200
rect 14642 24188 14648 24200
rect 13412 24160 13457 24188
rect 14603 24160 14648 24188
rect 13412 24148 13418 24160
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 14734 24188 14792 24194
rect 14734 24154 14746 24188
rect 14780 24154 14792 24188
rect 14734 24148 14792 24154
rect 14826 24148 14832 24200
rect 14884 24197 14890 24200
rect 14884 24188 14892 24197
rect 15013 24191 15071 24197
rect 14884 24160 14929 24188
rect 14884 24151 14892 24160
rect 15013 24157 15025 24191
rect 15059 24188 15071 24191
rect 15672 24188 15700 24364
rect 15930 24352 15936 24364
rect 15988 24352 15994 24404
rect 18230 24352 18236 24404
rect 18288 24392 18294 24404
rect 19245 24395 19303 24401
rect 19245 24392 19257 24395
rect 18288 24364 19257 24392
rect 18288 24352 18294 24364
rect 19245 24361 19257 24364
rect 19291 24361 19303 24395
rect 24581 24395 24639 24401
rect 19245 24355 19303 24361
rect 21284 24364 24348 24392
rect 16942 24284 16948 24336
rect 17000 24324 17006 24336
rect 20898 24324 20904 24336
rect 17000 24296 20904 24324
rect 17000 24284 17006 24296
rect 20898 24284 20904 24296
rect 20956 24284 20962 24336
rect 18046 24216 18052 24268
rect 18104 24256 18110 24268
rect 18141 24259 18199 24265
rect 18141 24256 18153 24259
rect 18104 24228 18153 24256
rect 18104 24216 18110 24228
rect 18141 24225 18153 24228
rect 18187 24225 18199 24259
rect 18141 24219 18199 24225
rect 18414 24188 18420 24200
rect 15059 24160 15700 24188
rect 18375 24160 18420 24188
rect 15059 24157 15071 24160
rect 15013 24151 15071 24157
rect 14884 24148 14890 24151
rect 18414 24148 18420 24160
rect 18472 24148 18478 24200
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24188 19487 24191
rect 19886 24188 19892 24200
rect 19475 24160 19892 24188
rect 19475 24157 19487 24160
rect 19429 24151 19487 24157
rect 19886 24148 19892 24160
rect 19944 24148 19950 24200
rect 20949 24191 21007 24197
rect 20949 24157 20961 24191
rect 20995 24157 21007 24191
rect 20949 24151 21007 24157
rect 21085 24191 21143 24197
rect 21085 24157 21097 24191
rect 21131 24188 21143 24191
rect 21284 24188 21312 24364
rect 21910 24284 21916 24336
rect 21968 24324 21974 24336
rect 21968 24296 22508 24324
rect 21968 24284 21974 24296
rect 21542 24256 21548 24268
rect 21376 24228 21548 24256
rect 21376 24197 21404 24228
rect 21542 24216 21548 24228
rect 21600 24216 21606 24268
rect 21131 24160 21312 24188
rect 21360 24191 21418 24197
rect 21131 24157 21143 24160
rect 21085 24151 21143 24157
rect 21360 24157 21372 24191
rect 21406 24157 21418 24191
rect 21360 24151 21418 24157
rect 7834 24120 7840 24132
rect 7747 24092 7840 24120
rect 7834 24080 7840 24092
rect 7892 24120 7898 24132
rect 10134 24120 10140 24132
rect 7892 24092 10140 24120
rect 7892 24080 7898 24092
rect 10134 24080 10140 24092
rect 10192 24080 10198 24132
rect 12268 24120 12296 24148
rect 13372 24120 13400 24148
rect 12268 24092 13400 24120
rect 8941 24055 8999 24061
rect 8941 24021 8953 24055
rect 8987 24052 8999 24055
rect 9030 24052 9036 24064
rect 8987 24024 9036 24052
rect 8987 24021 8999 24024
rect 8941 24015 8999 24021
rect 9030 24012 9036 24024
rect 9088 24052 9094 24064
rect 9950 24052 9956 24064
rect 9088 24024 9956 24052
rect 9088 24012 9094 24024
rect 9950 24012 9956 24024
rect 10008 24012 10014 24064
rect 11149 24055 11207 24061
rect 11149 24021 11161 24055
rect 11195 24052 11207 24055
rect 11238 24052 11244 24064
rect 11195 24024 11244 24052
rect 11195 24021 11207 24024
rect 11149 24015 11207 24021
rect 11238 24012 11244 24024
rect 11296 24012 11302 24064
rect 11606 24052 11612 24064
rect 11567 24024 11612 24052
rect 11606 24012 11612 24024
rect 11664 24012 11670 24064
rect 12713 24055 12771 24061
rect 12713 24021 12725 24055
rect 12759 24052 12771 24055
rect 12894 24052 12900 24064
rect 12759 24024 12900 24052
rect 12759 24021 12771 24024
rect 12713 24015 12771 24021
rect 12894 24012 12900 24024
rect 12952 24012 12958 24064
rect 13906 24012 13912 24064
rect 13964 24052 13970 24064
rect 14752 24052 14780 24148
rect 18230 24080 18236 24132
rect 18288 24120 18294 24132
rect 19242 24120 19248 24132
rect 18288 24092 19248 24120
rect 18288 24080 18294 24092
rect 19242 24080 19248 24092
rect 19300 24120 19306 24132
rect 19613 24123 19671 24129
rect 19613 24120 19625 24123
rect 19300 24092 19625 24120
rect 19300 24080 19306 24092
rect 19613 24089 19625 24092
rect 19659 24089 19671 24123
rect 20964 24120 20992 24151
rect 21450 24148 21456 24200
rect 21508 24188 21514 24200
rect 22094 24197 22100 24200
rect 22051 24191 22100 24197
rect 22051 24188 22063 24191
rect 21508 24160 21553 24188
rect 21744 24160 22063 24188
rect 21508 24148 21514 24160
rect 21177 24123 21235 24129
rect 20964 24092 21036 24120
rect 19613 24083 19671 24089
rect 16574 24052 16580 24064
rect 13964 24024 14780 24052
rect 16535 24024 16580 24052
rect 13964 24012 13970 24024
rect 16574 24012 16580 24024
rect 16632 24012 16638 24064
rect 20809 24055 20867 24061
rect 20809 24021 20821 24055
rect 20855 24052 20867 24055
rect 20898 24052 20904 24064
rect 20855 24024 20904 24052
rect 20855 24021 20867 24024
rect 20809 24015 20867 24021
rect 20898 24012 20904 24024
rect 20956 24012 20962 24064
rect 21008 24052 21036 24092
rect 21177 24089 21189 24123
rect 21223 24120 21235 24123
rect 21266 24120 21272 24132
rect 21223 24092 21272 24120
rect 21223 24089 21235 24092
rect 21177 24083 21235 24089
rect 21266 24080 21272 24092
rect 21324 24080 21330 24132
rect 21450 24052 21456 24064
rect 21008 24024 21456 24052
rect 21450 24012 21456 24024
rect 21508 24052 21514 24064
rect 21744 24052 21772 24160
rect 22051 24157 22063 24160
rect 22097 24157 22100 24191
rect 22051 24151 22100 24157
rect 22094 24148 22100 24151
rect 22152 24188 22158 24200
rect 22480 24197 22508 24296
rect 22554 24284 22560 24336
rect 22612 24284 22618 24336
rect 22572 24197 22600 24284
rect 22281 24191 22339 24197
rect 22152 24160 22199 24188
rect 22152 24148 22158 24160
rect 22281 24157 22293 24191
rect 22327 24188 22339 24191
rect 22464 24191 22522 24197
rect 22327 24160 22416 24188
rect 22327 24157 22339 24160
rect 22281 24151 22339 24157
rect 22189 24123 22247 24129
rect 22189 24089 22201 24123
rect 22235 24120 22247 24123
rect 22388 24120 22416 24160
rect 22464 24157 22476 24191
rect 22510 24157 22522 24191
rect 22464 24151 22522 24157
rect 22557 24191 22615 24197
rect 22557 24157 22569 24191
rect 22603 24157 22615 24191
rect 22557 24151 22615 24157
rect 22738 24120 22744 24132
rect 22235 24092 22324 24120
rect 22388 24092 22744 24120
rect 22235 24089 22247 24092
rect 22189 24083 22247 24089
rect 21910 24052 21916 24064
rect 21508 24024 21772 24052
rect 21871 24024 21916 24052
rect 21508 24012 21514 24024
rect 21910 24012 21916 24024
rect 21968 24012 21974 24064
rect 22296 24052 22324 24092
rect 22738 24080 22744 24092
rect 22796 24080 22802 24132
rect 24118 24052 24124 24064
rect 22296 24024 24124 24052
rect 24118 24012 24124 24024
rect 24176 24012 24182 24064
rect 24320 24052 24348 24364
rect 24581 24361 24593 24395
rect 24627 24392 24639 24395
rect 25038 24392 25044 24404
rect 24627 24364 25044 24392
rect 24627 24361 24639 24364
rect 24581 24355 24639 24361
rect 25038 24352 25044 24364
rect 25096 24352 25102 24404
rect 26786 24392 26792 24404
rect 25148 24364 26792 24392
rect 25148 24256 25176 24364
rect 26786 24352 26792 24364
rect 26844 24352 26850 24404
rect 28169 24395 28227 24401
rect 28169 24361 28181 24395
rect 28215 24392 28227 24395
rect 30006 24392 30012 24404
rect 28215 24364 30012 24392
rect 28215 24361 28227 24364
rect 28169 24355 28227 24361
rect 30006 24352 30012 24364
rect 30064 24352 30070 24404
rect 30098 24352 30104 24404
rect 30156 24392 30162 24404
rect 30193 24395 30251 24401
rect 30193 24392 30205 24395
rect 30156 24364 30205 24392
rect 30156 24352 30162 24364
rect 30193 24361 30205 24364
rect 30239 24361 30251 24395
rect 30193 24355 30251 24361
rect 28258 24284 28264 24336
rect 28316 24324 28322 24336
rect 30650 24324 30656 24336
rect 28316 24296 30656 24324
rect 28316 24284 28322 24296
rect 24780 24228 25176 24256
rect 24780 24197 24808 24228
rect 27798 24216 27804 24268
rect 27856 24256 27862 24268
rect 28626 24256 28632 24268
rect 27856 24228 28632 24256
rect 27856 24216 27862 24228
rect 28626 24216 28632 24228
rect 28684 24216 28690 24268
rect 24765 24191 24823 24197
rect 24765 24157 24777 24191
rect 24811 24157 24823 24191
rect 24946 24188 24952 24200
rect 24907 24160 24952 24188
rect 24765 24151 24823 24157
rect 24946 24148 24952 24160
rect 25004 24148 25010 24200
rect 25406 24188 25412 24200
rect 25367 24160 25412 24188
rect 25406 24148 25412 24160
rect 25464 24188 25470 24200
rect 27614 24188 27620 24200
rect 25464 24160 27620 24188
rect 25464 24148 25470 24160
rect 27614 24148 27620 24160
rect 27672 24148 27678 24200
rect 28810 24188 28816 24200
rect 27724 24160 28816 24188
rect 25498 24080 25504 24132
rect 25556 24120 25562 24132
rect 25654 24123 25712 24129
rect 25654 24120 25666 24123
rect 25556 24092 25666 24120
rect 25556 24080 25562 24092
rect 25654 24089 25666 24092
rect 25700 24089 25712 24123
rect 27724 24120 27752 24160
rect 28810 24148 28816 24160
rect 28868 24148 28874 24200
rect 29012 24188 29040 24296
rect 30650 24284 30656 24296
rect 30708 24284 30714 24336
rect 29086 24216 29092 24268
rect 29144 24256 29150 24268
rect 29144 24228 29855 24256
rect 29144 24216 29150 24228
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 29012 24160 29561 24188
rect 29549 24157 29561 24160
rect 29595 24157 29607 24191
rect 29712 24191 29770 24197
rect 29827 24194 29855 24228
rect 38654 24216 38660 24268
rect 38712 24256 38718 24268
rect 38712 24228 40264 24256
rect 38712 24216 38718 24228
rect 40236 24197 40264 24228
rect 29712 24188 29724 24191
rect 29549 24151 29607 24157
rect 29656 24160 29724 24188
rect 25654 24083 25712 24089
rect 25780 24092 27752 24120
rect 25780 24052 25808 24092
rect 27798 24080 27804 24132
rect 27856 24120 27862 24132
rect 27856 24092 27901 24120
rect 27856 24080 27862 24092
rect 27982 24080 27988 24132
rect 28040 24120 28046 24132
rect 28626 24120 28632 24132
rect 28040 24092 28085 24120
rect 28587 24092 28632 24120
rect 28040 24080 28046 24092
rect 28626 24080 28632 24092
rect 28684 24080 28690 24132
rect 29656 24120 29684 24160
rect 29712 24157 29724 24160
rect 29758 24157 29770 24191
rect 29712 24151 29770 24157
rect 29812 24188 29870 24194
rect 29812 24154 29824 24188
rect 29858 24154 29870 24188
rect 29812 24148 29870 24154
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24157 29975 24191
rect 29917 24151 29975 24157
rect 40221 24191 40279 24197
rect 40221 24157 40233 24191
rect 40267 24157 40279 24191
rect 41046 24188 41052 24200
rect 41007 24160 41052 24188
rect 40221 24151 40279 24157
rect 29012 24092 29684 24120
rect 24320 24024 25808 24052
rect 26786 24012 26792 24064
rect 26844 24052 26850 24064
rect 28166 24052 28172 24064
rect 26844 24024 28172 24052
rect 26844 24012 26850 24024
rect 28166 24012 28172 24024
rect 28224 24012 28230 24064
rect 29012 24061 29040 24092
rect 29932 24064 29960 24151
rect 41046 24148 41052 24160
rect 41104 24148 41110 24200
rect 58158 24188 58164 24200
rect 58119 24160 58164 24188
rect 58158 24148 58164 24160
rect 58216 24148 58222 24200
rect 39850 24080 39856 24132
rect 39908 24120 39914 24132
rect 40037 24123 40095 24129
rect 40037 24120 40049 24123
rect 39908 24092 40049 24120
rect 39908 24080 39914 24092
rect 40037 24089 40049 24092
rect 40083 24120 40095 24123
rect 40865 24123 40923 24129
rect 40865 24120 40877 24123
rect 40083 24092 40877 24120
rect 40083 24089 40095 24092
rect 40037 24083 40095 24089
rect 40865 24089 40877 24092
rect 40911 24089 40923 24123
rect 40865 24083 40923 24089
rect 28997 24055 29055 24061
rect 28997 24021 29009 24055
rect 29043 24021 29055 24055
rect 28997 24015 29055 24021
rect 29914 24012 29920 24064
rect 29972 24012 29978 24064
rect 40402 24052 40408 24064
rect 40363 24024 40408 24052
rect 40402 24012 40408 24024
rect 40460 24012 40466 24064
rect 41138 24012 41144 24064
rect 41196 24052 41202 24064
rect 41233 24055 41291 24061
rect 41233 24052 41245 24055
rect 41196 24024 41245 24052
rect 41196 24012 41202 24024
rect 41233 24021 41245 24024
rect 41279 24021 41291 24055
rect 41233 24015 41291 24021
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 9766 23808 9772 23860
rect 9824 23848 9830 23860
rect 10137 23851 10195 23857
rect 10137 23848 10149 23851
rect 9824 23820 10149 23848
rect 9824 23808 9830 23820
rect 10137 23817 10149 23820
rect 10183 23817 10195 23851
rect 10137 23811 10195 23817
rect 12066 23808 12072 23860
rect 12124 23848 12130 23860
rect 12161 23851 12219 23857
rect 12161 23848 12173 23851
rect 12124 23820 12173 23848
rect 12124 23808 12130 23820
rect 12161 23817 12173 23820
rect 12207 23817 12219 23851
rect 13722 23848 13728 23860
rect 12161 23811 12219 23817
rect 12406 23820 13728 23848
rect 11054 23780 11060 23792
rect 8312 23752 11060 23780
rect 2222 23712 2228 23724
rect 2183 23684 2228 23712
rect 2222 23672 2228 23684
rect 2280 23672 2286 23724
rect 2409 23715 2467 23721
rect 2409 23681 2421 23715
rect 2455 23712 2467 23715
rect 3234 23712 3240 23724
rect 2455 23684 3240 23712
rect 2455 23681 2467 23684
rect 2409 23675 2467 23681
rect 3234 23672 3240 23684
rect 3292 23672 3298 23724
rect 7653 23715 7711 23721
rect 7653 23681 7665 23715
rect 7699 23712 7711 23715
rect 7834 23712 7840 23724
rect 7699 23684 7840 23712
rect 7699 23681 7711 23684
rect 7653 23675 7711 23681
rect 7834 23672 7840 23684
rect 7892 23672 7898 23724
rect 8312 23721 8340 23752
rect 11054 23740 11060 23752
rect 11112 23740 11118 23792
rect 12406 23780 12434 23820
rect 13722 23808 13728 23820
rect 13780 23808 13786 23860
rect 14182 23848 14188 23860
rect 14143 23820 14188 23848
rect 14182 23808 14188 23820
rect 14240 23808 14246 23860
rect 14642 23848 14648 23860
rect 14603 23820 14648 23848
rect 14642 23808 14648 23820
rect 14700 23808 14706 23860
rect 18230 23848 18236 23860
rect 18191 23820 18236 23848
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 18598 23808 18604 23860
rect 18656 23848 18662 23860
rect 18656 23820 24992 23848
rect 18656 23808 18662 23820
rect 15194 23780 15200 23792
rect 11808 23752 12434 23780
rect 12820 23752 15200 23780
rect 8570 23721 8576 23724
rect 8297 23715 8355 23721
rect 8297 23681 8309 23715
rect 8343 23681 8355 23715
rect 8564 23712 8576 23721
rect 8531 23684 8576 23712
rect 8297 23675 8355 23681
rect 8564 23675 8576 23684
rect 8570 23672 8576 23675
rect 8628 23672 8634 23724
rect 10134 23672 10140 23724
rect 10192 23712 10198 23724
rect 11808 23721 11836 23752
rect 10321 23715 10379 23721
rect 10321 23712 10333 23715
rect 10192 23684 10333 23712
rect 10192 23672 10198 23684
rect 10321 23681 10333 23684
rect 10367 23681 10379 23715
rect 10321 23675 10379 23681
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23712 10563 23715
rect 11793 23715 11851 23721
rect 11793 23712 11805 23715
rect 10551 23684 11805 23712
rect 10551 23681 10563 23684
rect 10505 23675 10563 23681
rect 11793 23681 11805 23684
rect 11839 23681 11851 23715
rect 11974 23712 11980 23724
rect 11935 23684 11980 23712
rect 11793 23675 11851 23681
rect 7006 23604 7012 23656
rect 7064 23644 7070 23656
rect 7377 23647 7435 23653
rect 7377 23644 7389 23647
rect 7064 23616 7389 23644
rect 7064 23604 7070 23616
rect 7377 23613 7389 23616
rect 7423 23613 7435 23647
rect 7377 23607 7435 23613
rect 9582 23604 9588 23656
rect 9640 23644 9646 23656
rect 10520 23644 10548 23675
rect 11974 23672 11980 23684
rect 12032 23672 12038 23724
rect 12820 23721 12848 23752
rect 15194 23740 15200 23752
rect 15252 23740 15258 23792
rect 20622 23780 20628 23792
rect 15304 23752 20628 23780
rect 12805 23715 12863 23721
rect 12805 23681 12817 23715
rect 12851 23681 12863 23715
rect 12805 23675 12863 23681
rect 12894 23672 12900 23724
rect 12952 23712 12958 23724
rect 13061 23715 13119 23721
rect 13061 23712 13073 23715
rect 12952 23684 13073 23712
rect 12952 23672 12958 23684
rect 13061 23681 13073 23684
rect 13107 23681 13119 23715
rect 13061 23675 13119 23681
rect 13538 23672 13544 23724
rect 13596 23712 13602 23724
rect 15304 23712 15332 23752
rect 20622 23740 20628 23752
rect 20680 23740 20686 23792
rect 21266 23740 21272 23792
rect 21324 23780 21330 23792
rect 21726 23780 21732 23792
rect 21324 23752 21732 23780
rect 21324 23740 21330 23752
rect 21726 23740 21732 23752
rect 21784 23780 21790 23792
rect 22738 23780 22744 23792
rect 21784 23752 22744 23780
rect 21784 23740 21790 23752
rect 22738 23740 22744 23752
rect 22796 23740 22802 23792
rect 23106 23780 23112 23792
rect 22940 23752 23112 23780
rect 13596 23684 15332 23712
rect 13596 23672 13602 23684
rect 17954 23672 17960 23724
rect 18012 23712 18018 23724
rect 18049 23715 18107 23721
rect 18049 23712 18061 23715
rect 18012 23684 18061 23712
rect 18012 23672 18018 23684
rect 18049 23681 18061 23684
rect 18095 23681 18107 23715
rect 18049 23675 18107 23681
rect 21450 23672 21456 23724
rect 21508 23712 21514 23724
rect 22940 23721 22968 23752
rect 23106 23740 23112 23752
rect 23164 23740 23170 23792
rect 24302 23780 24308 23792
rect 24263 23752 24308 23780
rect 24302 23740 24308 23752
rect 24360 23740 24366 23792
rect 24964 23789 24992 23820
rect 27982 23808 27988 23860
rect 28040 23848 28046 23860
rect 28537 23851 28595 23857
rect 28537 23848 28549 23851
rect 28040 23820 28549 23848
rect 28040 23808 28046 23820
rect 28537 23817 28549 23820
rect 28583 23817 28595 23851
rect 32490 23848 32496 23860
rect 32451 23820 32496 23848
rect 28537 23811 28595 23817
rect 32490 23808 32496 23820
rect 32548 23848 32554 23860
rect 33134 23848 33140 23860
rect 32548 23820 33140 23848
rect 32548 23808 32554 23820
rect 33134 23808 33140 23820
rect 33192 23808 33198 23860
rect 39942 23808 39948 23860
rect 40000 23848 40006 23860
rect 40000 23820 40172 23848
rect 40000 23808 40006 23820
rect 24949 23783 25007 23789
rect 24949 23749 24961 23783
rect 24995 23780 25007 23783
rect 24995 23752 25820 23780
rect 24995 23749 25007 23752
rect 24949 23743 25007 23749
rect 22511 23715 22569 23721
rect 22511 23712 22523 23715
rect 21508 23684 22523 23712
rect 21508 23672 21514 23684
rect 22511 23681 22523 23684
rect 22557 23681 22569 23715
rect 22511 23675 22569 23681
rect 22649 23715 22707 23721
rect 22649 23681 22661 23715
rect 22695 23712 22707 23715
rect 22924 23715 22982 23721
rect 22695 23684 22876 23712
rect 22695 23681 22707 23684
rect 22649 23675 22707 23681
rect 22848 23644 22876 23684
rect 22924 23681 22936 23715
rect 22970 23681 22982 23715
rect 22924 23675 22982 23681
rect 23014 23672 23020 23724
rect 23072 23712 23078 23724
rect 24320 23712 24348 23740
rect 25409 23715 25467 23721
rect 25409 23712 25421 23715
rect 23072 23684 23117 23712
rect 24320 23684 25421 23712
rect 23072 23672 23078 23684
rect 25409 23681 25421 23684
rect 25455 23681 25467 23715
rect 25590 23712 25596 23724
rect 25551 23684 25596 23712
rect 25409 23675 25467 23681
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 25792 23721 25820 23752
rect 27614 23740 27620 23792
rect 27672 23780 27678 23792
rect 28902 23780 28908 23792
rect 27672 23752 28908 23780
rect 27672 23740 27678 23752
rect 28902 23740 28908 23752
rect 28960 23780 28966 23792
rect 28960 23752 29960 23780
rect 28960 23740 28966 23752
rect 25685 23715 25743 23721
rect 25685 23681 25697 23715
rect 25731 23681 25743 23715
rect 25685 23675 25743 23681
rect 25777 23715 25835 23721
rect 25777 23681 25789 23715
rect 25823 23681 25835 23715
rect 25777 23675 25835 23681
rect 24670 23644 24676 23656
rect 9640 23616 10548 23644
rect 22296 23616 22692 23644
rect 22848 23616 24676 23644
rect 9640 23604 9646 23616
rect 17770 23576 17776 23588
rect 14568 23548 17776 23576
rect 2590 23508 2596 23520
rect 2551 23480 2596 23508
rect 2590 23468 2596 23480
rect 2648 23468 2654 23520
rect 9677 23511 9735 23517
rect 9677 23477 9689 23511
rect 9723 23508 9735 23511
rect 10134 23508 10140 23520
rect 9723 23480 10140 23508
rect 9723 23477 9735 23480
rect 9677 23471 9735 23477
rect 10134 23468 10140 23480
rect 10192 23468 10198 23520
rect 11882 23468 11888 23520
rect 11940 23508 11946 23520
rect 14568 23508 14596 23548
rect 17770 23536 17776 23548
rect 17828 23536 17834 23588
rect 11940 23480 14596 23508
rect 11940 23468 11946 23480
rect 14642 23468 14648 23520
rect 14700 23508 14706 23520
rect 22296 23508 22324 23616
rect 22373 23579 22431 23585
rect 22373 23545 22385 23579
rect 22419 23576 22431 23579
rect 22554 23576 22560 23588
rect 22419 23548 22560 23576
rect 22419 23545 22431 23548
rect 22373 23539 22431 23545
rect 22554 23536 22560 23548
rect 22612 23536 22618 23588
rect 22664 23576 22692 23616
rect 24670 23604 24676 23616
rect 24728 23604 24734 23656
rect 23750 23576 23756 23588
rect 22664 23548 23756 23576
rect 23750 23536 23756 23548
rect 23808 23536 23814 23588
rect 24118 23536 24124 23588
rect 24176 23576 24182 23588
rect 24762 23576 24768 23588
rect 24176 23548 24768 23576
rect 24176 23536 24182 23548
rect 24762 23536 24768 23548
rect 24820 23576 24826 23588
rect 25700 23576 25728 23675
rect 29638 23672 29644 23724
rect 29696 23721 29702 23724
rect 29932 23721 29960 23752
rect 30650 23740 30656 23792
rect 30708 23780 30714 23792
rect 33502 23780 33508 23792
rect 30708 23752 33508 23780
rect 30708 23740 30714 23752
rect 33502 23740 33508 23752
rect 33560 23740 33566 23792
rect 33689 23783 33747 23789
rect 33689 23749 33701 23783
rect 33735 23780 33747 23783
rect 34330 23780 34336 23792
rect 33735 23752 34336 23780
rect 33735 23749 33747 23752
rect 33689 23743 33747 23749
rect 34330 23740 34336 23752
rect 34388 23740 34394 23792
rect 36081 23783 36139 23789
rect 36081 23749 36093 23783
rect 36127 23780 36139 23783
rect 36127 23752 38792 23780
rect 36127 23749 36139 23752
rect 36081 23743 36139 23749
rect 29696 23712 29708 23721
rect 29917 23715 29975 23721
rect 29696 23684 29741 23712
rect 29696 23675 29708 23684
rect 29917 23681 29929 23715
rect 29963 23681 29975 23715
rect 29917 23675 29975 23681
rect 33413 23715 33471 23721
rect 33413 23681 33425 23715
rect 33459 23712 33471 23715
rect 35526 23712 35532 23724
rect 33459 23684 35532 23712
rect 33459 23681 33471 23684
rect 33413 23675 33471 23681
rect 29696 23672 29702 23675
rect 35526 23672 35532 23684
rect 35584 23672 35590 23724
rect 35986 23712 35992 23724
rect 35947 23684 35992 23712
rect 35986 23672 35992 23684
rect 36044 23672 36050 23724
rect 36173 23715 36231 23721
rect 36173 23681 36185 23715
rect 36219 23712 36231 23715
rect 36262 23712 36268 23724
rect 36219 23684 36268 23712
rect 36219 23681 36231 23684
rect 36173 23675 36231 23681
rect 36262 23672 36268 23684
rect 36320 23672 36326 23724
rect 36357 23715 36415 23721
rect 36357 23681 36369 23715
rect 36403 23712 36415 23715
rect 36906 23712 36912 23724
rect 36403 23684 36912 23712
rect 36403 23681 36415 23684
rect 36357 23675 36415 23681
rect 36906 23672 36912 23684
rect 36964 23672 36970 23724
rect 33502 23644 33508 23656
rect 33463 23616 33508 23644
rect 33502 23604 33508 23616
rect 33560 23604 33566 23656
rect 24820 23548 25728 23576
rect 24820 23536 24826 23548
rect 30006 23536 30012 23588
rect 30064 23576 30070 23588
rect 33229 23579 33287 23585
rect 33229 23576 33241 23579
rect 30064 23548 33241 23576
rect 30064 23536 30070 23548
rect 33229 23545 33241 23548
rect 33275 23545 33287 23579
rect 33229 23539 33287 23545
rect 33318 23536 33324 23588
rect 33376 23576 33382 23588
rect 35805 23579 35863 23585
rect 35805 23576 35817 23579
rect 33376 23548 35817 23576
rect 33376 23536 33382 23548
rect 35805 23545 35817 23548
rect 35851 23545 35863 23579
rect 35805 23539 35863 23545
rect 14700 23480 22324 23508
rect 14700 23468 14706 23480
rect 25866 23468 25872 23520
rect 25924 23508 25930 23520
rect 26053 23511 26111 23517
rect 26053 23508 26065 23511
rect 25924 23480 26065 23508
rect 25924 23468 25930 23480
rect 26053 23477 26065 23480
rect 26099 23477 26111 23511
rect 33686 23508 33692 23520
rect 33647 23480 33692 23508
rect 26053 23471 26111 23477
rect 33686 23468 33692 23480
rect 33744 23468 33750 23520
rect 38764 23517 38792 23752
rect 40144 23721 40172 23820
rect 39873 23715 39931 23721
rect 39873 23681 39885 23715
rect 39919 23712 39931 23715
rect 40129 23715 40187 23721
rect 39919 23684 40080 23712
rect 39919 23681 39931 23684
rect 39873 23675 39931 23681
rect 40052 23644 40080 23684
rect 40129 23681 40141 23715
rect 40175 23681 40187 23715
rect 40862 23712 40868 23724
rect 40823 23684 40868 23712
rect 40129 23675 40187 23681
rect 40862 23672 40868 23684
rect 40920 23672 40926 23724
rect 40957 23715 41015 23721
rect 40957 23681 40969 23715
rect 41003 23681 41015 23715
rect 40957 23675 41015 23681
rect 41049 23715 41107 23721
rect 41049 23681 41061 23715
rect 41095 23712 41107 23715
rect 41138 23712 41144 23724
rect 41095 23684 41144 23712
rect 41095 23681 41107 23684
rect 41049 23675 41107 23681
rect 40589 23647 40647 23653
rect 40589 23644 40601 23647
rect 40052 23616 40601 23644
rect 40589 23613 40601 23616
rect 40635 23613 40647 23647
rect 40589 23607 40647 23613
rect 40678 23604 40684 23656
rect 40736 23644 40742 23656
rect 40972 23644 41000 23675
rect 41138 23672 41144 23684
rect 41196 23672 41202 23724
rect 41230 23672 41236 23724
rect 41288 23712 41294 23724
rect 41288 23684 41333 23712
rect 41288 23672 41294 23684
rect 40736 23616 41000 23644
rect 40736 23604 40742 23616
rect 38749 23511 38807 23517
rect 38749 23477 38761 23511
rect 38795 23508 38807 23511
rect 41046 23508 41052 23520
rect 38795 23480 41052 23508
rect 38795 23477 38807 23480
rect 38749 23471 38807 23477
rect 41046 23468 41052 23480
rect 41104 23468 41110 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 8113 23307 8171 23313
rect 8113 23273 8125 23307
rect 8159 23304 8171 23307
rect 11330 23304 11336 23316
rect 8159 23276 11336 23304
rect 8159 23273 8171 23276
rect 8113 23267 8171 23273
rect 2958 23196 2964 23248
rect 3016 23196 3022 23248
rect 2976 23168 3004 23196
rect 3786 23168 3792 23180
rect 2424 23140 3792 23168
rect 2424 23100 2452 23140
rect 3786 23128 3792 23140
rect 3844 23128 3850 23180
rect 7561 23171 7619 23177
rect 7561 23137 7573 23171
rect 7607 23168 7619 23171
rect 8128 23168 8156 23267
rect 11330 23264 11336 23276
rect 11388 23264 11394 23316
rect 11974 23264 11980 23316
rect 12032 23304 12038 23316
rect 12345 23307 12403 23313
rect 12345 23304 12357 23307
rect 12032 23276 12357 23304
rect 12032 23264 12038 23276
rect 12345 23273 12357 23276
rect 12391 23273 12403 23307
rect 16298 23304 16304 23316
rect 12345 23267 12403 23273
rect 14660 23276 16304 23304
rect 13814 23168 13820 23180
rect 7607 23140 8156 23168
rect 13004 23140 13820 23168
rect 7607 23137 7619 23140
rect 7561 23131 7619 23137
rect 2547 23103 2605 23109
rect 2547 23100 2559 23103
rect 2424 23072 2559 23100
rect 2547 23069 2559 23072
rect 2593 23069 2605 23103
rect 2682 23100 2688 23112
rect 2643 23072 2688 23100
rect 2547 23063 2605 23069
rect 2682 23060 2688 23072
rect 2740 23060 2746 23112
rect 2777 23103 2835 23109
rect 2777 23069 2789 23103
rect 2823 23069 2835 23103
rect 2777 23063 2835 23069
rect 2961 23103 3019 23109
rect 2961 23069 2973 23103
rect 3007 23100 3019 23103
rect 7282 23100 7288 23112
rect 3007 23072 7288 23100
rect 3007 23069 3019 23072
rect 2961 23063 3019 23069
rect 1578 22992 1584 23044
rect 1636 23032 1642 23044
rect 2792 23032 2820 23063
rect 7282 23060 7288 23072
rect 7340 23060 7346 23112
rect 10965 23103 11023 23109
rect 10965 23069 10977 23103
rect 11011 23100 11023 23103
rect 11054 23100 11060 23112
rect 11011 23072 11060 23100
rect 11011 23069 11023 23072
rect 10965 23063 11023 23069
rect 11054 23060 11060 23072
rect 11112 23060 11118 23112
rect 11232 23103 11290 23109
rect 11232 23069 11244 23103
rect 11278 23100 11290 23103
rect 11606 23100 11612 23112
rect 11278 23072 11612 23100
rect 11278 23069 11290 23072
rect 11232 23063 11290 23069
rect 11606 23060 11612 23072
rect 11664 23060 11670 23112
rect 12618 23060 12624 23112
rect 12676 23100 12682 23112
rect 13004 23109 13032 23140
rect 13814 23128 13820 23140
rect 13872 23168 13878 23180
rect 14093 23171 14151 23177
rect 14093 23168 14105 23171
rect 13872 23140 14105 23168
rect 13872 23128 13878 23140
rect 14093 23137 14105 23140
rect 14139 23168 14151 23171
rect 14366 23168 14372 23180
rect 14139 23140 14372 23168
rect 14139 23137 14151 23140
rect 14093 23131 14151 23137
rect 14366 23128 14372 23140
rect 14424 23128 14430 23180
rect 12805 23103 12863 23109
rect 12805 23100 12817 23103
rect 12676 23072 12817 23100
rect 12676 23060 12682 23072
rect 12805 23069 12817 23072
rect 12851 23069 12863 23103
rect 12805 23063 12863 23069
rect 12989 23103 13047 23109
rect 12989 23069 13001 23103
rect 13035 23069 13047 23103
rect 12989 23063 13047 23069
rect 13173 23103 13231 23109
rect 13173 23069 13185 23103
rect 13219 23100 13231 23103
rect 14660 23100 14688 23276
rect 16298 23264 16304 23276
rect 16356 23264 16362 23316
rect 16850 23304 16856 23316
rect 16811 23276 16856 23304
rect 16850 23264 16856 23276
rect 16908 23264 16914 23316
rect 20254 23264 20260 23316
rect 20312 23304 20318 23316
rect 20312 23276 20668 23304
rect 20312 23264 20318 23276
rect 15933 23239 15991 23245
rect 15933 23236 15945 23239
rect 15028 23208 15945 23236
rect 14826 23100 14832 23112
rect 13219 23072 14688 23100
rect 14787 23072 14832 23100
rect 13219 23069 13231 23072
rect 13173 23063 13231 23069
rect 1636 23004 2820 23032
rect 1636 22992 1642 23004
rect 11698 22992 11704 23044
rect 11756 23032 11762 23044
rect 13188 23032 13216 23063
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 14918 23060 14924 23112
rect 14976 23100 14982 23112
rect 15028 23109 15056 23208
rect 15933 23205 15945 23208
rect 15979 23236 15991 23239
rect 20640 23236 20668 23276
rect 21358 23264 21364 23316
rect 21416 23304 21422 23316
rect 21545 23307 21603 23313
rect 21545 23304 21557 23307
rect 21416 23276 21557 23304
rect 21416 23264 21422 23276
rect 21545 23273 21557 23276
rect 21591 23273 21603 23307
rect 22373 23307 22431 23313
rect 22373 23304 22385 23307
rect 21545 23267 21603 23273
rect 22066 23276 22385 23304
rect 22066 23236 22094 23276
rect 22373 23273 22385 23276
rect 22419 23273 22431 23307
rect 22373 23267 22431 23273
rect 22462 23264 22468 23316
rect 22520 23264 22526 23316
rect 29638 23304 29644 23316
rect 29551 23276 29644 23304
rect 29638 23264 29644 23276
rect 29696 23304 29702 23316
rect 29914 23304 29920 23316
rect 29696 23276 29920 23304
rect 29696 23264 29702 23276
rect 29914 23264 29920 23276
rect 29972 23264 29978 23316
rect 33870 23264 33876 23316
rect 33928 23304 33934 23316
rect 33928 23276 39344 23304
rect 33928 23264 33934 23276
rect 22480 23236 22508 23264
rect 39316 23245 39344 23276
rect 39758 23264 39764 23316
rect 39816 23304 39822 23316
rect 39945 23307 40003 23313
rect 39945 23304 39957 23307
rect 39816 23276 39957 23304
rect 39816 23264 39822 23276
rect 39945 23273 39957 23276
rect 39991 23273 40003 23307
rect 39945 23267 40003 23273
rect 40862 23264 40868 23316
rect 40920 23304 40926 23316
rect 41049 23307 41107 23313
rect 41049 23304 41061 23307
rect 40920 23276 41061 23304
rect 40920 23264 40926 23276
rect 41049 23273 41061 23276
rect 41095 23273 41107 23307
rect 41049 23267 41107 23273
rect 15979 23208 20576 23236
rect 20640 23208 22094 23236
rect 22388 23208 22508 23236
rect 39301 23239 39359 23245
rect 15979 23205 15991 23208
rect 15933 23199 15991 23205
rect 20548 23168 20576 23208
rect 22388 23168 22416 23208
rect 39301 23205 39313 23239
rect 39347 23236 39359 23239
rect 40770 23236 40776 23248
rect 39347 23208 40776 23236
rect 39347 23205 39359 23208
rect 39301 23199 39359 23205
rect 20548 23140 22416 23168
rect 22465 23171 22523 23177
rect 22465 23137 22477 23171
rect 22511 23168 22523 23171
rect 22511 23140 25360 23168
rect 22511 23137 22523 23140
rect 22465 23131 22523 23137
rect 15013 23103 15071 23109
rect 15013 23100 15025 23103
rect 14976 23072 15025 23100
rect 14976 23060 14982 23072
rect 15013 23069 15025 23072
rect 15059 23069 15071 23103
rect 15013 23063 15071 23069
rect 15197 23103 15255 23109
rect 15197 23069 15209 23103
rect 15243 23100 15255 23103
rect 16114 23100 16120 23112
rect 15243 23072 16120 23100
rect 15243 23069 15255 23072
rect 15197 23063 15255 23069
rect 16114 23060 16120 23072
rect 16172 23100 16178 23112
rect 22554 23100 22560 23112
rect 16172 23072 22094 23100
rect 22515 23072 22560 23100
rect 16172 23060 16178 23072
rect 11756 23004 13216 23032
rect 15105 23035 15163 23041
rect 11756 22992 11762 23004
rect 15105 23001 15117 23035
rect 15151 23032 15163 23035
rect 15838 23032 15844 23044
rect 15151 23004 15844 23032
rect 15151 23001 15163 23004
rect 15105 22995 15163 23001
rect 15838 22992 15844 23004
rect 15896 22992 15902 23044
rect 17954 22992 17960 23044
rect 18012 23032 18018 23044
rect 19245 23035 19303 23041
rect 19245 23032 19257 23035
rect 18012 23004 19257 23032
rect 18012 22992 18018 23004
rect 19245 23001 19257 23004
rect 19291 23001 19303 23035
rect 19245 22995 19303 23001
rect 19429 23035 19487 23041
rect 19429 23001 19441 23035
rect 19475 23032 19487 23035
rect 20070 23032 20076 23044
rect 19475 23004 20076 23032
rect 19475 23001 19487 23004
rect 19429 22995 19487 23001
rect 20070 22992 20076 23004
rect 20128 22992 20134 23044
rect 22066 23032 22094 23072
rect 22554 23060 22560 23072
rect 22612 23060 22618 23112
rect 22646 23032 22652 23044
rect 22066 23004 22652 23032
rect 22646 22992 22652 23004
rect 22704 22992 22710 23044
rect 24857 23035 24915 23041
rect 24857 23001 24869 23035
rect 24903 23001 24915 23035
rect 25332 23032 25360 23140
rect 25406 23128 25412 23180
rect 25464 23168 25470 23180
rect 25593 23171 25651 23177
rect 25593 23168 25605 23171
rect 25464 23140 25605 23168
rect 25464 23128 25470 23140
rect 25593 23137 25605 23140
rect 25639 23137 25651 23171
rect 25593 23131 25651 23137
rect 34054 23128 34060 23180
rect 34112 23168 34118 23180
rect 35710 23168 35716 23180
rect 34112 23140 35716 23168
rect 34112 23128 34118 23140
rect 35710 23128 35716 23140
rect 35768 23168 35774 23180
rect 35897 23171 35955 23177
rect 35897 23168 35909 23171
rect 35768 23140 35909 23168
rect 35768 23128 35774 23140
rect 35897 23137 35909 23140
rect 35943 23137 35955 23171
rect 35897 23131 35955 23137
rect 25866 23109 25872 23112
rect 25860 23100 25872 23109
rect 25827 23072 25872 23100
rect 25860 23063 25872 23072
rect 25866 23060 25872 23063
rect 25924 23060 25930 23112
rect 26234 23060 26240 23112
rect 26292 23100 26298 23112
rect 34238 23100 34244 23112
rect 26292 23072 34244 23100
rect 26292 23060 26298 23072
rect 34238 23060 34244 23072
rect 34296 23060 34302 23112
rect 40144 23100 40172 23208
rect 40770 23196 40776 23208
rect 40828 23196 40834 23248
rect 40221 23103 40279 23109
rect 40221 23100 40233 23103
rect 40144 23072 40233 23100
rect 40221 23069 40233 23072
rect 40267 23069 40279 23103
rect 40221 23063 40279 23069
rect 40313 23103 40371 23109
rect 40313 23069 40325 23103
rect 40359 23069 40371 23103
rect 40313 23063 40371 23069
rect 28810 23032 28816 23044
rect 25332 23004 28816 23032
rect 24857 22995 24915 23001
rect 2314 22964 2320 22976
rect 2275 22936 2320 22964
rect 2314 22924 2320 22936
rect 2372 22924 2378 22976
rect 3786 22964 3792 22976
rect 3747 22936 3792 22964
rect 3786 22924 3792 22936
rect 3844 22924 3850 22976
rect 9858 22924 9864 22976
rect 9916 22964 9922 22976
rect 14734 22964 14740 22976
rect 9916 22936 14740 22964
rect 9916 22924 9922 22936
rect 14734 22924 14740 22936
rect 14792 22924 14798 22976
rect 15378 22964 15384 22976
rect 15339 22936 15384 22964
rect 15378 22924 15384 22936
rect 15436 22924 15442 22976
rect 19334 22924 19340 22976
rect 19392 22964 19398 22976
rect 19613 22967 19671 22973
rect 19613 22964 19625 22967
rect 19392 22936 19625 22964
rect 19392 22924 19398 22936
rect 19613 22933 19625 22936
rect 19659 22933 19671 22967
rect 19613 22927 19671 22933
rect 22189 22967 22247 22973
rect 22189 22933 22201 22967
rect 22235 22964 22247 22967
rect 22462 22964 22468 22976
rect 22235 22936 22468 22964
rect 22235 22933 22247 22936
rect 22189 22927 22247 22933
rect 22462 22924 22468 22936
rect 22520 22924 22526 22976
rect 23750 22964 23756 22976
rect 23711 22936 23756 22964
rect 23750 22924 23756 22936
rect 23808 22964 23814 22976
rect 24872 22964 24900 22995
rect 28810 22992 28816 23004
rect 28868 22992 28874 23044
rect 31849 23035 31907 23041
rect 31849 23001 31861 23035
rect 31895 23032 31907 23035
rect 31938 23032 31944 23044
rect 31895 23004 31944 23032
rect 31895 23001 31907 23004
rect 31849 22995 31907 23001
rect 31938 22992 31944 23004
rect 31996 22992 32002 23044
rect 32030 22992 32036 23044
rect 32088 23032 32094 23044
rect 32088 23004 32720 23032
rect 32088 22992 32094 23004
rect 23808 22936 24900 22964
rect 24949 22967 25007 22973
rect 23808 22924 23814 22936
rect 24949 22933 24961 22967
rect 24995 22964 25007 22967
rect 26326 22964 26332 22976
rect 24995 22936 26332 22964
rect 24995 22933 25007 22936
rect 24949 22927 25007 22933
rect 26326 22924 26332 22936
rect 26384 22924 26390 22976
rect 26973 22967 27031 22973
rect 26973 22933 26985 22967
rect 27019 22964 27031 22967
rect 27338 22964 27344 22976
rect 27019 22936 27344 22964
rect 27019 22933 27031 22936
rect 26973 22927 27031 22933
rect 27338 22924 27344 22936
rect 27396 22924 27402 22976
rect 32214 22964 32220 22976
rect 32175 22936 32220 22964
rect 32214 22924 32220 22936
rect 32272 22924 32278 22976
rect 32692 22973 32720 23004
rect 33226 22992 33232 23044
rect 33284 23032 33290 23044
rect 36170 23041 36176 23044
rect 33790 23035 33848 23041
rect 33790 23032 33802 23035
rect 33284 23004 33802 23032
rect 33284 22992 33290 23004
rect 33790 23001 33802 23004
rect 33836 23001 33848 23035
rect 33790 22995 33848 23001
rect 36164 22995 36176 23041
rect 36228 23032 36234 23044
rect 40328 23032 40356 23063
rect 40402 23060 40408 23112
rect 40460 23100 40466 23112
rect 40589 23103 40647 23109
rect 40460 23072 40505 23100
rect 40460 23060 40466 23072
rect 40589 23069 40601 23103
rect 40635 23100 40647 23103
rect 41138 23100 41144 23112
rect 40635 23072 41144 23100
rect 40635 23069 40647 23072
rect 40589 23063 40647 23069
rect 41138 23060 41144 23072
rect 41196 23060 41202 23112
rect 40678 23032 40684 23044
rect 36228 23004 36264 23032
rect 40328 23004 40684 23032
rect 36170 22992 36176 22995
rect 36228 22992 36234 23004
rect 40420 22976 40448 23004
rect 40678 22992 40684 23004
rect 40736 22992 40742 23044
rect 32677 22967 32735 22973
rect 32677 22933 32689 22967
rect 32723 22933 32735 22967
rect 32677 22927 32735 22933
rect 35437 22967 35495 22973
rect 35437 22933 35449 22967
rect 35483 22964 35495 22967
rect 36722 22964 36728 22976
rect 35483 22936 36728 22964
rect 35483 22933 35495 22936
rect 35437 22927 35495 22933
rect 36722 22924 36728 22936
rect 36780 22924 36786 22976
rect 37274 22964 37280 22976
rect 37235 22936 37280 22964
rect 37274 22924 37280 22936
rect 37332 22924 37338 22976
rect 40402 22924 40408 22976
rect 40460 22924 40466 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1578 22760 1584 22772
rect 1539 22732 1584 22760
rect 1578 22720 1584 22732
rect 1636 22720 1642 22772
rect 5994 22760 6000 22772
rect 5460 22732 6000 22760
rect 2314 22652 2320 22704
rect 2372 22692 2378 22704
rect 2654 22695 2712 22701
rect 2654 22692 2666 22695
rect 2372 22664 2666 22692
rect 2372 22652 2378 22664
rect 2654 22661 2666 22664
rect 2700 22661 2712 22695
rect 2654 22655 2712 22661
rect 4433 22695 4491 22701
rect 4433 22661 4445 22695
rect 4479 22692 4491 22695
rect 5166 22692 5172 22704
rect 4479 22664 5172 22692
rect 4479 22661 4491 22664
rect 4433 22655 4491 22661
rect 5166 22652 5172 22664
rect 5224 22652 5230 22704
rect 5460 22701 5488 22732
rect 5994 22720 6000 22732
rect 6052 22760 6058 22772
rect 8481 22763 8539 22769
rect 8481 22760 8493 22763
rect 6052 22732 8493 22760
rect 6052 22720 6058 22732
rect 8481 22729 8493 22732
rect 8527 22729 8539 22763
rect 8481 22723 8539 22729
rect 9677 22763 9735 22769
rect 9677 22729 9689 22763
rect 9723 22760 9735 22763
rect 10410 22760 10416 22772
rect 9723 22732 10416 22760
rect 9723 22729 9735 22732
rect 9677 22723 9735 22729
rect 10410 22720 10416 22732
rect 10468 22760 10474 22772
rect 15565 22763 15623 22769
rect 15565 22760 15577 22763
rect 10468 22732 12434 22760
rect 10468 22720 10474 22732
rect 5445 22695 5503 22701
rect 5445 22661 5457 22695
rect 5491 22661 5503 22695
rect 5445 22655 5503 22661
rect 5629 22695 5687 22701
rect 5629 22661 5641 22695
rect 5675 22692 5687 22695
rect 11793 22695 11851 22701
rect 5675 22664 8064 22692
rect 5675 22661 5687 22664
rect 5629 22655 5687 22661
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22593 1823 22627
rect 1765 22587 1823 22593
rect 1949 22627 2007 22633
rect 1949 22593 1961 22627
rect 1995 22593 2007 22627
rect 2406 22624 2412 22636
rect 2367 22596 2412 22624
rect 1949 22587 2007 22593
rect 1780 22420 1808 22587
rect 1964 22556 1992 22587
rect 2406 22584 2412 22596
rect 2464 22584 2470 22636
rect 4617 22627 4675 22633
rect 4617 22624 4629 22627
rect 2516 22596 4629 22624
rect 2222 22556 2228 22568
rect 1964 22528 2228 22556
rect 2222 22516 2228 22528
rect 2280 22556 2286 22568
rect 2516 22556 2544 22596
rect 4617 22593 4629 22596
rect 4663 22624 4675 22627
rect 5460 22624 5488 22655
rect 4663 22596 5488 22624
rect 4663 22593 4675 22596
rect 4617 22587 4675 22593
rect 6362 22584 6368 22636
rect 6420 22624 6426 22636
rect 6914 22633 6920 22636
rect 6641 22627 6699 22633
rect 6641 22624 6653 22627
rect 6420 22596 6653 22624
rect 6420 22584 6426 22596
rect 6641 22593 6653 22596
rect 6687 22593 6699 22627
rect 6641 22587 6699 22593
rect 6908 22587 6920 22633
rect 6972 22624 6978 22636
rect 6972 22596 7008 22624
rect 6914 22584 6920 22587
rect 6972 22584 6978 22596
rect 2280 22528 2544 22556
rect 2280 22516 2286 22528
rect 8036 22497 8064 22664
rect 11793 22661 11805 22695
rect 11839 22692 11851 22695
rect 11974 22692 11980 22704
rect 11839 22664 11980 22692
rect 11839 22661 11851 22664
rect 11793 22655 11851 22661
rect 11974 22652 11980 22664
rect 12032 22652 12038 22704
rect 8662 22624 8668 22636
rect 8623 22596 8668 22624
rect 8662 22584 8668 22596
rect 8720 22584 8726 22636
rect 9214 22584 9220 22636
rect 9272 22624 9278 22636
rect 9585 22627 9643 22633
rect 9585 22624 9597 22627
rect 9272 22596 9597 22624
rect 9272 22584 9278 22596
rect 9585 22593 9597 22596
rect 9631 22624 9643 22627
rect 10318 22624 10324 22636
rect 9631 22596 10324 22624
rect 9631 22593 9643 22596
rect 9585 22587 9643 22593
rect 10318 22584 10324 22596
rect 10376 22584 10382 22636
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 10428 22596 11529 22624
rect 8110 22516 8116 22568
rect 8168 22556 8174 22568
rect 10428 22556 10456 22596
rect 11517 22593 11529 22596
rect 11563 22593 11575 22627
rect 11698 22624 11704 22636
rect 11659 22596 11704 22624
rect 11517 22587 11575 22593
rect 11698 22584 11704 22596
rect 11756 22584 11762 22636
rect 11882 22584 11888 22636
rect 11940 22624 11946 22636
rect 11940 22596 12033 22624
rect 11940 22584 11946 22596
rect 8168 22528 10456 22556
rect 8168 22516 8174 22528
rect 11054 22516 11060 22568
rect 11112 22556 11118 22568
rect 11900 22556 11928 22584
rect 11112 22528 11928 22556
rect 12406 22556 12434 22732
rect 14108 22732 15577 22760
rect 14108 22624 14136 22732
rect 15565 22729 15577 22732
rect 15611 22760 15623 22763
rect 16114 22760 16120 22772
rect 15611 22732 16120 22760
rect 15611 22729 15623 22732
rect 15565 22723 15623 22729
rect 16114 22720 16120 22732
rect 16172 22720 16178 22772
rect 18049 22763 18107 22769
rect 18049 22760 18061 22763
rect 17926 22732 18061 22760
rect 14182 22652 14188 22704
rect 14240 22692 14246 22704
rect 14369 22695 14427 22701
rect 14369 22692 14381 22695
rect 14240 22664 14381 22692
rect 14240 22652 14246 22664
rect 14369 22661 14381 22664
rect 14415 22661 14427 22695
rect 14369 22655 14427 22661
rect 14461 22695 14519 22701
rect 14461 22661 14473 22695
rect 14507 22692 14519 22695
rect 14918 22692 14924 22704
rect 14507 22664 14924 22692
rect 14507 22661 14519 22664
rect 14461 22655 14519 22661
rect 14918 22652 14924 22664
rect 14976 22652 14982 22704
rect 17926 22692 17954 22732
rect 18049 22729 18061 22732
rect 18095 22760 18107 22763
rect 18598 22760 18604 22772
rect 18095 22732 18604 22760
rect 18095 22729 18107 22732
rect 18049 22723 18107 22729
rect 18598 22720 18604 22732
rect 18656 22760 18662 22772
rect 18782 22760 18788 22772
rect 18656 22732 18788 22760
rect 18656 22720 18662 22732
rect 18782 22720 18788 22732
rect 18840 22720 18846 22772
rect 20162 22720 20168 22772
rect 20220 22760 20226 22772
rect 23750 22760 23756 22772
rect 20220 22732 23756 22760
rect 20220 22720 20226 22732
rect 23750 22720 23756 22732
rect 23808 22720 23814 22772
rect 24946 22720 24952 22772
rect 25004 22760 25010 22772
rect 25317 22763 25375 22769
rect 25317 22760 25329 22763
rect 25004 22732 25329 22760
rect 25004 22720 25010 22732
rect 25317 22729 25329 22732
rect 25363 22729 25375 22763
rect 25317 22723 25375 22729
rect 23934 22692 23940 22704
rect 16408 22664 17954 22692
rect 20732 22664 23940 22692
rect 14277 22627 14335 22633
rect 14277 22624 14289 22627
rect 14108 22596 14289 22624
rect 14277 22593 14289 22596
rect 14323 22593 14335 22627
rect 14642 22624 14648 22636
rect 14603 22596 14648 22624
rect 14277 22587 14335 22593
rect 14642 22584 14648 22596
rect 14700 22584 14706 22636
rect 16408 22556 16436 22664
rect 16482 22584 16488 22636
rect 16540 22624 16546 22636
rect 18693 22627 18751 22633
rect 18693 22624 18705 22627
rect 16540 22596 18705 22624
rect 16540 22584 16546 22596
rect 18693 22593 18705 22596
rect 18739 22593 18751 22627
rect 18693 22587 18751 22593
rect 18782 22584 18788 22636
rect 18840 22624 18846 22636
rect 20732 22633 20760 22664
rect 23934 22652 23940 22664
rect 23992 22652 23998 22704
rect 18949 22627 19007 22633
rect 18949 22624 18961 22627
rect 18840 22596 18961 22624
rect 18840 22584 18846 22596
rect 18949 22593 18961 22596
rect 18995 22593 19007 22627
rect 18949 22587 19007 22593
rect 20717 22627 20775 22633
rect 20717 22593 20729 22627
rect 20763 22593 20775 22627
rect 20898 22624 20904 22636
rect 20859 22596 20904 22624
rect 20717 22587 20775 22593
rect 20898 22584 20904 22596
rect 20956 22584 20962 22636
rect 22186 22624 22192 22636
rect 22147 22596 22192 22624
rect 22186 22584 22192 22596
rect 22244 22584 22250 22636
rect 24118 22624 24124 22636
rect 24079 22596 24124 22624
rect 24118 22584 24124 22596
rect 24176 22584 24182 22636
rect 24762 22584 24768 22636
rect 24820 22624 24826 22636
rect 25133 22627 25191 22633
rect 25133 22624 25145 22627
rect 24820 22596 25145 22624
rect 24820 22584 24826 22596
rect 25133 22593 25145 22596
rect 25179 22593 25191 22627
rect 25332 22624 25360 22723
rect 25590 22720 25596 22772
rect 25648 22760 25654 22772
rect 25961 22763 26019 22769
rect 25961 22760 25973 22763
rect 25648 22732 25973 22760
rect 25648 22720 25654 22732
rect 25961 22729 25973 22732
rect 26007 22729 26019 22763
rect 27798 22760 27804 22772
rect 25961 22723 26019 22729
rect 26068 22732 27804 22760
rect 25866 22652 25872 22704
rect 25924 22692 25930 22704
rect 26068 22692 26096 22732
rect 27798 22720 27804 22732
rect 27856 22760 27862 22772
rect 27856 22732 27936 22760
rect 27856 22720 27862 22732
rect 25924 22664 26096 22692
rect 26145 22695 26203 22701
rect 25924 22652 25930 22664
rect 26145 22661 26157 22695
rect 26191 22692 26203 22695
rect 27338 22692 27344 22704
rect 26191 22664 27344 22692
rect 26191 22661 26203 22664
rect 26145 22655 26203 22661
rect 27338 22652 27344 22664
rect 27396 22652 27402 22704
rect 27908 22701 27936 22732
rect 33042 22720 33048 22772
rect 33100 22720 33106 22772
rect 33226 22760 33232 22772
rect 33187 22732 33232 22760
rect 33226 22720 33232 22732
rect 33284 22720 33290 22772
rect 33686 22760 33692 22772
rect 33647 22732 33692 22760
rect 33686 22720 33692 22732
rect 33744 22720 33750 22772
rect 36081 22763 36139 22769
rect 36081 22729 36093 22763
rect 36127 22760 36139 22763
rect 36170 22760 36176 22772
rect 36127 22732 36176 22760
rect 36127 22729 36139 22732
rect 36081 22723 36139 22729
rect 36170 22720 36176 22732
rect 36228 22720 36234 22772
rect 27893 22695 27951 22701
rect 27893 22661 27905 22695
rect 27939 22661 27951 22695
rect 27893 22655 27951 22661
rect 31205 22695 31263 22701
rect 31205 22661 31217 22695
rect 31251 22692 31263 22695
rect 32122 22692 32128 22704
rect 31251 22664 32128 22692
rect 31251 22661 31263 22664
rect 31205 22655 31263 22661
rect 32122 22652 32128 22664
rect 32180 22652 32186 22704
rect 32214 22652 32220 22704
rect 32272 22692 32278 22704
rect 33060 22692 33088 22720
rect 34054 22692 34060 22704
rect 32272 22664 32720 22692
rect 33060 22664 33916 22692
rect 34015 22664 34060 22692
rect 32272 22652 32278 22664
rect 26329 22627 26387 22633
rect 26329 22624 26341 22627
rect 25332 22596 26341 22624
rect 25133 22587 25191 22593
rect 26329 22593 26341 22596
rect 26375 22593 26387 22627
rect 26329 22587 26387 22593
rect 28077 22627 28135 22633
rect 28077 22593 28089 22627
rect 28123 22593 28135 22627
rect 28077 22587 28135 22593
rect 16666 22556 16672 22568
rect 12406 22528 16436 22556
rect 16627 22528 16672 22556
rect 11112 22516 11118 22528
rect 16666 22516 16672 22528
rect 16724 22516 16730 22568
rect 16945 22559 17003 22565
rect 16945 22525 16957 22559
rect 16991 22525 17003 22559
rect 16945 22519 17003 22525
rect 22097 22559 22155 22565
rect 22097 22525 22109 22559
rect 22143 22525 22155 22559
rect 22097 22519 22155 22525
rect 3789 22491 3847 22497
rect 3789 22457 3801 22491
rect 3835 22488 3847 22491
rect 8021 22491 8079 22497
rect 3835 22460 6500 22488
rect 3835 22457 3847 22460
rect 3789 22451 3847 22457
rect 3804 22420 3832 22451
rect 1780 22392 3832 22420
rect 4249 22423 4307 22429
rect 4249 22389 4261 22423
rect 4295 22420 4307 22423
rect 4614 22420 4620 22432
rect 4295 22392 4620 22420
rect 4295 22389 4307 22392
rect 4249 22383 4307 22389
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 5813 22423 5871 22429
rect 5813 22389 5825 22423
rect 5859 22420 5871 22423
rect 6362 22420 6368 22432
rect 5859 22392 6368 22420
rect 5859 22389 5871 22392
rect 5813 22383 5871 22389
rect 6362 22380 6368 22392
rect 6420 22380 6426 22432
rect 6472 22420 6500 22460
rect 8021 22457 8033 22491
rect 8067 22488 8079 22491
rect 14826 22488 14832 22500
rect 8067 22460 14832 22488
rect 8067 22457 8079 22460
rect 8021 22451 8079 22457
rect 14826 22448 14832 22460
rect 14884 22448 14890 22500
rect 16298 22448 16304 22500
rect 16356 22488 16362 22500
rect 16960 22488 16988 22519
rect 20070 22488 20076 22500
rect 16356 22460 16988 22488
rect 19983 22460 20076 22488
rect 16356 22448 16362 22460
rect 20070 22448 20076 22460
rect 20128 22488 20134 22500
rect 20622 22488 20628 22500
rect 20128 22460 20628 22488
rect 20128 22448 20134 22460
rect 20622 22448 20628 22460
rect 20680 22448 20686 22500
rect 21358 22448 21364 22500
rect 21416 22488 21422 22500
rect 22112 22488 22140 22519
rect 23566 22516 23572 22568
rect 23624 22556 23630 22568
rect 23845 22559 23903 22565
rect 23845 22556 23857 22559
rect 23624 22528 23857 22556
rect 23624 22516 23630 22528
rect 23845 22525 23857 22528
rect 23891 22525 23903 22559
rect 23845 22519 23903 22525
rect 24670 22516 24676 22568
rect 24728 22556 24734 22568
rect 28092 22556 28120 22587
rect 28166 22584 28172 22636
rect 28224 22624 28230 22636
rect 31021 22627 31079 22633
rect 31021 22624 31033 22627
rect 28224 22596 31033 22624
rect 28224 22584 28230 22596
rect 31021 22593 31033 22596
rect 31067 22593 31079 22627
rect 31021 22587 31079 22593
rect 31297 22627 31355 22633
rect 31297 22593 31309 22627
rect 31343 22593 31355 22627
rect 31297 22587 31355 22593
rect 28902 22556 28908 22568
rect 24728 22528 28908 22556
rect 24728 22516 24734 22528
rect 28902 22516 28908 22528
rect 28960 22516 28966 22568
rect 23658 22488 23664 22500
rect 21416 22460 22048 22488
rect 22112 22460 23664 22488
rect 21416 22448 21422 22460
rect 8386 22420 8392 22432
rect 6472 22392 8392 22420
rect 8386 22380 8392 22392
rect 8444 22380 8450 22432
rect 10318 22420 10324 22432
rect 10279 22392 10324 22420
rect 10318 22380 10324 22392
rect 10376 22380 10382 22432
rect 12069 22423 12127 22429
rect 12069 22389 12081 22423
rect 12115 22420 12127 22423
rect 12894 22420 12900 22432
rect 12115 22392 12900 22420
rect 12115 22389 12127 22392
rect 12069 22383 12127 22389
rect 12894 22380 12900 22392
rect 12952 22380 12958 22432
rect 14093 22423 14151 22429
rect 14093 22389 14105 22423
rect 14139 22420 14151 22423
rect 14458 22420 14464 22432
rect 14139 22392 14464 22420
rect 14139 22389 14151 22392
rect 14093 22383 14151 22389
rect 14458 22380 14464 22392
rect 14516 22380 14522 22432
rect 14734 22380 14740 22432
rect 14792 22420 14798 22432
rect 20533 22423 20591 22429
rect 20533 22420 20545 22423
rect 14792 22392 20545 22420
rect 14792 22380 14798 22392
rect 20533 22389 20545 22392
rect 20579 22389 20591 22423
rect 20533 22383 20591 22389
rect 20901 22423 20959 22429
rect 20901 22389 20913 22423
rect 20947 22420 20959 22423
rect 21082 22420 21088 22432
rect 20947 22392 21088 22420
rect 20947 22389 20959 22392
rect 20901 22383 20959 22389
rect 21082 22380 21088 22392
rect 21140 22380 21146 22432
rect 21634 22380 21640 22432
rect 21692 22420 21698 22432
rect 22020 22429 22048 22460
rect 23658 22448 23664 22460
rect 23716 22448 23722 22500
rect 31312 22488 31340 22587
rect 31386 22584 31392 22636
rect 31444 22624 31450 22636
rect 31444 22596 31489 22624
rect 31444 22584 31450 22596
rect 32306 22584 32312 22636
rect 32364 22624 32370 22636
rect 32585 22627 32643 22633
rect 32585 22624 32597 22627
rect 32364 22596 32597 22624
rect 32364 22584 32370 22596
rect 32585 22593 32597 22596
rect 32631 22593 32643 22627
rect 32692 22627 32720 22664
rect 32748 22630 32806 22636
rect 32748 22627 32760 22630
rect 32692 22599 32760 22627
rect 32585 22587 32643 22593
rect 32748 22596 32760 22599
rect 32794 22596 32806 22630
rect 32748 22590 32806 22596
rect 32858 22584 32864 22636
rect 32916 22624 32922 22636
rect 32999 22627 33057 22633
rect 32916 22596 32961 22624
rect 32916 22584 32922 22596
rect 32999 22593 33011 22627
rect 33045 22624 33057 22627
rect 33134 22624 33140 22636
rect 33045 22596 33140 22624
rect 33045 22593 33057 22596
rect 32999 22587 33057 22593
rect 33134 22584 33140 22596
rect 33192 22584 33198 22636
rect 33888 22633 33916 22664
rect 34054 22652 34060 22664
rect 34112 22652 34118 22704
rect 35345 22695 35403 22701
rect 35345 22661 35357 22695
rect 35391 22692 35403 22695
rect 37274 22692 37280 22704
rect 35391 22664 37280 22692
rect 35391 22661 35403 22664
rect 35345 22655 35403 22661
rect 37274 22652 37280 22664
rect 37332 22692 37338 22704
rect 37461 22695 37519 22701
rect 37461 22692 37473 22695
rect 37332 22664 37473 22692
rect 37332 22652 37338 22664
rect 37461 22661 37473 22664
rect 37507 22661 37519 22695
rect 37461 22655 37519 22661
rect 38562 22652 38568 22704
rect 38620 22692 38626 22704
rect 39669 22695 39727 22701
rect 39669 22692 39681 22695
rect 38620 22664 39681 22692
rect 38620 22652 38626 22664
rect 39669 22661 39681 22664
rect 39715 22661 39727 22695
rect 39669 22655 39727 22661
rect 33873 22627 33931 22633
rect 33873 22593 33885 22627
rect 33919 22593 33931 22627
rect 33873 22587 33931 22593
rect 33962 22584 33968 22636
rect 34020 22624 34026 22636
rect 34238 22624 34244 22636
rect 34020 22596 34065 22624
rect 34199 22596 34244 22624
rect 34020 22584 34026 22596
rect 34238 22584 34244 22596
rect 34296 22584 34302 22636
rect 35253 22627 35311 22633
rect 35253 22593 35265 22627
rect 35299 22624 35311 22627
rect 35437 22627 35495 22633
rect 35299 22596 35388 22624
rect 35299 22593 35311 22596
rect 35253 22587 35311 22593
rect 33778 22488 33784 22500
rect 31312 22460 33784 22488
rect 33778 22448 33784 22460
rect 33836 22448 33842 22500
rect 21821 22423 21879 22429
rect 21821 22420 21833 22423
rect 21692 22392 21833 22420
rect 21692 22380 21698 22392
rect 21821 22389 21833 22392
rect 21867 22389 21879 22423
rect 21821 22383 21879 22389
rect 22005 22423 22063 22429
rect 22005 22389 22017 22423
rect 22051 22389 22063 22423
rect 22005 22383 22063 22389
rect 22554 22380 22560 22432
rect 22612 22420 22618 22432
rect 22833 22423 22891 22429
rect 22833 22420 22845 22423
rect 22612 22392 22845 22420
rect 22612 22380 22618 22392
rect 22833 22389 22845 22392
rect 22879 22389 22891 22423
rect 22833 22383 22891 22389
rect 28074 22380 28080 22432
rect 28132 22420 28138 22432
rect 28261 22423 28319 22429
rect 28261 22420 28273 22423
rect 28132 22392 28273 22420
rect 28132 22380 28138 22392
rect 28261 22389 28273 22392
rect 28307 22389 28319 22423
rect 28261 22383 28319 22389
rect 31573 22423 31631 22429
rect 31573 22389 31585 22423
rect 31619 22420 31631 22423
rect 32950 22420 32956 22432
rect 31619 22392 32956 22420
rect 31619 22389 31631 22392
rect 31573 22383 31631 22389
rect 32950 22380 32956 22392
rect 33008 22380 33014 22432
rect 33134 22380 33140 22432
rect 33192 22420 33198 22432
rect 35069 22423 35127 22429
rect 35069 22420 35081 22423
rect 33192 22392 35081 22420
rect 33192 22380 33198 22392
rect 35069 22389 35081 22392
rect 35115 22389 35127 22423
rect 35360 22420 35388 22596
rect 35437 22593 35449 22627
rect 35483 22593 35495 22627
rect 35618 22624 35624 22636
rect 35579 22596 35624 22624
rect 35437 22587 35495 22593
rect 35452 22488 35480 22587
rect 35618 22584 35624 22596
rect 35676 22584 35682 22636
rect 36354 22624 36360 22636
rect 36315 22596 36360 22624
rect 36354 22584 36360 22596
rect 36412 22584 36418 22636
rect 36449 22627 36507 22633
rect 36449 22593 36461 22627
rect 36495 22593 36507 22627
rect 36449 22587 36507 22593
rect 36541 22627 36599 22633
rect 36541 22593 36553 22627
rect 36587 22593 36599 22627
rect 36722 22624 36728 22636
rect 36683 22596 36728 22624
rect 36541 22587 36599 22593
rect 36262 22488 36268 22500
rect 35452 22460 36268 22488
rect 36262 22448 36268 22460
rect 36320 22448 36326 22500
rect 36464 22488 36492 22587
rect 36556 22556 36584 22587
rect 36722 22584 36728 22596
rect 36780 22624 36786 22636
rect 36998 22624 37004 22636
rect 36780 22596 37004 22624
rect 36780 22584 36786 22596
rect 36998 22584 37004 22596
rect 37056 22584 37062 22636
rect 37645 22627 37703 22633
rect 37645 22593 37657 22627
rect 37691 22593 37703 22627
rect 37645 22587 37703 22593
rect 37277 22559 37335 22565
rect 37277 22556 37289 22559
rect 36556 22528 37289 22556
rect 37277 22525 37289 22528
rect 37323 22525 37335 22559
rect 37660 22556 37688 22587
rect 38470 22584 38476 22636
rect 38528 22624 38534 22636
rect 38930 22624 38936 22636
rect 38528 22596 38936 22624
rect 38528 22584 38534 22596
rect 38930 22584 38936 22596
rect 38988 22624 38994 22636
rect 39485 22627 39543 22633
rect 39485 22624 39497 22627
rect 38988 22596 39497 22624
rect 38988 22584 38994 22596
rect 39485 22593 39497 22596
rect 39531 22593 39543 22627
rect 39485 22587 39543 22593
rect 39758 22556 39764 22568
rect 37660 22528 39764 22556
rect 37277 22519 37335 22525
rect 39758 22516 39764 22528
rect 39816 22516 39822 22568
rect 40402 22488 40408 22500
rect 36464 22460 40408 22488
rect 40402 22448 40408 22460
rect 40460 22448 40466 22500
rect 58158 22488 58164 22500
rect 58119 22460 58164 22488
rect 58158 22448 58164 22460
rect 58216 22448 58222 22500
rect 35986 22420 35992 22432
rect 35360 22392 35992 22420
rect 35069 22383 35127 22389
rect 35986 22380 35992 22392
rect 36044 22380 36050 22432
rect 39853 22423 39911 22429
rect 39853 22389 39865 22423
rect 39899 22420 39911 22423
rect 40310 22420 40316 22432
rect 39899 22392 40316 22420
rect 39899 22389 39911 22392
rect 39853 22383 39911 22389
rect 40310 22380 40316 22392
rect 40368 22380 40374 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 3234 22216 3240 22228
rect 3147 22188 3240 22216
rect 3234 22176 3240 22188
rect 3292 22216 3298 22228
rect 8110 22216 8116 22228
rect 3292 22188 8116 22216
rect 3292 22176 3298 22188
rect 8110 22176 8116 22188
rect 8168 22176 8174 22228
rect 8662 22176 8668 22228
rect 8720 22216 8726 22228
rect 8941 22219 8999 22225
rect 8941 22216 8953 22219
rect 8720 22188 8953 22216
rect 8720 22176 8726 22188
rect 8941 22185 8953 22188
rect 8987 22185 8999 22219
rect 14918 22216 14924 22228
rect 14879 22188 14924 22216
rect 8941 22179 8999 22185
rect 6086 22040 6092 22092
rect 6144 22080 6150 22092
rect 6825 22083 6883 22089
rect 6144 22052 6776 22080
rect 6144 22040 6150 22052
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 2866 22012 2872 22024
rect 1903 21984 2872 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 2866 21972 2872 21984
rect 2924 22012 2930 22024
rect 3789 22015 3847 22021
rect 3789 22012 3801 22015
rect 2924 21984 3801 22012
rect 2924 21972 2930 21984
rect 3789 21981 3801 21984
rect 3835 21981 3847 22015
rect 3789 21975 3847 21981
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 21981 6239 22015
rect 6362 22012 6368 22024
rect 6323 21984 6368 22012
rect 6181 21975 6239 21981
rect 2130 21953 2136 21956
rect 2124 21907 2136 21953
rect 2188 21944 2194 21956
rect 2188 21916 2224 21944
rect 2130 21904 2136 21907
rect 2188 21904 2194 21916
rect 3694 21904 3700 21956
rect 3752 21944 3758 21956
rect 4034 21947 4092 21953
rect 4034 21944 4046 21947
rect 3752 21916 4046 21944
rect 3752 21904 3758 21916
rect 4034 21913 4046 21916
rect 4080 21913 4092 21947
rect 4034 21907 4092 21913
rect 4154 21904 4160 21956
rect 4212 21944 4218 21956
rect 5074 21944 5080 21956
rect 4212 21916 5080 21944
rect 4212 21904 4218 21916
rect 5074 21904 5080 21916
rect 5132 21904 5138 21956
rect 6196 21944 6224 21975
rect 6362 21972 6368 21984
rect 6420 21972 6426 22024
rect 6472 22021 6500 22052
rect 6457 22015 6515 22021
rect 6457 21981 6469 22015
rect 6503 21981 6515 22015
rect 6457 21975 6515 21981
rect 6546 21972 6552 22024
rect 6604 22012 6610 22024
rect 6748 22012 6776 22052
rect 6825 22049 6837 22083
rect 6871 22080 6883 22083
rect 6914 22080 6920 22092
rect 6871 22052 6920 22080
rect 6871 22049 6883 22052
rect 6825 22043 6883 22049
rect 6914 22040 6920 22052
rect 6972 22040 6978 22092
rect 8956 22080 8984 22179
rect 14918 22176 14924 22188
rect 14976 22176 14982 22228
rect 15194 22176 15200 22228
rect 15252 22216 15258 22228
rect 16574 22216 16580 22228
rect 15252 22188 16580 22216
rect 15252 22176 15258 22188
rect 16574 22176 16580 22188
rect 16632 22216 16638 22228
rect 17678 22216 17684 22228
rect 16632 22188 17684 22216
rect 16632 22176 16638 22188
rect 17678 22176 17684 22188
rect 17736 22176 17742 22228
rect 18693 22219 18751 22225
rect 18693 22185 18705 22219
rect 18739 22216 18751 22219
rect 18782 22216 18788 22228
rect 18739 22188 18788 22216
rect 18739 22185 18751 22188
rect 18693 22179 18751 22185
rect 18782 22176 18788 22188
rect 18840 22176 18846 22228
rect 19429 22219 19487 22225
rect 19429 22185 19441 22219
rect 19475 22185 19487 22219
rect 19429 22179 19487 22185
rect 10318 22108 10324 22160
rect 10376 22148 10382 22160
rect 12802 22148 12808 22160
rect 10376 22120 12808 22148
rect 10376 22108 10382 22120
rect 12802 22108 12808 22120
rect 12860 22108 12866 22160
rect 16117 22151 16175 22157
rect 16117 22148 16129 22151
rect 15948 22120 16129 22148
rect 12345 22083 12403 22089
rect 7024 22052 7604 22080
rect 8956 22052 11560 22080
rect 7024 22024 7052 22052
rect 7006 22012 7012 22024
rect 6604 21984 6649 22012
rect 6748 21984 7012 22012
rect 6604 21972 6610 21984
rect 7006 21972 7012 21984
rect 7064 21972 7070 22024
rect 7282 22012 7288 22024
rect 7243 21984 7288 22012
rect 7282 21972 7288 21984
rect 7340 21972 7346 22024
rect 7466 22012 7472 22024
rect 7427 21984 7472 22012
rect 7466 21972 7472 21984
rect 7524 21972 7530 22024
rect 7576 22021 7604 22052
rect 7561 22015 7619 22021
rect 7561 21981 7573 22015
rect 7607 21981 7619 22015
rect 7561 21975 7619 21981
rect 7653 22015 7711 22021
rect 7653 21981 7665 22015
rect 7699 21981 7711 22015
rect 7653 21975 7711 21981
rect 6914 21944 6920 21956
rect 6196 21916 6920 21944
rect 6914 21904 6920 21916
rect 6972 21944 6978 21956
rect 7300 21944 7328 21972
rect 7668 21944 7696 21975
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 9861 22015 9919 22021
rect 9861 22012 9873 22015
rect 8444 21984 9873 22012
rect 8444 21972 8450 21984
rect 9861 21981 9873 21984
rect 9907 21981 9919 22015
rect 9861 21975 9919 21981
rect 9950 21972 9956 22024
rect 10008 22012 10014 22024
rect 10137 22015 10195 22021
rect 10137 22012 10149 22015
rect 10008 21984 10149 22012
rect 10008 21972 10014 21984
rect 10137 21981 10149 21984
rect 10183 21981 10195 22015
rect 10137 21975 10195 21981
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 22012 10287 22015
rect 11054 22012 11060 22024
rect 10275 21984 11060 22012
rect 10275 21981 10287 21984
rect 10229 21975 10287 21981
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 8294 21944 8300 21956
rect 6972 21916 7328 21944
rect 7576 21916 8300 21944
rect 6972 21904 6978 21916
rect 5166 21876 5172 21888
rect 5127 21848 5172 21876
rect 5166 21836 5172 21848
rect 5224 21836 5230 21888
rect 6730 21836 6736 21888
rect 6788 21876 6794 21888
rect 7576 21876 7604 21916
rect 8294 21904 8300 21916
rect 8352 21904 8358 21956
rect 10042 21944 10048 21956
rect 9955 21916 10048 21944
rect 10042 21904 10048 21916
rect 10100 21944 10106 21956
rect 11532 21944 11560 22052
rect 12345 22049 12357 22083
rect 12391 22080 12403 22083
rect 15838 22080 15844 22092
rect 12391 22052 15844 22080
rect 12391 22049 12403 22052
rect 12345 22043 12403 22049
rect 15838 22040 15844 22052
rect 15896 22040 15902 22092
rect 11609 22015 11667 22021
rect 11609 21981 11621 22015
rect 11655 22012 11667 22015
rect 12161 22015 12219 22021
rect 12161 22012 12173 22015
rect 11655 21984 12173 22012
rect 11655 21981 11667 21984
rect 11609 21975 11667 21981
rect 12161 21981 12173 21984
rect 12207 22012 12219 22015
rect 15194 22012 15200 22024
rect 12207 21984 15200 22012
rect 12207 21981 12219 21984
rect 12161 21975 12219 21981
rect 15194 21972 15200 21984
rect 15252 21972 15258 22024
rect 15948 21944 15976 22120
rect 16117 22117 16129 22120
rect 16163 22148 16175 22151
rect 16163 22120 16804 22148
rect 16163 22117 16175 22120
rect 16117 22111 16175 22117
rect 16776 22080 16804 22120
rect 17586 22108 17592 22160
rect 17644 22148 17650 22160
rect 19444 22148 19472 22179
rect 20806 22176 20812 22228
rect 20864 22216 20870 22228
rect 20990 22216 20996 22228
rect 20864 22188 20996 22216
rect 20864 22176 20870 22188
rect 20990 22176 20996 22188
rect 21048 22176 21054 22228
rect 22002 22176 22008 22228
rect 22060 22216 22066 22228
rect 22097 22219 22155 22225
rect 22097 22216 22109 22219
rect 22060 22188 22109 22216
rect 22060 22176 22066 22188
rect 22097 22185 22109 22188
rect 22143 22185 22155 22219
rect 22097 22179 22155 22185
rect 24302 22176 24308 22228
rect 24360 22216 24366 22228
rect 24397 22219 24455 22225
rect 24397 22216 24409 22219
rect 24360 22188 24409 22216
rect 24360 22176 24366 22188
rect 24397 22185 24409 22188
rect 24443 22185 24455 22219
rect 24397 22179 24455 22185
rect 28902 22176 28908 22228
rect 28960 22216 28966 22228
rect 28997 22219 29055 22225
rect 28997 22216 29009 22219
rect 28960 22188 29009 22216
rect 28960 22176 28966 22188
rect 28997 22185 29009 22188
rect 29043 22185 29055 22219
rect 28997 22179 29055 22185
rect 32493 22219 32551 22225
rect 32493 22185 32505 22219
rect 32539 22216 32551 22219
rect 33137 22219 33195 22225
rect 33137 22216 33149 22219
rect 32539 22188 33149 22216
rect 32539 22185 32551 22188
rect 32493 22179 32551 22185
rect 33137 22185 33149 22188
rect 33183 22185 33195 22219
rect 33137 22179 33195 22185
rect 22646 22148 22652 22160
rect 17644 22120 19472 22148
rect 20732 22120 22652 22148
rect 17644 22108 17650 22120
rect 17126 22080 17132 22092
rect 16132 22052 16528 22080
rect 16776 22052 17132 22080
rect 16132 22024 16160 22052
rect 16114 21972 16120 22024
rect 16172 21972 16178 22024
rect 16298 22012 16304 22024
rect 16259 21984 16304 22012
rect 16298 21972 16304 21984
rect 16356 21972 16362 22024
rect 16393 22015 16451 22021
rect 16393 21981 16405 22015
rect 16439 21981 16451 22015
rect 16393 21975 16451 21981
rect 16408 21944 16436 21975
rect 10100 21916 11468 21944
rect 11532 21916 15976 21944
rect 16316 21916 16436 21944
rect 16500 21944 16528 22052
rect 17126 22040 17132 22052
rect 17184 22040 17190 22092
rect 19334 22080 19340 22092
rect 18248 22052 19340 22080
rect 16942 21972 16948 22024
rect 17000 22012 17006 22024
rect 17218 22012 17224 22024
rect 17000 21984 17224 22012
rect 17000 21972 17006 21984
rect 17218 21972 17224 21984
rect 17276 21972 17282 22024
rect 17313 22015 17371 22021
rect 17313 21981 17325 22015
rect 17359 21981 17371 22015
rect 17313 21975 17371 21981
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 22012 17463 22015
rect 17494 22012 17500 22024
rect 17451 21984 17500 22012
rect 17451 21981 17463 21984
rect 17405 21975 17463 21981
rect 17328 21944 17356 21975
rect 17494 21972 17500 21984
rect 17552 21972 17558 22024
rect 17589 22015 17647 22021
rect 17589 21981 17601 22015
rect 17635 22012 17647 22015
rect 18046 22012 18052 22024
rect 17635 21984 18052 22012
rect 17635 21981 17647 21984
rect 17589 21975 17647 21981
rect 18046 21972 18052 21984
rect 18104 21972 18110 22024
rect 18248 22021 18276 22052
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 20732 22080 20760 22120
rect 22646 22108 22652 22120
rect 22704 22108 22710 22160
rect 19444 22052 20760 22080
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 18325 22015 18383 22021
rect 18325 21981 18337 22015
rect 18371 21981 18383 22015
rect 18325 21975 18383 21981
rect 18463 22015 18521 22021
rect 18463 21981 18475 22015
rect 18509 22012 18521 22015
rect 18598 22012 18604 22024
rect 18509 21984 18604 22012
rect 18509 21981 18521 21984
rect 18463 21975 18521 21981
rect 16500 21916 17954 21944
rect 10100 21904 10106 21916
rect 7926 21876 7932 21888
rect 6788 21848 7604 21876
rect 7887 21848 7932 21876
rect 6788 21836 6794 21848
rect 7926 21836 7932 21848
rect 7984 21836 7990 21888
rect 10413 21879 10471 21885
rect 10413 21845 10425 21879
rect 10459 21876 10471 21879
rect 10594 21876 10600 21888
rect 10459 21848 10600 21876
rect 10459 21845 10471 21848
rect 10413 21839 10471 21845
rect 10594 21836 10600 21848
rect 10652 21836 10658 21888
rect 11440 21876 11468 21916
rect 11698 21876 11704 21888
rect 11440 21848 11704 21876
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 15654 21876 15660 21888
rect 15615 21848 15660 21876
rect 15654 21836 15660 21848
rect 15712 21876 15718 21888
rect 16316 21876 16344 21916
rect 16942 21876 16948 21888
rect 15712 21848 16344 21876
rect 16903 21848 16948 21876
rect 15712 21836 15718 21848
rect 16942 21836 16948 21848
rect 17000 21836 17006 21888
rect 17926 21876 17954 21916
rect 18340 21876 18368 21975
rect 18598 21972 18604 21984
rect 18656 22012 18662 22024
rect 19444 22012 19472 22052
rect 20806 22040 20812 22092
rect 20864 22080 20870 22092
rect 22370 22080 22376 22092
rect 20864 22052 22376 22080
rect 20864 22040 20870 22052
rect 22370 22040 22376 22052
rect 22428 22040 22434 22092
rect 23566 22080 23572 22092
rect 23400 22052 23572 22080
rect 18656 21984 19472 22012
rect 19521 22015 19579 22021
rect 18656 21972 18662 21984
rect 19521 21981 19533 22015
rect 19567 21981 19579 22015
rect 19521 21975 19579 21981
rect 19613 22015 19671 22021
rect 19613 21981 19625 22015
rect 19659 22012 19671 22015
rect 21910 22012 21916 22024
rect 19659 21984 21916 22012
rect 19659 21981 19671 21984
rect 19613 21975 19671 21981
rect 19536 21944 19564 21975
rect 21910 21972 21916 21984
rect 21968 21972 21974 22024
rect 22554 21972 22560 22024
rect 22612 22012 22618 22024
rect 23400 22021 23428 22052
rect 23566 22040 23572 22052
rect 23624 22040 23630 22092
rect 25958 22040 25964 22092
rect 26016 22080 26022 22092
rect 29914 22080 29920 22092
rect 26016 22052 27752 22080
rect 26016 22040 26022 22052
rect 23293 22015 23351 22021
rect 23293 22012 23305 22015
rect 22612 21984 23305 22012
rect 22612 21972 22618 21984
rect 23293 21981 23305 21984
rect 23339 21981 23351 22015
rect 23293 21975 23351 21981
rect 23382 22015 23440 22021
rect 23382 21981 23394 22015
rect 23428 21981 23440 22015
rect 23382 21975 23440 21981
rect 23474 21972 23480 22024
rect 23532 22012 23538 22024
rect 23661 22015 23719 22021
rect 23532 21984 23577 22012
rect 23532 21972 23538 21984
rect 23661 21981 23673 22015
rect 23707 22012 23719 22015
rect 24302 22012 24308 22024
rect 23707 21984 24308 22012
rect 23707 21981 23719 21984
rect 23661 21975 23719 21981
rect 20714 21944 20720 21956
rect 19536 21916 20720 21944
rect 20714 21904 20720 21916
rect 20772 21904 20778 21956
rect 20809 21947 20867 21953
rect 20809 21913 20821 21947
rect 20855 21913 20867 21947
rect 20809 21907 20867 21913
rect 18414 21876 18420 21888
rect 17926 21848 18420 21876
rect 18414 21836 18420 21848
rect 18472 21836 18478 21888
rect 19058 21836 19064 21888
rect 19116 21876 19122 21888
rect 19245 21879 19303 21885
rect 19245 21876 19257 21879
rect 19116 21848 19257 21876
rect 19116 21836 19122 21848
rect 19245 21845 19257 21848
rect 19291 21845 19303 21879
rect 20254 21876 20260 21888
rect 20215 21848 20260 21876
rect 19245 21839 19303 21845
rect 20254 21836 20260 21848
rect 20312 21876 20318 21888
rect 20824 21876 20852 21907
rect 22094 21904 22100 21956
rect 22152 21944 22158 21956
rect 23676 21944 23704 21975
rect 24302 21972 24308 21984
rect 24360 21972 24366 22024
rect 26602 21972 26608 22024
rect 26660 22012 26666 22024
rect 27617 22015 27675 22021
rect 27617 22012 27629 22015
rect 26660 21984 27629 22012
rect 26660 21972 26666 21984
rect 27617 21981 27629 21984
rect 27663 21981 27675 22015
rect 27724 22012 27752 22052
rect 28644 22052 29920 22080
rect 28644 22012 28672 22052
rect 29914 22040 29920 22052
rect 29972 22040 29978 22092
rect 31386 22040 31392 22092
rect 31444 22080 31450 22092
rect 33318 22080 33324 22092
rect 31444 22052 32352 22080
rect 31444 22040 31450 22052
rect 27724 21984 28672 22012
rect 27617 21975 27675 21981
rect 29270 21972 29276 22024
rect 29328 22012 29334 22024
rect 31941 22015 31999 22021
rect 31941 22012 31953 22015
rect 29328 21984 31953 22012
rect 29328 21972 29334 21984
rect 31941 21981 31953 21984
rect 31987 21981 31999 22015
rect 31941 21975 31999 21981
rect 32030 21972 32036 22024
rect 32088 22012 32094 22024
rect 32324 22021 32352 22052
rect 33152 22052 33324 22080
rect 32217 22015 32275 22021
rect 32217 22012 32229 22015
rect 32088 21984 32229 22012
rect 32088 21972 32094 21984
rect 32217 21981 32229 21984
rect 32263 21981 32275 22015
rect 32217 21975 32275 21981
rect 32309 22015 32367 22021
rect 32309 21981 32321 22015
rect 32355 22012 32367 22015
rect 33042 22012 33048 22024
rect 32355 21984 33048 22012
rect 32355 21981 32367 21984
rect 32309 21975 32367 21981
rect 33042 21972 33048 21984
rect 33100 21972 33106 22024
rect 33152 22021 33180 22052
rect 33318 22040 33324 22052
rect 33376 22040 33382 22092
rect 33137 22015 33195 22021
rect 33137 21981 33149 22015
rect 33183 21981 33195 22015
rect 33137 21975 33195 21981
rect 33229 22015 33287 22021
rect 33229 21981 33241 22015
rect 33275 21981 33287 22015
rect 33410 22012 33416 22024
rect 33371 21984 33416 22012
rect 33229 21975 33287 21981
rect 22152 21916 23704 21944
rect 25332 21916 27016 21944
rect 22152 21904 22158 21916
rect 23014 21876 23020 21888
rect 20312 21848 20852 21876
rect 22975 21848 23020 21876
rect 20312 21836 20318 21848
rect 23014 21836 23020 21848
rect 23072 21836 23078 21888
rect 23658 21836 23664 21888
rect 23716 21876 23722 21888
rect 25332 21876 25360 21916
rect 26878 21876 26884 21888
rect 23716 21848 25360 21876
rect 26839 21848 26884 21876
rect 23716 21836 23722 21848
rect 26878 21836 26884 21848
rect 26936 21836 26942 21888
rect 26988 21876 27016 21916
rect 27706 21904 27712 21956
rect 27764 21944 27770 21956
rect 27862 21947 27920 21953
rect 27862 21944 27874 21947
rect 27764 21916 27874 21944
rect 27764 21904 27770 21916
rect 27862 21913 27874 21916
rect 27908 21913 27920 21947
rect 32122 21944 32128 21956
rect 32083 21916 32128 21944
rect 27862 21907 27920 21913
rect 32122 21904 32128 21916
rect 32180 21904 32186 21956
rect 33244 21944 33272 21975
rect 33410 21972 33416 21984
rect 33468 21972 33474 22024
rect 35986 22012 35992 22024
rect 35947 21984 35992 22012
rect 35986 21972 35992 21984
rect 36044 21972 36050 22024
rect 36078 21972 36084 22024
rect 36136 22012 36142 22024
rect 36357 22015 36415 22021
rect 36136 21984 36181 22012
rect 36136 21972 36142 21984
rect 36357 21981 36369 22015
rect 36403 22012 36415 22015
rect 37182 22012 37188 22024
rect 36403 21984 37188 22012
rect 36403 21981 36415 21984
rect 36357 21975 36415 21981
rect 37182 21972 37188 21984
rect 37240 21972 37246 22024
rect 39301 22015 39359 22021
rect 39301 21981 39313 22015
rect 39347 22012 39359 22015
rect 40034 22012 40040 22024
rect 39347 21984 40040 22012
rect 39347 21981 39359 21984
rect 39301 21975 39359 21981
rect 40034 21972 40040 21984
rect 40092 22012 40098 22024
rect 40129 22015 40187 22021
rect 40129 22012 40141 22015
rect 40092 21984 40141 22012
rect 40092 21972 40098 21984
rect 40129 21981 40141 21984
rect 40175 21981 40187 22015
rect 40129 21975 40187 21981
rect 40218 22012 40276 22018
rect 40218 21978 40230 22012
rect 40264 21978 40276 22012
rect 40218 21972 40276 21978
rect 33686 21944 33692 21956
rect 33244 21916 33692 21944
rect 33686 21904 33692 21916
rect 33744 21904 33750 21956
rect 36173 21947 36231 21953
rect 36173 21913 36185 21947
rect 36219 21944 36231 21947
rect 36262 21944 36268 21956
rect 36219 21916 36268 21944
rect 36219 21913 36231 21916
rect 36173 21907 36231 21913
rect 36262 21904 36268 21916
rect 36320 21904 36326 21956
rect 40233 21888 40261 21972
rect 40310 21969 40316 22021
rect 40368 22009 40374 22021
rect 40494 22012 40500 22024
rect 40368 21981 40410 22009
rect 40455 21984 40500 22012
rect 40368 21969 40374 21981
rect 40494 21972 40500 21984
rect 40552 21972 40558 22024
rect 32953 21879 33011 21885
rect 32953 21876 32965 21879
rect 26988 21848 32965 21876
rect 32953 21845 32965 21848
rect 32999 21845 33011 21879
rect 32953 21839 33011 21845
rect 35526 21836 35532 21888
rect 35584 21876 35590 21888
rect 35805 21879 35863 21885
rect 35805 21876 35817 21879
rect 35584 21848 35817 21876
rect 35584 21836 35590 21848
rect 35805 21845 35817 21848
rect 35851 21845 35863 21879
rect 39850 21876 39856 21888
rect 39811 21848 39856 21876
rect 35805 21839 35863 21845
rect 39850 21836 39856 21848
rect 39908 21836 39914 21888
rect 40218 21876 40224 21888
rect 40131 21848 40224 21876
rect 40218 21836 40224 21848
rect 40276 21876 40282 21888
rect 40954 21876 40960 21888
rect 40276 21848 40960 21876
rect 40276 21836 40282 21848
rect 40954 21836 40960 21848
rect 41012 21836 41018 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 2041 21675 2099 21681
rect 2041 21641 2053 21675
rect 2087 21672 2099 21675
rect 2130 21672 2136 21684
rect 2087 21644 2136 21672
rect 2087 21641 2099 21644
rect 2041 21635 2099 21641
rect 2130 21632 2136 21644
rect 2188 21632 2194 21684
rect 3694 21672 3700 21684
rect 3655 21644 3700 21672
rect 3694 21632 3700 21644
rect 3752 21632 3758 21684
rect 6086 21672 6092 21684
rect 4080 21644 6092 21672
rect 2774 21604 2780 21616
rect 2424 21576 2780 21604
rect 2424 21545 2452 21576
rect 2774 21564 2780 21576
rect 2832 21604 2838 21616
rect 4080 21604 4108 21644
rect 6086 21632 6092 21644
rect 6144 21632 6150 21684
rect 6178 21632 6184 21684
rect 6236 21672 6242 21684
rect 6365 21675 6423 21681
rect 6365 21672 6377 21675
rect 6236 21644 6377 21672
rect 6236 21632 6242 21644
rect 6365 21641 6377 21644
rect 6411 21672 6423 21675
rect 14642 21672 14648 21684
rect 6411 21644 14648 21672
rect 6411 21641 6423 21644
rect 6365 21635 6423 21641
rect 14642 21632 14648 21644
rect 14700 21632 14706 21684
rect 15930 21632 15936 21684
rect 15988 21672 15994 21684
rect 16298 21672 16304 21684
rect 15988 21644 16304 21672
rect 15988 21632 15994 21644
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 18046 21632 18052 21684
rect 18104 21672 18110 21684
rect 18104 21644 20668 21672
rect 18104 21632 18110 21644
rect 4614 21604 4620 21616
rect 2832 21576 4108 21604
rect 2832 21564 2838 21576
rect 2317 21539 2375 21545
rect 2317 21505 2329 21539
rect 2363 21505 2375 21539
rect 2317 21499 2375 21505
rect 2409 21539 2467 21545
rect 2409 21505 2421 21539
rect 2455 21505 2467 21539
rect 2409 21499 2467 21505
rect 2501 21539 2559 21545
rect 2501 21505 2513 21539
rect 2547 21536 2559 21539
rect 2590 21536 2596 21548
rect 2547 21508 2596 21536
rect 2547 21505 2559 21508
rect 2501 21499 2559 21505
rect 2332 21468 2360 21499
rect 2590 21496 2596 21508
rect 2648 21496 2654 21548
rect 2685 21539 2743 21545
rect 2685 21505 2697 21539
rect 2731 21505 2743 21539
rect 3970 21536 3976 21548
rect 3931 21508 3976 21536
rect 2685 21499 2743 21505
rect 2332 21440 2452 21468
rect 2424 21332 2452 21440
rect 2700 21400 2728 21499
rect 3970 21496 3976 21508
rect 4028 21496 4034 21548
rect 4080 21545 4108 21576
rect 4172 21576 4620 21604
rect 4172 21545 4200 21576
rect 4614 21564 4620 21576
rect 4672 21564 4678 21616
rect 4893 21607 4951 21613
rect 4893 21573 4905 21607
rect 4939 21604 4951 21607
rect 5074 21604 5080 21616
rect 4939 21576 5080 21604
rect 4939 21573 4951 21576
rect 4893 21567 4951 21573
rect 5074 21564 5080 21576
rect 5132 21564 5138 21616
rect 5166 21564 5172 21616
rect 5224 21604 5230 21616
rect 7500 21607 7558 21613
rect 5224 21576 7374 21604
rect 5224 21564 5230 21576
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 4157 21539 4215 21545
rect 4157 21505 4169 21539
rect 4203 21505 4215 21539
rect 4341 21539 4399 21545
rect 4341 21536 4353 21539
rect 4157 21499 4215 21505
rect 4264 21508 4353 21536
rect 4264 21400 4292 21508
rect 4341 21505 4353 21508
rect 4387 21536 4399 21539
rect 6914 21536 6920 21548
rect 4387 21508 6920 21536
rect 4387 21505 4399 21508
rect 4341 21499 4399 21505
rect 6914 21496 6920 21508
rect 6972 21496 6978 21548
rect 7346 21536 7374 21576
rect 7500 21573 7512 21607
rect 7546 21604 7558 21607
rect 7926 21604 7932 21616
rect 7546 21576 7932 21604
rect 7546 21573 7558 21576
rect 7500 21567 7558 21573
rect 7926 21564 7932 21576
rect 7984 21564 7990 21616
rect 8294 21604 8300 21616
rect 8255 21576 8300 21604
rect 8294 21564 8300 21576
rect 8352 21564 8358 21616
rect 10134 21604 10140 21616
rect 10095 21576 10140 21604
rect 10134 21564 10140 21576
rect 10192 21564 10198 21616
rect 15749 21607 15807 21613
rect 15749 21573 15761 21607
rect 15795 21604 15807 21607
rect 16390 21604 16396 21616
rect 15795 21576 16396 21604
rect 15795 21573 15807 21576
rect 15749 21567 15807 21573
rect 16390 21564 16396 21576
rect 16448 21564 16454 21616
rect 16942 21613 16948 21616
rect 16936 21604 16948 21613
rect 16903 21576 16948 21604
rect 16936 21567 16948 21576
rect 16942 21564 16948 21567
rect 17000 21564 17006 21616
rect 20640 21604 20668 21644
rect 20714 21632 20720 21684
rect 20772 21672 20778 21684
rect 25958 21672 25964 21684
rect 20772 21644 25964 21672
rect 20772 21632 20778 21644
rect 25958 21632 25964 21644
rect 26016 21632 26022 21684
rect 27617 21675 27675 21681
rect 27617 21641 27629 21675
rect 27663 21672 27675 21675
rect 27706 21672 27712 21684
rect 27663 21644 27712 21672
rect 27663 21641 27675 21644
rect 27617 21635 27675 21641
rect 27706 21632 27712 21644
rect 27764 21632 27770 21684
rect 28810 21632 28816 21684
rect 28868 21672 28874 21684
rect 29549 21675 29607 21681
rect 29549 21672 29561 21675
rect 28868 21644 29561 21672
rect 28868 21632 28874 21644
rect 29549 21641 29561 21644
rect 29595 21641 29607 21675
rect 29549 21635 29607 21641
rect 29638 21632 29644 21684
rect 29696 21672 29702 21684
rect 32030 21672 32036 21684
rect 29696 21644 32036 21672
rect 29696 21632 29702 21644
rect 32030 21632 32036 21644
rect 32088 21632 32094 21684
rect 32769 21675 32827 21681
rect 32769 21641 32781 21675
rect 32815 21641 32827 21675
rect 34606 21672 34612 21684
rect 32769 21635 32827 21641
rect 32876 21644 34612 21672
rect 20993 21607 21051 21613
rect 20993 21604 21005 21607
rect 20640 21576 21005 21604
rect 20993 21573 21005 21576
rect 21039 21604 21051 21607
rect 21818 21604 21824 21616
rect 21039 21576 21824 21604
rect 21039 21573 21051 21576
rect 20993 21567 21051 21573
rect 21818 21564 21824 21576
rect 21876 21564 21882 21616
rect 23014 21564 23020 21616
rect 23072 21604 23078 21616
rect 23302 21607 23360 21613
rect 23302 21604 23314 21607
rect 23072 21576 23314 21604
rect 23072 21564 23078 21576
rect 23302 21573 23314 21576
rect 23348 21573 23360 21607
rect 23302 21567 23360 21573
rect 23934 21564 23940 21616
rect 23992 21604 23998 21616
rect 32784 21604 32812 21635
rect 23992 21576 29040 21604
rect 23992 21564 23998 21576
rect 9861 21539 9919 21545
rect 9861 21536 9873 21539
rect 7346 21508 9873 21536
rect 9861 21505 9873 21508
rect 9907 21505 9919 21539
rect 10042 21536 10048 21548
rect 10003 21508 10048 21536
rect 9861 21499 9919 21505
rect 10042 21496 10048 21508
rect 10100 21496 10106 21548
rect 10229 21539 10287 21545
rect 10229 21505 10241 21539
rect 10275 21536 10287 21539
rect 11054 21536 11060 21548
rect 10275 21508 11060 21536
rect 10275 21505 10287 21508
rect 10229 21499 10287 21505
rect 11054 21496 11060 21508
rect 11112 21496 11118 21548
rect 15378 21536 15384 21548
rect 15339 21508 15384 21536
rect 15378 21496 15384 21508
rect 15436 21496 15442 21548
rect 15474 21539 15532 21545
rect 15474 21505 15486 21539
rect 15520 21505 15532 21539
rect 15474 21499 15532 21505
rect 15657 21539 15715 21545
rect 15657 21505 15669 21539
rect 15703 21505 15715 21539
rect 15657 21499 15715 21505
rect 15887 21539 15945 21545
rect 15887 21505 15899 21539
rect 15933 21536 15945 21539
rect 16298 21536 16304 21548
rect 15933 21508 16304 21536
rect 15933 21505 15945 21508
rect 15887 21499 15945 21505
rect 7745 21471 7803 21477
rect 7745 21437 7757 21471
rect 7791 21468 7803 21471
rect 8294 21468 8300 21480
rect 7791 21440 8300 21468
rect 7791 21437 7803 21440
rect 7745 21431 7803 21437
rect 8294 21428 8300 21440
rect 8352 21428 8358 21480
rect 13998 21428 14004 21480
rect 14056 21468 14062 21480
rect 15488 21468 15516 21499
rect 14056 21440 15516 21468
rect 15672 21468 15700 21499
rect 16298 21496 16304 21508
rect 16356 21496 16362 21548
rect 16482 21496 16488 21548
rect 16540 21536 16546 21548
rect 16669 21539 16727 21545
rect 16669 21536 16681 21539
rect 16540 21508 16681 21536
rect 16540 21496 16546 21508
rect 16669 21505 16681 21508
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 17218 21496 17224 21548
rect 17276 21536 17282 21548
rect 17276 21508 17724 21536
rect 17276 21496 17282 21508
rect 17696 21468 17724 21508
rect 20438 21496 20444 21548
rect 20496 21536 20502 21548
rect 21177 21539 21235 21545
rect 21177 21536 21189 21539
rect 20496 21508 21189 21536
rect 20496 21496 20502 21508
rect 21177 21505 21189 21508
rect 21223 21505 21235 21539
rect 21177 21499 21235 21505
rect 21542 21496 21548 21548
rect 21600 21536 21606 21548
rect 26694 21536 26700 21548
rect 21600 21508 26700 21536
rect 21600 21496 21606 21508
rect 26694 21496 26700 21508
rect 26752 21496 26758 21548
rect 27893 21539 27951 21545
rect 27893 21536 27905 21539
rect 27264 21508 27905 21536
rect 23569 21471 23627 21477
rect 15672 21440 16160 21468
rect 17696 21440 21128 21468
rect 14056 21428 14062 21440
rect 2700 21372 4292 21400
rect 8110 21360 8116 21412
rect 8168 21400 8174 21412
rect 12434 21400 12440 21412
rect 8168 21372 12440 21400
rect 8168 21360 8174 21372
rect 12434 21360 12440 21372
rect 12492 21360 12498 21412
rect 13630 21360 13636 21412
rect 13688 21400 13694 21412
rect 16025 21403 16083 21409
rect 16025 21400 16037 21403
rect 13688 21372 16037 21400
rect 13688 21360 13694 21372
rect 16025 21369 16037 21372
rect 16071 21369 16083 21403
rect 16025 21363 16083 21369
rect 2498 21332 2504 21344
rect 2411 21304 2504 21332
rect 2498 21292 2504 21304
rect 2556 21332 2562 21344
rect 3234 21332 3240 21344
rect 2556 21304 3240 21332
rect 2556 21292 2562 21304
rect 3234 21292 3240 21304
rect 3292 21292 3298 21344
rect 10413 21335 10471 21341
rect 10413 21301 10425 21335
rect 10459 21332 10471 21335
rect 11422 21332 11428 21344
rect 10459 21304 11428 21332
rect 10459 21301 10471 21304
rect 10413 21295 10471 21301
rect 11422 21292 11428 21304
rect 11480 21292 11486 21344
rect 14274 21332 14280 21344
rect 14235 21304 14280 21332
rect 14274 21292 14280 21304
rect 14332 21292 14338 21344
rect 16132 21332 16160 21440
rect 20438 21400 20444 21412
rect 17604 21372 20444 21400
rect 17604 21344 17632 21372
rect 20438 21360 20444 21372
rect 20496 21360 20502 21412
rect 21100 21400 21128 21440
rect 23569 21437 23581 21471
rect 23615 21468 23627 21471
rect 26602 21468 26608 21480
rect 23615 21440 26608 21468
rect 23615 21437 23627 21440
rect 23569 21431 23627 21437
rect 22554 21400 22560 21412
rect 21100 21372 22560 21400
rect 22554 21360 22560 21372
rect 22612 21360 22618 21412
rect 16942 21332 16948 21344
rect 16132 21304 16948 21332
rect 16942 21292 16948 21304
rect 17000 21292 17006 21344
rect 17586 21292 17592 21344
rect 17644 21292 17650 21344
rect 18046 21332 18052 21344
rect 18007 21304 18052 21332
rect 18046 21292 18052 21304
rect 18104 21292 18110 21344
rect 22186 21332 22192 21344
rect 22147 21304 22192 21332
rect 22186 21292 22192 21304
rect 22244 21292 22250 21344
rect 23198 21292 23204 21344
rect 23256 21332 23262 21344
rect 23584 21332 23612 21431
rect 26602 21428 26608 21440
rect 26660 21428 26666 21480
rect 27264 21344 27292 21508
rect 27893 21505 27905 21508
rect 27939 21505 27951 21539
rect 27893 21499 27951 21505
rect 27985 21539 28043 21545
rect 27985 21505 27997 21539
rect 28031 21505 28043 21539
rect 27985 21499 28043 21505
rect 27430 21428 27436 21480
rect 27488 21468 27494 21480
rect 28000 21468 28028 21499
rect 28074 21496 28080 21548
rect 28132 21536 28138 21548
rect 28258 21536 28264 21548
rect 28132 21508 28177 21536
rect 28219 21508 28264 21536
rect 28132 21496 28138 21508
rect 28258 21496 28264 21508
rect 28316 21496 28322 21548
rect 28442 21496 28448 21548
rect 28500 21536 28506 21548
rect 28905 21539 28963 21545
rect 28905 21536 28917 21539
rect 28500 21508 28917 21536
rect 28500 21496 28506 21508
rect 28905 21505 28917 21508
rect 28951 21505 28963 21539
rect 29012 21536 29040 21576
rect 29656 21576 32812 21604
rect 29656 21536 29684 21576
rect 29012 21508 29684 21536
rect 29733 21539 29791 21545
rect 28905 21499 28963 21505
rect 29733 21505 29745 21539
rect 29779 21505 29791 21539
rect 29733 21499 29791 21505
rect 30009 21539 30067 21545
rect 30009 21505 30021 21539
rect 30055 21536 30067 21539
rect 32876 21536 32904 21644
rect 34606 21632 34612 21644
rect 34664 21632 34670 21684
rect 33229 21607 33287 21613
rect 33229 21573 33241 21607
rect 33275 21604 33287 21607
rect 33594 21604 33600 21616
rect 33275 21576 33600 21604
rect 33275 21573 33287 21576
rect 33229 21567 33287 21573
rect 33594 21564 33600 21576
rect 33652 21564 33658 21616
rect 39700 21607 39758 21613
rect 39700 21573 39712 21607
rect 39746 21604 39758 21607
rect 39850 21604 39856 21616
rect 39746 21576 39856 21604
rect 39746 21573 39758 21576
rect 39700 21567 39758 21573
rect 39850 21564 39856 21576
rect 39908 21564 39914 21616
rect 30055 21508 32904 21536
rect 32953 21539 33011 21545
rect 30055 21505 30067 21508
rect 30009 21499 30067 21505
rect 32953 21505 32965 21539
rect 32999 21536 33011 21539
rect 33134 21536 33140 21548
rect 32999 21508 33140 21536
rect 32999 21505 33011 21508
rect 32953 21499 33011 21505
rect 28994 21468 29000 21480
rect 27488 21440 29000 21468
rect 27488 21428 27494 21440
rect 28994 21428 29000 21440
rect 29052 21428 29058 21480
rect 29089 21471 29147 21477
rect 29089 21437 29101 21471
rect 29135 21468 29147 21471
rect 29638 21468 29644 21480
rect 29135 21440 29644 21468
rect 29135 21437 29147 21440
rect 29089 21431 29147 21437
rect 29638 21428 29644 21440
rect 29696 21428 29702 21480
rect 29748 21400 29776 21499
rect 33134 21496 33140 21508
rect 33192 21496 33198 21548
rect 29822 21428 29828 21480
rect 29880 21468 29886 21480
rect 29880 21440 29925 21468
rect 29880 21428 29886 21440
rect 31846 21428 31852 21480
rect 31904 21468 31910 21480
rect 33045 21471 33103 21477
rect 33045 21468 33057 21471
rect 31904 21440 33057 21468
rect 31904 21428 31910 21440
rect 33045 21437 33057 21440
rect 33091 21437 33103 21471
rect 39942 21468 39948 21480
rect 39903 21440 39948 21468
rect 33045 21431 33103 21437
rect 39942 21428 39948 21440
rect 40000 21428 40006 21480
rect 37274 21400 37280 21412
rect 29748 21372 37280 21400
rect 37274 21360 37280 21372
rect 37332 21360 37338 21412
rect 23256 21304 23612 21332
rect 27157 21335 27215 21341
rect 23256 21292 23262 21304
rect 27157 21301 27169 21335
rect 27203 21332 27215 21335
rect 27246 21332 27252 21344
rect 27203 21304 27252 21332
rect 27203 21301 27215 21304
rect 27157 21295 27215 21301
rect 27246 21292 27252 21304
rect 27304 21292 27310 21344
rect 29730 21332 29736 21344
rect 29691 21304 29736 21332
rect 29730 21292 29736 21304
rect 29788 21292 29794 21344
rect 32950 21332 32956 21344
rect 32911 21304 32956 21332
rect 32950 21292 32956 21304
rect 33008 21292 33014 21344
rect 35894 21332 35900 21344
rect 35855 21304 35900 21332
rect 35894 21292 35900 21304
rect 35952 21332 35958 21344
rect 36354 21332 36360 21344
rect 35952 21304 36360 21332
rect 35952 21292 35958 21304
rect 36354 21292 36360 21304
rect 36412 21292 36418 21344
rect 37826 21292 37832 21344
rect 37884 21332 37890 21344
rect 38562 21332 38568 21344
rect 37884 21304 38568 21332
rect 37884 21292 37890 21304
rect 38562 21292 38568 21304
rect 38620 21292 38626 21344
rect 58158 21332 58164 21344
rect 58119 21304 58164 21332
rect 58158 21292 58164 21304
rect 58216 21292 58222 21344
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 6365 21131 6423 21137
rect 6365 21097 6377 21131
rect 6411 21128 6423 21131
rect 7466 21128 7472 21140
rect 6411 21100 7472 21128
rect 6411 21097 6423 21100
rect 6365 21091 6423 21097
rect 7466 21088 7472 21100
rect 7524 21088 7530 21140
rect 10597 21131 10655 21137
rect 10597 21097 10609 21131
rect 10643 21128 10655 21131
rect 10686 21128 10692 21140
rect 10643 21100 10692 21128
rect 10643 21097 10655 21100
rect 10597 21091 10655 21097
rect 10686 21088 10692 21100
rect 10744 21088 10750 21140
rect 15841 21131 15899 21137
rect 15841 21097 15853 21131
rect 15887 21128 15899 21131
rect 16482 21128 16488 21140
rect 15887 21100 16488 21128
rect 15887 21097 15899 21100
rect 15841 21091 15899 21097
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 17494 21088 17500 21140
rect 17552 21128 17558 21140
rect 17589 21131 17647 21137
rect 17589 21128 17601 21131
rect 17552 21100 17601 21128
rect 17552 21088 17558 21100
rect 17589 21097 17601 21100
rect 17635 21097 17647 21131
rect 17589 21091 17647 21097
rect 22281 21131 22339 21137
rect 22281 21097 22293 21131
rect 22327 21128 22339 21131
rect 23474 21128 23480 21140
rect 22327 21100 23480 21128
rect 22327 21097 22339 21100
rect 22281 21091 22339 21097
rect 23474 21088 23480 21100
rect 23532 21088 23538 21140
rect 26326 21088 26332 21140
rect 26384 21128 26390 21140
rect 26694 21128 26700 21140
rect 26384 21100 26700 21128
rect 26384 21088 26390 21100
rect 26694 21088 26700 21100
rect 26752 21088 26758 21140
rect 32030 21088 32036 21140
rect 32088 21128 32094 21140
rect 35894 21128 35900 21140
rect 32088 21100 35900 21128
rect 32088 21088 32094 21100
rect 35894 21088 35900 21100
rect 35952 21088 35958 21140
rect 6638 21020 6644 21072
rect 6696 21060 6702 21072
rect 6917 21063 6975 21069
rect 6917 21060 6929 21063
rect 6696 21032 6929 21060
rect 6696 21020 6702 21032
rect 6917 21029 6929 21032
rect 6963 21029 6975 21063
rect 8110 21060 8116 21072
rect 8071 21032 8116 21060
rect 6917 21023 6975 21029
rect 8110 21020 8116 21032
rect 8168 21020 8174 21072
rect 11606 21060 11612 21072
rect 11567 21032 11612 21060
rect 11606 21020 11612 21032
rect 11664 21020 11670 21072
rect 12437 21063 12495 21069
rect 12437 21029 12449 21063
rect 12483 21060 12495 21063
rect 13906 21060 13912 21072
rect 12483 21032 13912 21060
rect 12483 21029 12495 21032
rect 12437 21023 12495 21029
rect 12452 20992 12480 21023
rect 13906 21020 13912 21032
rect 13964 21020 13970 21072
rect 16298 21020 16304 21072
rect 16356 21060 16362 21072
rect 20257 21063 20315 21069
rect 20257 21060 20269 21063
rect 16356 21032 20269 21060
rect 16356 21020 16362 21032
rect 20257 21029 20269 21032
rect 20303 21060 20315 21063
rect 21450 21060 21456 21072
rect 20303 21032 21456 21060
rect 20303 21029 20315 21032
rect 20257 21023 20315 21029
rect 21450 21020 21456 21032
rect 21508 21020 21514 21072
rect 24762 21060 24768 21072
rect 21928 21032 24768 21060
rect 11808 20964 12480 20992
rect 5994 20924 6000 20936
rect 5955 20896 6000 20924
rect 5994 20884 6000 20896
rect 6052 20884 6058 20936
rect 6178 20924 6184 20936
rect 6139 20896 6184 20924
rect 6178 20884 6184 20896
rect 6236 20884 6242 20936
rect 11808 20933 11836 20964
rect 13446 20952 13452 21004
rect 13504 20992 13510 21004
rect 14737 20995 14795 21001
rect 14737 20992 14749 20995
rect 13504 20964 14749 20992
rect 13504 20952 13510 20964
rect 14737 20961 14749 20964
rect 14783 20992 14795 20995
rect 18138 20992 18144 21004
rect 14783 20964 18144 20992
rect 14783 20961 14795 20964
rect 14737 20955 14795 20961
rect 18138 20952 18144 20964
rect 18196 20952 18202 21004
rect 11793 20927 11851 20933
rect 11793 20893 11805 20927
rect 11839 20893 11851 20927
rect 11793 20887 11851 20893
rect 12989 20927 13047 20933
rect 12989 20893 13001 20927
rect 13035 20924 13047 20927
rect 13354 20924 13360 20936
rect 13035 20896 13360 20924
rect 13035 20893 13047 20896
rect 12989 20887 13047 20893
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 13906 20884 13912 20936
rect 13964 20924 13970 20936
rect 14274 20924 14280 20936
rect 13964 20896 14280 20924
rect 13964 20884 13970 20896
rect 14274 20884 14280 20896
rect 14332 20924 14338 20936
rect 14553 20927 14611 20933
rect 14553 20924 14565 20927
rect 14332 20896 14565 20924
rect 14332 20884 14338 20896
rect 14553 20893 14565 20896
rect 14599 20924 14611 20927
rect 17586 20924 17592 20936
rect 14599 20896 17592 20924
rect 14599 20893 14611 20896
rect 14553 20887 14611 20893
rect 17586 20884 17592 20896
rect 17644 20884 17650 20936
rect 17773 20927 17831 20933
rect 17773 20893 17785 20927
rect 17819 20924 17831 20927
rect 18046 20924 18052 20936
rect 17819 20896 18052 20924
rect 17819 20893 17831 20896
rect 17773 20887 17831 20893
rect 18046 20884 18052 20896
rect 18104 20924 18110 20936
rect 19334 20924 19340 20936
rect 18104 20896 19340 20924
rect 18104 20884 18110 20896
rect 19334 20884 19340 20896
rect 19392 20884 19398 20936
rect 8297 20859 8355 20865
rect 8297 20825 8309 20859
rect 8343 20856 8355 20859
rect 8386 20856 8392 20868
rect 8343 20828 8392 20856
rect 8343 20825 8355 20828
rect 8297 20819 8355 20825
rect 8386 20816 8392 20828
rect 8444 20816 8450 20868
rect 9861 20859 9919 20865
rect 9861 20825 9873 20859
rect 9907 20856 9919 20859
rect 10689 20859 10747 20865
rect 10689 20856 10701 20859
rect 9907 20828 10701 20856
rect 9907 20825 9919 20828
rect 9861 20819 9919 20825
rect 10689 20825 10701 20828
rect 10735 20856 10747 20859
rect 10962 20856 10968 20868
rect 10735 20828 10968 20856
rect 10735 20825 10747 20828
rect 10689 20819 10747 20825
rect 10962 20816 10968 20828
rect 11020 20816 11026 20868
rect 13173 20859 13231 20865
rect 13173 20825 13185 20859
rect 13219 20856 13231 20859
rect 13998 20856 14004 20868
rect 13219 20828 14004 20856
rect 13219 20825 13231 20828
rect 13173 20819 13231 20825
rect 13998 20816 14004 20828
rect 14056 20816 14062 20868
rect 16022 20816 16028 20868
rect 16080 20856 16086 20868
rect 17129 20859 17187 20865
rect 17129 20856 17141 20859
rect 16080 20828 17141 20856
rect 16080 20816 16086 20828
rect 17129 20825 17141 20828
rect 17175 20825 17187 20859
rect 17954 20856 17960 20868
rect 17915 20828 17960 20856
rect 17129 20819 17187 20825
rect 17954 20816 17960 20828
rect 18012 20816 18018 20868
rect 20162 20816 20168 20868
rect 20220 20856 20226 20868
rect 20441 20859 20499 20865
rect 20441 20856 20453 20859
rect 20220 20828 20453 20856
rect 20220 20816 20226 20828
rect 20441 20825 20453 20828
rect 20487 20825 20499 20859
rect 20441 20819 20499 20825
rect 21266 20816 21272 20868
rect 21324 20856 21330 20868
rect 21928 20865 21956 21032
rect 24762 21020 24768 21032
rect 24820 21020 24826 21072
rect 22094 20952 22100 21004
rect 22152 20952 22158 21004
rect 23032 20964 23345 20992
rect 22112 20924 22140 20952
rect 22747 20927 22805 20933
rect 23032 20930 23060 20964
rect 22747 20924 22759 20927
rect 22112 20896 22759 20924
rect 22747 20893 22759 20896
rect 22793 20893 22805 20927
rect 22904 20921 22962 20927
rect 22904 20918 22916 20921
rect 22747 20887 22805 20893
rect 22848 20890 22916 20918
rect 21913 20859 21971 20865
rect 21913 20856 21925 20859
rect 21324 20828 21925 20856
rect 21324 20816 21330 20828
rect 21913 20825 21925 20828
rect 21959 20825 21971 20859
rect 21913 20819 21971 20825
rect 22097 20859 22155 20865
rect 22097 20825 22109 20859
rect 22143 20856 22155 20859
rect 22186 20856 22192 20868
rect 22143 20828 22192 20856
rect 22143 20825 22155 20828
rect 22097 20819 22155 20825
rect 22186 20816 22192 20828
rect 22244 20816 22250 20868
rect 22848 20800 22876 20890
rect 22904 20887 22916 20890
rect 22950 20887 22962 20921
rect 22904 20881 22962 20887
rect 23004 20924 23062 20930
rect 23004 20890 23016 20924
rect 23050 20890 23062 20924
rect 23004 20884 23062 20890
rect 23106 20884 23112 20936
rect 23164 20924 23170 20936
rect 23164 20896 23209 20924
rect 23317 20921 23345 20964
rect 23566 20924 23572 20936
rect 23391 20921 23572 20924
rect 23317 20896 23572 20921
rect 23164 20884 23170 20896
rect 23317 20893 23419 20896
rect 23566 20884 23572 20896
rect 23624 20884 23630 20936
rect 24780 20933 24808 21020
rect 27154 20952 27160 21004
rect 27212 20992 27218 21004
rect 28997 20995 29055 21001
rect 28997 20992 29009 20995
rect 27212 20964 29009 20992
rect 27212 20952 27218 20964
rect 28997 20961 29009 20964
rect 29043 20992 29055 20995
rect 29178 20992 29184 21004
rect 29043 20964 29184 20992
rect 29043 20961 29055 20964
rect 28997 20955 29055 20961
rect 29178 20952 29184 20964
rect 29236 20952 29242 21004
rect 24765 20927 24823 20933
rect 24765 20893 24777 20927
rect 24811 20893 24823 20927
rect 26602 20924 26608 20936
rect 26563 20896 26608 20924
rect 24765 20887 24823 20893
rect 26602 20884 26608 20896
rect 26660 20884 26666 20936
rect 27246 20884 27252 20936
rect 27304 20924 27310 20936
rect 27341 20927 27399 20933
rect 27341 20924 27353 20927
rect 27304 20896 27353 20924
rect 27304 20884 27310 20896
rect 27341 20893 27353 20896
rect 27387 20924 27399 20927
rect 27387 20896 31754 20924
rect 27387 20893 27399 20896
rect 27341 20887 27399 20893
rect 23474 20816 23480 20868
rect 23532 20856 23538 20868
rect 24397 20859 24455 20865
rect 24397 20856 24409 20859
rect 23532 20828 24409 20856
rect 23532 20816 23538 20828
rect 24397 20825 24409 20828
rect 24443 20825 24455 20859
rect 24578 20856 24584 20868
rect 24539 20828 24584 20856
rect 24397 20819 24455 20825
rect 24578 20816 24584 20828
rect 24636 20816 24642 20868
rect 26360 20859 26418 20865
rect 26360 20825 26372 20859
rect 26406 20856 26418 20859
rect 26970 20856 26976 20868
rect 26406 20828 26976 20856
rect 26406 20825 26418 20828
rect 26360 20819 26418 20825
rect 26970 20816 26976 20828
rect 27028 20816 27034 20868
rect 27157 20859 27215 20865
rect 27157 20825 27169 20859
rect 27203 20825 27215 20859
rect 27157 20819 27215 20825
rect 13262 20748 13268 20800
rect 13320 20788 13326 20800
rect 13357 20791 13415 20797
rect 13357 20788 13369 20791
rect 13320 20760 13369 20788
rect 13320 20748 13326 20760
rect 13357 20757 13369 20760
rect 13403 20757 13415 20791
rect 13357 20751 13415 20757
rect 16942 20748 16948 20800
rect 17000 20788 17006 20800
rect 21726 20788 21732 20800
rect 17000 20760 21732 20788
rect 17000 20748 17006 20760
rect 21726 20748 21732 20760
rect 21784 20748 21790 20800
rect 22830 20748 22836 20800
rect 22888 20748 22894 20800
rect 23382 20788 23388 20800
rect 23343 20760 23388 20788
rect 23382 20748 23388 20760
rect 23440 20748 23446 20800
rect 25222 20788 25228 20800
rect 25183 20760 25228 20788
rect 25222 20748 25228 20760
rect 25280 20748 25286 20800
rect 26234 20748 26240 20800
rect 26292 20788 26298 20800
rect 26878 20788 26884 20800
rect 26292 20760 26884 20788
rect 26292 20748 26298 20760
rect 26878 20748 26884 20760
rect 26936 20788 26942 20800
rect 27172 20788 27200 20819
rect 29178 20816 29184 20868
rect 29236 20856 29242 20868
rect 30009 20859 30067 20865
rect 30009 20856 30021 20859
rect 29236 20828 30021 20856
rect 29236 20816 29242 20828
rect 30009 20825 30021 20828
rect 30055 20825 30067 20859
rect 31726 20856 31754 20896
rect 31726 20828 32260 20856
rect 30009 20819 30067 20825
rect 32232 20800 32260 20828
rect 26936 20760 27200 20788
rect 26936 20748 26942 20760
rect 27246 20748 27252 20800
rect 27304 20788 27310 20800
rect 27801 20791 27859 20797
rect 27801 20788 27813 20791
rect 27304 20760 27813 20788
rect 27304 20748 27310 20760
rect 27801 20757 27813 20760
rect 27847 20757 27859 20791
rect 28442 20788 28448 20800
rect 28403 20760 28448 20788
rect 27801 20751 27859 20757
rect 28442 20748 28448 20760
rect 28500 20748 28506 20800
rect 28994 20748 29000 20800
rect 29052 20788 29058 20800
rect 29822 20788 29828 20800
rect 29052 20760 29828 20788
rect 29052 20748 29058 20760
rect 29822 20748 29828 20760
rect 29880 20748 29886 20800
rect 30098 20788 30104 20800
rect 30059 20760 30104 20788
rect 30098 20748 30104 20760
rect 30156 20788 30162 20800
rect 30374 20788 30380 20800
rect 30156 20760 30380 20788
rect 30156 20748 30162 20760
rect 30374 20748 30380 20760
rect 30432 20748 30438 20800
rect 32214 20788 32220 20800
rect 32175 20760 32220 20788
rect 32214 20748 32220 20760
rect 32272 20748 32278 20800
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 7561 20587 7619 20593
rect 7561 20584 7573 20587
rect 6886 20556 7573 20584
rect 3050 20476 3056 20528
rect 3108 20516 3114 20528
rect 6886 20516 6914 20556
rect 7561 20553 7573 20556
rect 7607 20584 7619 20587
rect 11238 20584 11244 20596
rect 7607 20556 11244 20584
rect 7607 20553 7619 20556
rect 7561 20547 7619 20553
rect 11238 20544 11244 20556
rect 11296 20544 11302 20596
rect 11606 20544 11612 20596
rect 11664 20584 11670 20596
rect 11882 20584 11888 20596
rect 11664 20556 11888 20584
rect 11664 20544 11670 20556
rect 11882 20544 11888 20556
rect 11940 20584 11946 20596
rect 11977 20587 12035 20593
rect 11977 20584 11989 20587
rect 11940 20556 11989 20584
rect 11940 20544 11946 20556
rect 11977 20553 11989 20556
rect 12023 20553 12035 20587
rect 13998 20584 14004 20596
rect 13959 20556 14004 20584
rect 11977 20547 12035 20553
rect 13998 20544 14004 20556
rect 14056 20544 14062 20596
rect 16022 20584 16028 20596
rect 15983 20556 16028 20584
rect 16022 20544 16028 20556
rect 16080 20544 16086 20596
rect 16942 20584 16948 20596
rect 16903 20556 16948 20584
rect 16942 20544 16948 20556
rect 17000 20544 17006 20596
rect 17788 20556 22600 20584
rect 16482 20516 16488 20528
rect 3108 20488 6914 20516
rect 12636 20488 16488 20516
rect 3108 20476 3114 20488
rect 4798 20448 4804 20460
rect 4711 20420 4804 20448
rect 4798 20408 4804 20420
rect 4856 20448 4862 20460
rect 12636 20457 12664 20488
rect 16482 20476 16488 20488
rect 16540 20476 16546 20528
rect 6825 20451 6883 20457
rect 6825 20448 6837 20451
rect 4856 20420 6837 20448
rect 4856 20408 4862 20420
rect 6825 20417 6837 20420
rect 6871 20448 6883 20451
rect 7653 20451 7711 20457
rect 7653 20448 7665 20451
rect 6871 20420 7665 20448
rect 6871 20417 6883 20420
rect 6825 20411 6883 20417
rect 7653 20417 7665 20420
rect 7699 20417 7711 20451
rect 7653 20411 7711 20417
rect 12621 20451 12679 20457
rect 12621 20417 12633 20451
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 12877 20451 12935 20457
rect 12877 20448 12889 20451
rect 12768 20420 12889 20448
rect 12768 20408 12774 20420
rect 12877 20417 12889 20420
rect 12923 20417 12935 20451
rect 12877 20411 12935 20417
rect 13354 20408 13360 20460
rect 13412 20448 13418 20460
rect 15197 20451 15255 20457
rect 15197 20448 15209 20451
rect 13412 20420 15209 20448
rect 13412 20408 13418 20420
rect 15197 20417 15209 20420
rect 15243 20417 15255 20451
rect 15197 20411 15255 20417
rect 15746 20408 15752 20460
rect 15804 20448 15810 20460
rect 17788 20457 17816 20556
rect 18782 20516 18788 20528
rect 17880 20488 18788 20516
rect 17037 20451 17095 20457
rect 17037 20448 17049 20451
rect 15804 20420 17049 20448
rect 15804 20408 15810 20420
rect 17037 20417 17049 20420
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 17773 20451 17831 20457
rect 17773 20417 17785 20451
rect 17819 20417 17831 20451
rect 17773 20411 17831 20417
rect 15473 20383 15531 20389
rect 15473 20349 15485 20383
rect 15519 20349 15531 20383
rect 17052 20380 17080 20411
rect 17880 20380 17908 20488
rect 18782 20476 18788 20488
rect 18840 20516 18846 20528
rect 19337 20519 19395 20525
rect 19337 20516 19349 20519
rect 18840 20488 19349 20516
rect 18840 20476 18846 20488
rect 19337 20485 19349 20488
rect 19383 20485 19395 20519
rect 20806 20516 20812 20528
rect 19337 20479 19395 20485
rect 19628 20488 20812 20516
rect 17957 20451 18015 20457
rect 17957 20417 17969 20451
rect 18003 20438 18015 20451
rect 19148 20451 19206 20457
rect 18003 20417 18092 20438
rect 17957 20411 18092 20417
rect 19148 20417 19160 20451
rect 19194 20417 19206 20451
rect 19148 20411 19206 20417
rect 17972 20410 18092 20411
rect 17052 20352 17908 20380
rect 18064 20380 18092 20410
rect 19163 20380 19191 20411
rect 19242 20408 19248 20460
rect 19300 20448 19306 20460
rect 19300 20420 19345 20448
rect 19300 20408 19306 20420
rect 19426 20408 19432 20460
rect 19484 20457 19490 20460
rect 19628 20457 19656 20488
rect 20806 20476 20812 20488
rect 20864 20476 20870 20528
rect 22572 20516 22600 20556
rect 22646 20544 22652 20596
rect 22704 20584 22710 20596
rect 23106 20584 23112 20596
rect 22704 20556 23112 20584
rect 22704 20544 22710 20556
rect 23106 20544 23112 20556
rect 23164 20544 23170 20596
rect 26970 20584 26976 20596
rect 23216 20556 26188 20584
rect 26931 20556 26976 20584
rect 23216 20516 23244 20556
rect 22572 20488 23244 20516
rect 25222 20476 25228 20528
rect 25280 20516 25286 20528
rect 26053 20519 26111 20525
rect 26053 20516 26065 20519
rect 25280 20488 26065 20516
rect 25280 20476 25286 20488
rect 26053 20485 26065 20488
rect 26099 20485 26111 20519
rect 26160 20516 26188 20556
rect 26970 20544 26976 20556
rect 27028 20544 27034 20596
rect 29730 20584 29736 20596
rect 29691 20556 29736 20584
rect 29730 20544 29736 20556
rect 29788 20544 29794 20596
rect 30193 20587 30251 20593
rect 30193 20553 30205 20587
rect 30239 20553 30251 20587
rect 36906 20584 36912 20596
rect 30193 20547 30251 20553
rect 30392 20556 36912 20584
rect 30208 20516 30236 20547
rect 26160 20488 30236 20516
rect 26053 20479 26111 20485
rect 19484 20451 19523 20457
rect 19511 20417 19523 20451
rect 19484 20411 19523 20417
rect 19613 20451 19671 20457
rect 19613 20417 19625 20451
rect 19659 20417 19671 20451
rect 19613 20411 19671 20417
rect 20252 20451 20310 20457
rect 20252 20417 20264 20451
rect 20298 20417 20310 20451
rect 20252 20411 20310 20417
rect 20349 20451 20407 20457
rect 20349 20417 20361 20451
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 19484 20408 19490 20411
rect 20162 20380 20168 20392
rect 18064 20352 19012 20380
rect 15473 20343 15531 20349
rect 15488 20312 15516 20343
rect 15562 20312 15568 20324
rect 15475 20284 15568 20312
rect 15562 20272 15568 20284
rect 15620 20312 15626 20324
rect 17954 20312 17960 20324
rect 15620 20284 17960 20312
rect 15620 20272 15626 20284
rect 17954 20272 17960 20284
rect 18012 20272 18018 20324
rect 18984 20321 19012 20352
rect 19076 20352 19191 20380
rect 19251 20352 20168 20380
rect 18969 20315 19027 20321
rect 18969 20281 18981 20315
rect 19015 20281 19027 20315
rect 19076 20312 19104 20352
rect 19251 20312 19279 20352
rect 20162 20340 20168 20352
rect 20220 20380 20226 20392
rect 20267 20380 20295 20411
rect 20220 20352 20295 20380
rect 20364 20380 20392 20411
rect 20438 20408 20444 20460
rect 20496 20448 20502 20460
rect 20622 20448 20628 20460
rect 20496 20420 20541 20448
rect 20583 20420 20628 20448
rect 20496 20408 20502 20420
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 20717 20451 20775 20457
rect 20717 20417 20729 20451
rect 20763 20448 20775 20451
rect 20898 20448 20904 20460
rect 20763 20420 20904 20448
rect 20763 20417 20775 20420
rect 20717 20411 20775 20417
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 22094 20448 22100 20460
rect 22055 20420 22100 20448
rect 22094 20408 22100 20420
rect 22152 20408 22158 20460
rect 23106 20448 23112 20460
rect 23067 20420 23112 20448
rect 23106 20408 23112 20420
rect 23164 20408 23170 20460
rect 23382 20457 23388 20460
rect 23376 20448 23388 20457
rect 23343 20420 23388 20448
rect 23376 20411 23388 20420
rect 23382 20408 23388 20411
rect 23440 20408 23446 20460
rect 23842 20408 23848 20460
rect 23900 20448 23906 20460
rect 25866 20448 25872 20460
rect 23900 20420 25872 20448
rect 23900 20408 23906 20420
rect 25866 20408 25872 20420
rect 25924 20408 25930 20460
rect 27062 20408 27068 20460
rect 27120 20448 27126 20460
rect 27246 20448 27252 20460
rect 27120 20420 27252 20448
rect 27120 20408 27126 20420
rect 27246 20408 27252 20420
rect 27304 20408 27310 20460
rect 27341 20451 27399 20457
rect 27341 20417 27353 20451
rect 27387 20417 27399 20451
rect 27341 20411 27399 20417
rect 27433 20451 27491 20457
rect 27433 20417 27445 20451
rect 27479 20448 27491 20451
rect 27617 20451 27675 20457
rect 27479 20420 27568 20448
rect 27479 20417 27491 20420
rect 27433 20411 27491 20417
rect 21910 20380 21916 20392
rect 20364 20352 21916 20380
rect 20220 20340 20226 20352
rect 21910 20340 21916 20352
rect 21968 20340 21974 20392
rect 20438 20312 20444 20324
rect 19076 20284 19279 20312
rect 19904 20284 20444 20312
rect 18969 20275 19027 20281
rect 19904 20256 19932 20284
rect 20438 20272 20444 20284
rect 20496 20272 20502 20324
rect 26878 20272 26884 20324
rect 26936 20312 26942 20324
rect 27356 20312 27384 20411
rect 27430 20312 27436 20324
rect 26936 20284 27436 20312
rect 26936 20272 26942 20284
rect 27430 20272 27436 20284
rect 27488 20272 27494 20324
rect 7926 20204 7932 20256
rect 7984 20244 7990 20256
rect 8297 20247 8355 20253
rect 8297 20244 8309 20247
rect 7984 20216 8309 20244
rect 7984 20204 7990 20216
rect 8297 20213 8309 20216
rect 8343 20244 8355 20247
rect 8386 20244 8392 20256
rect 8343 20216 8392 20244
rect 8343 20213 8355 20216
rect 8297 20207 8355 20213
rect 8386 20204 8392 20216
rect 8444 20204 8450 20256
rect 17586 20244 17592 20256
rect 17547 20216 17592 20244
rect 17586 20204 17592 20216
rect 17644 20204 17650 20256
rect 17862 20244 17868 20256
rect 17823 20216 17868 20244
rect 17862 20204 17868 20216
rect 17920 20204 17926 20256
rect 18782 20204 18788 20256
rect 18840 20244 18846 20256
rect 19886 20244 19892 20256
rect 18840 20216 19892 20244
rect 18840 20204 18846 20216
rect 19886 20204 19892 20216
rect 19944 20204 19950 20256
rect 20070 20244 20076 20256
rect 20031 20216 20076 20244
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 24489 20247 24547 20253
rect 24489 20213 24501 20247
rect 24535 20244 24547 20247
rect 24578 20244 24584 20256
rect 24535 20216 24584 20244
rect 24535 20213 24547 20216
rect 24489 20207 24547 20213
rect 24578 20204 24584 20216
rect 24636 20204 24642 20256
rect 26237 20247 26295 20253
rect 26237 20213 26249 20247
rect 26283 20244 26295 20247
rect 27540 20244 27568 20420
rect 27617 20417 27629 20451
rect 27663 20448 27675 20451
rect 27890 20448 27896 20460
rect 27663 20420 27896 20448
rect 27663 20417 27675 20420
rect 27617 20411 27675 20417
rect 27890 20408 27896 20420
rect 27948 20408 27954 20460
rect 28626 20408 28632 20460
rect 28684 20448 28690 20460
rect 29181 20451 29239 20457
rect 29181 20448 29193 20451
rect 28684 20420 29193 20448
rect 28684 20408 28690 20420
rect 29181 20417 29193 20420
rect 29227 20417 29239 20451
rect 29362 20448 29368 20460
rect 29323 20420 29368 20448
rect 29181 20411 29239 20417
rect 29362 20408 29368 20420
rect 29420 20408 29426 20460
rect 29457 20451 29515 20457
rect 29457 20417 29469 20451
rect 29503 20417 29515 20451
rect 29457 20411 29515 20417
rect 29472 20312 29500 20411
rect 29546 20408 29552 20460
rect 29604 20448 29610 20460
rect 30392 20457 30420 20556
rect 36906 20544 36912 20556
rect 36964 20544 36970 20596
rect 37274 20584 37280 20596
rect 37235 20556 37280 20584
rect 37274 20544 37280 20556
rect 37332 20544 37338 20596
rect 38289 20587 38347 20593
rect 38289 20584 38301 20587
rect 37568 20556 38301 20584
rect 30650 20516 30656 20528
rect 30611 20488 30656 20516
rect 30650 20476 30656 20488
rect 30708 20476 30714 20528
rect 33045 20519 33103 20525
rect 33045 20485 33057 20519
rect 33091 20516 33103 20519
rect 34618 20519 34676 20525
rect 34618 20516 34630 20519
rect 33091 20488 34630 20516
rect 33091 20485 33103 20488
rect 33045 20479 33103 20485
rect 34618 20485 34630 20488
rect 34664 20485 34676 20519
rect 34618 20479 34676 20485
rect 30377 20451 30435 20457
rect 29604 20420 29649 20448
rect 29604 20408 29610 20420
rect 30377 20417 30389 20451
rect 30423 20417 30435 20451
rect 30377 20411 30435 20417
rect 32306 20408 32312 20460
rect 32364 20448 32370 20460
rect 32401 20451 32459 20457
rect 32401 20448 32413 20451
rect 32364 20420 32413 20448
rect 32364 20408 32370 20420
rect 32401 20417 32413 20420
rect 32447 20417 32459 20451
rect 32401 20411 32459 20417
rect 32585 20451 32643 20457
rect 32585 20417 32597 20451
rect 32631 20417 32643 20451
rect 32585 20411 32643 20417
rect 30466 20380 30472 20392
rect 30427 20352 30472 20380
rect 30466 20340 30472 20352
rect 30524 20340 30530 20392
rect 32600 20312 32628 20411
rect 32674 20408 32680 20460
rect 32732 20448 32738 20460
rect 32858 20457 32864 20460
rect 32815 20451 32864 20457
rect 32732 20420 32777 20448
rect 32732 20408 32738 20420
rect 32815 20417 32827 20451
rect 32861 20417 32864 20451
rect 32815 20411 32864 20417
rect 32858 20408 32864 20411
rect 32916 20408 32922 20460
rect 34885 20451 34943 20457
rect 34885 20417 34897 20451
rect 34931 20417 34943 20451
rect 34885 20411 34943 20417
rect 36173 20451 36231 20457
rect 36173 20417 36185 20451
rect 36219 20448 36231 20451
rect 36262 20448 36268 20460
rect 36219 20420 36268 20448
rect 36219 20417 36231 20420
rect 36173 20411 36231 20417
rect 33042 20312 33048 20324
rect 29472 20284 31754 20312
rect 32600 20284 33048 20312
rect 26283 20216 27568 20244
rect 26283 20213 26295 20216
rect 26237 20207 26295 20213
rect 27890 20204 27896 20256
rect 27948 20244 27954 20256
rect 28258 20244 28264 20256
rect 27948 20216 28264 20244
rect 27948 20204 27954 20216
rect 28258 20204 28264 20216
rect 28316 20244 28322 20256
rect 28353 20247 28411 20253
rect 28353 20244 28365 20247
rect 28316 20216 28365 20244
rect 28316 20204 28322 20216
rect 28353 20213 28365 20216
rect 28399 20213 28411 20247
rect 30374 20244 30380 20256
rect 30335 20216 30380 20244
rect 28353 20207 28411 20213
rect 30374 20204 30380 20216
rect 30432 20204 30438 20256
rect 31726 20244 31754 20284
rect 33042 20272 33048 20284
rect 33100 20272 33106 20324
rect 32858 20244 32864 20256
rect 31726 20216 32864 20244
rect 32858 20204 32864 20216
rect 32916 20244 32922 20256
rect 33505 20247 33563 20253
rect 33505 20244 33517 20247
rect 32916 20216 33517 20244
rect 32916 20204 32922 20216
rect 33505 20213 33517 20216
rect 33551 20213 33563 20247
rect 33505 20207 33563 20213
rect 34238 20204 34244 20256
rect 34296 20244 34302 20256
rect 34900 20244 34928 20411
rect 36262 20408 36268 20420
rect 36320 20408 36326 20460
rect 37182 20408 37188 20460
rect 37240 20448 37246 20460
rect 37568 20457 37596 20556
rect 38289 20553 38301 20556
rect 38335 20584 38347 20587
rect 38335 20556 40356 20584
rect 38335 20553 38347 20556
rect 38289 20547 38347 20553
rect 40328 20525 40356 20556
rect 40313 20519 40371 20525
rect 40313 20485 40325 20519
rect 40359 20485 40371 20519
rect 40313 20479 40371 20485
rect 37461 20451 37519 20457
rect 37461 20448 37473 20451
rect 37240 20420 37473 20448
rect 37240 20408 37246 20420
rect 37461 20417 37473 20420
rect 37507 20417 37519 20451
rect 37461 20411 37519 20417
rect 37553 20451 37611 20457
rect 37553 20417 37565 20451
rect 37599 20417 37611 20451
rect 37553 20411 37611 20417
rect 37645 20451 37703 20457
rect 37645 20417 37657 20451
rect 37691 20417 37703 20451
rect 37826 20448 37832 20460
rect 37787 20420 37832 20448
rect 37645 20411 37703 20417
rect 35897 20383 35955 20389
rect 35897 20349 35909 20383
rect 35943 20380 35955 20383
rect 37090 20380 37096 20392
rect 35943 20352 37096 20380
rect 35943 20349 35955 20352
rect 35897 20343 35955 20349
rect 37090 20340 37096 20352
rect 37148 20380 37154 20392
rect 37660 20380 37688 20411
rect 37826 20408 37832 20420
rect 37884 20408 37890 20460
rect 39413 20451 39471 20457
rect 39413 20417 39425 20451
rect 39459 20448 39471 20451
rect 39574 20448 39580 20460
rect 39459 20420 39580 20448
rect 39459 20417 39471 20420
rect 39413 20411 39471 20417
rect 39574 20408 39580 20420
rect 39632 20408 39638 20460
rect 39758 20408 39764 20460
rect 39816 20448 39822 20460
rect 40129 20451 40187 20457
rect 40129 20448 40141 20451
rect 39816 20420 40141 20448
rect 39816 20408 39822 20420
rect 40129 20417 40141 20420
rect 40175 20417 40187 20451
rect 40129 20411 40187 20417
rect 37148 20352 37688 20380
rect 39669 20383 39727 20389
rect 37148 20340 37154 20352
rect 39669 20349 39681 20383
rect 39715 20380 39727 20383
rect 39942 20380 39948 20392
rect 39715 20352 39948 20380
rect 39715 20349 39727 20352
rect 39669 20343 39727 20349
rect 39684 20244 39712 20343
rect 39942 20340 39948 20352
rect 40000 20340 40006 20392
rect 34296 20216 39712 20244
rect 40497 20247 40555 20253
rect 34296 20204 34302 20216
rect 40497 20213 40509 20247
rect 40543 20244 40555 20247
rect 40678 20244 40684 20256
rect 40543 20216 40684 20244
rect 40543 20213 40555 20216
rect 40497 20207 40555 20213
rect 40678 20204 40684 20216
rect 40736 20204 40742 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 7190 20000 7196 20052
rect 7248 20040 7254 20052
rect 7285 20043 7343 20049
rect 7285 20040 7297 20043
rect 7248 20012 7297 20040
rect 7248 20000 7254 20012
rect 7285 20009 7297 20012
rect 7331 20009 7343 20043
rect 12710 20040 12716 20052
rect 12671 20012 12716 20040
rect 7285 20003 7343 20009
rect 12710 20000 12716 20012
rect 12768 20000 12774 20052
rect 15562 20040 15568 20052
rect 15523 20012 15568 20040
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 21821 20043 21879 20049
rect 21821 20009 21833 20043
rect 21867 20040 21879 20043
rect 22094 20040 22100 20052
rect 21867 20012 22100 20040
rect 21867 20009 21879 20012
rect 21821 20003 21879 20009
rect 22094 20000 22100 20012
rect 22152 20040 22158 20052
rect 23566 20040 23572 20052
rect 22152 20012 23572 20040
rect 22152 20000 22158 20012
rect 23566 20000 23572 20012
rect 23624 20000 23630 20052
rect 33042 20040 33048 20052
rect 33003 20012 33048 20040
rect 33042 20000 33048 20012
rect 33100 20000 33106 20052
rect 36906 20000 36912 20052
rect 36964 20040 36970 20052
rect 37553 20043 37611 20049
rect 37553 20040 37565 20043
rect 36964 20012 37565 20040
rect 36964 20000 36970 20012
rect 37553 20009 37565 20012
rect 37599 20009 37611 20043
rect 37553 20003 37611 20009
rect 39574 20000 39580 20052
rect 39632 20040 39638 20052
rect 40221 20043 40279 20049
rect 40221 20040 40233 20043
rect 39632 20012 40233 20040
rect 39632 20000 39638 20012
rect 40221 20009 40233 20012
rect 40267 20009 40279 20043
rect 40221 20003 40279 20009
rect 3234 19932 3240 19984
rect 3292 19972 3298 19984
rect 4617 19975 4675 19981
rect 4617 19972 4629 19975
rect 3292 19944 4629 19972
rect 3292 19932 3298 19944
rect 4617 19941 4629 19944
rect 4663 19972 4675 19975
rect 9398 19972 9404 19984
rect 4663 19944 9404 19972
rect 4663 19941 4675 19944
rect 4617 19935 4675 19941
rect 9398 19932 9404 19944
rect 9456 19932 9462 19984
rect 18046 19932 18052 19984
rect 18104 19972 18110 19984
rect 26326 19972 26332 19984
rect 18104 19944 26332 19972
rect 18104 19932 18110 19944
rect 26326 19932 26332 19944
rect 26384 19932 26390 19984
rect 27154 19932 27160 19984
rect 27212 19972 27218 19984
rect 36722 19972 36728 19984
rect 27212 19944 36728 19972
rect 27212 19932 27218 19944
rect 36722 19932 36728 19944
rect 36780 19932 36786 19984
rect 12434 19904 12440 19916
rect 11624 19876 12440 19904
rect 2590 19836 2596 19848
rect 2551 19808 2596 19836
rect 2590 19796 2596 19808
rect 2648 19796 2654 19848
rect 4433 19839 4491 19845
rect 4433 19805 4445 19839
rect 4479 19836 4491 19839
rect 4798 19836 4804 19848
rect 4479 19808 4804 19836
rect 4479 19805 4491 19808
rect 4433 19799 4491 19805
rect 4798 19796 4804 19808
rect 4856 19796 4862 19848
rect 8294 19796 8300 19848
rect 8352 19836 8358 19848
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 8352 19808 9413 19836
rect 8352 19796 8358 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 11330 19796 11336 19848
rect 11388 19836 11394 19848
rect 11624 19845 11652 19876
rect 12434 19864 12440 19876
rect 12492 19904 12498 19916
rect 14369 19907 14427 19913
rect 14369 19904 14381 19907
rect 12492 19876 14381 19904
rect 12492 19864 12498 19876
rect 11517 19839 11575 19845
rect 11517 19836 11529 19839
rect 11388 19808 11529 19836
rect 11388 19796 11394 19808
rect 11517 19805 11529 19808
rect 11563 19805 11575 19839
rect 11517 19799 11575 19805
rect 11609 19839 11667 19845
rect 11609 19805 11621 19839
rect 11655 19805 11667 19839
rect 11609 19799 11667 19805
rect 11698 19796 11704 19848
rect 11756 19836 11762 19848
rect 11756 19808 11801 19836
rect 11756 19796 11762 19808
rect 11882 19796 11888 19848
rect 11940 19836 11946 19848
rect 12158 19836 12164 19848
rect 11940 19808 12164 19836
rect 11940 19796 11946 19808
rect 12158 19796 12164 19808
rect 12216 19796 12222 19848
rect 12710 19796 12716 19848
rect 12768 19836 12774 19848
rect 13096 19845 13124 19876
rect 14369 19873 14381 19876
rect 14415 19873 14427 19907
rect 16114 19904 16120 19916
rect 14369 19867 14427 19873
rect 15580 19876 16120 19904
rect 12989 19839 13047 19845
rect 12989 19836 13001 19839
rect 12768 19808 13001 19836
rect 12768 19796 12774 19808
rect 12989 19805 13001 19808
rect 13035 19805 13047 19839
rect 12989 19799 13047 19805
rect 13081 19839 13139 19845
rect 13081 19805 13093 19839
rect 13127 19805 13139 19839
rect 13081 19799 13139 19805
rect 13173 19839 13231 19845
rect 13173 19805 13185 19839
rect 13219 19836 13231 19839
rect 13262 19836 13268 19848
rect 13219 19808 13268 19836
rect 13219 19805 13231 19808
rect 13173 19799 13231 19805
rect 13262 19796 13268 19808
rect 13320 19796 13326 19848
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19836 13415 19839
rect 13446 19836 13452 19848
rect 13403 19808 13452 19836
rect 13403 19805 13415 19808
rect 13357 19799 13415 19805
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19836 14151 19839
rect 14182 19836 14188 19848
rect 14139 19808 14188 19836
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 14182 19796 14188 19808
rect 14240 19836 14246 19848
rect 15580 19836 15608 19876
rect 16114 19864 16120 19876
rect 16172 19864 16178 19916
rect 20346 19904 20352 19916
rect 19720 19876 20352 19904
rect 15746 19836 15752 19848
rect 14240 19808 15608 19836
rect 15707 19808 15752 19836
rect 14240 19796 14246 19808
rect 15746 19796 15752 19808
rect 15804 19796 15810 19848
rect 15838 19796 15844 19848
rect 15896 19836 15902 19848
rect 19720 19845 19748 19876
rect 20346 19864 20352 19876
rect 20404 19864 20410 19916
rect 22373 19907 22431 19913
rect 22373 19904 22385 19907
rect 21744 19876 22385 19904
rect 19705 19839 19763 19845
rect 15896 19808 15941 19836
rect 15896 19796 15902 19808
rect 19705 19805 19717 19839
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 19798 19839 19856 19845
rect 19798 19805 19810 19839
rect 19844 19805 19856 19839
rect 19798 19799 19856 19805
rect 5994 19728 6000 19780
rect 6052 19768 6058 19780
rect 6641 19771 6699 19777
rect 6641 19768 6653 19771
rect 6052 19740 6653 19768
rect 6052 19728 6058 19740
rect 6641 19737 6653 19740
rect 6687 19768 6699 19771
rect 7561 19771 7619 19777
rect 7561 19768 7573 19771
rect 6687 19740 7573 19768
rect 6687 19737 6699 19740
rect 6641 19731 6699 19737
rect 7561 19737 7573 19740
rect 7607 19737 7619 19771
rect 7561 19731 7619 19737
rect 9668 19771 9726 19777
rect 9668 19737 9680 19771
rect 9714 19768 9726 19771
rect 11241 19771 11299 19777
rect 11241 19768 11253 19771
rect 9714 19740 11253 19768
rect 9714 19737 9726 19740
rect 9668 19731 9726 19737
rect 11241 19737 11253 19740
rect 11287 19737 11299 19771
rect 11241 19731 11299 19737
rect 19334 19728 19340 19780
rect 19392 19768 19398 19780
rect 19812 19768 19840 19799
rect 19886 19796 19892 19848
rect 19944 19836 19950 19848
rect 19981 19839 20039 19845
rect 19981 19836 19993 19839
rect 19944 19808 19993 19836
rect 19944 19796 19950 19808
rect 19981 19805 19993 19808
rect 20027 19805 20039 19839
rect 19981 19799 20039 19805
rect 20162 19796 20168 19848
rect 20220 19845 20226 19848
rect 20220 19836 20228 19845
rect 20220 19808 20265 19836
rect 20220 19799 20228 19808
rect 20220 19796 20226 19799
rect 21174 19796 21180 19848
rect 21232 19836 21238 19848
rect 21744 19845 21772 19876
rect 22373 19873 22385 19876
rect 22419 19873 22431 19907
rect 29914 19904 29920 19916
rect 29827 19876 29920 19904
rect 22373 19867 22431 19873
rect 29914 19864 29920 19876
rect 29972 19904 29978 19916
rect 30834 19904 30840 19916
rect 29972 19876 30840 19904
rect 29972 19864 29978 19876
rect 30834 19864 30840 19876
rect 30892 19904 30898 19916
rect 31386 19904 31392 19916
rect 30892 19876 31392 19904
rect 30892 19864 30898 19876
rect 31386 19864 31392 19876
rect 31444 19864 31450 19916
rect 35986 19864 35992 19916
rect 36044 19904 36050 19916
rect 36541 19907 36599 19913
rect 36541 19904 36553 19907
rect 36044 19876 36553 19904
rect 36044 19864 36050 19876
rect 36541 19873 36553 19876
rect 36587 19873 36599 19907
rect 36541 19867 36599 19873
rect 40402 19864 40408 19916
rect 40460 19904 40466 19916
rect 40770 19904 40776 19916
rect 40460 19876 40776 19904
rect 40460 19864 40466 19876
rect 21729 19839 21787 19845
rect 21729 19836 21741 19839
rect 21232 19808 21741 19836
rect 21232 19796 21238 19808
rect 21729 19805 21741 19808
rect 21775 19805 21787 19839
rect 21729 19799 21787 19805
rect 21913 19839 21971 19845
rect 21913 19805 21925 19839
rect 21959 19836 21971 19839
rect 21959 19808 22094 19836
rect 21959 19805 21971 19808
rect 21913 19799 21971 19805
rect 19392 19740 19840 19768
rect 20073 19771 20131 19777
rect 19392 19728 19398 19740
rect 20073 19737 20085 19771
rect 20119 19768 20131 19771
rect 20714 19768 20720 19780
rect 20119 19740 20720 19768
rect 20119 19737 20131 19740
rect 20073 19731 20131 19737
rect 20714 19728 20720 19740
rect 20772 19728 20778 19780
rect 22066 19768 22094 19808
rect 22186 19796 22192 19848
rect 22244 19836 22250 19848
rect 24394 19836 24400 19848
rect 22244 19808 24400 19836
rect 22244 19796 22250 19808
rect 24394 19796 24400 19808
rect 24452 19796 24458 19848
rect 25682 19796 25688 19848
rect 25740 19836 25746 19848
rect 28810 19836 28816 19848
rect 25740 19808 28816 19836
rect 25740 19796 25746 19808
rect 28810 19796 28816 19808
rect 28868 19836 28874 19848
rect 29546 19836 29552 19848
rect 28868 19808 29552 19836
rect 28868 19796 28874 19808
rect 29546 19796 29552 19808
rect 29604 19836 29610 19848
rect 29641 19839 29699 19845
rect 29641 19836 29653 19839
rect 29604 19808 29653 19836
rect 29604 19796 29610 19808
rect 29641 19805 29653 19808
rect 29687 19805 29699 19839
rect 29641 19799 29699 19805
rect 31938 19796 31944 19848
rect 31996 19836 32002 19848
rect 32677 19839 32735 19845
rect 32677 19836 32689 19839
rect 31996 19808 32689 19836
rect 31996 19796 32002 19808
rect 32677 19805 32689 19808
rect 32723 19805 32735 19839
rect 32858 19836 32864 19848
rect 32819 19808 32864 19836
rect 32677 19799 32735 19805
rect 32858 19796 32864 19808
rect 32916 19796 32922 19848
rect 36265 19839 36323 19845
rect 36265 19805 36277 19839
rect 36311 19836 36323 19839
rect 37182 19836 37188 19848
rect 36311 19808 37188 19836
rect 36311 19805 36323 19808
rect 36265 19799 36323 19805
rect 37182 19796 37188 19808
rect 37240 19836 37246 19848
rect 37737 19839 37795 19845
rect 37737 19836 37749 19839
rect 37240 19808 37749 19836
rect 37240 19796 37246 19808
rect 37737 19805 37749 19808
rect 37783 19805 37795 19839
rect 37737 19799 37795 19805
rect 37829 19839 37887 19845
rect 37829 19805 37841 19839
rect 37875 19836 37887 19839
rect 38105 19839 38163 19845
rect 37875 19808 38056 19836
rect 37875 19805 37887 19808
rect 37829 19799 37887 19805
rect 22370 19768 22376 19780
rect 22066 19740 22376 19768
rect 22370 19728 22376 19740
rect 22428 19728 22434 19780
rect 27430 19768 27436 19780
rect 27391 19740 27436 19768
rect 27430 19728 27436 19740
rect 27488 19728 27494 19780
rect 37090 19728 37096 19780
rect 37148 19768 37154 19780
rect 37921 19771 37979 19777
rect 37921 19768 37933 19771
rect 37148 19740 37933 19768
rect 37148 19728 37154 19740
rect 37921 19737 37933 19740
rect 37967 19737 37979 19771
rect 38028 19768 38056 19808
rect 38105 19805 38117 19839
rect 38151 19836 38163 19839
rect 38746 19836 38752 19848
rect 38151 19808 38752 19836
rect 38151 19805 38163 19808
rect 38105 19799 38163 19805
rect 38746 19796 38752 19808
rect 38804 19796 38810 19848
rect 40034 19796 40040 19848
rect 40092 19836 40098 19848
rect 40604 19845 40632 19876
rect 40770 19864 40776 19876
rect 40828 19864 40834 19916
rect 40497 19839 40555 19845
rect 40497 19836 40509 19839
rect 40092 19808 40509 19836
rect 40092 19796 40098 19808
rect 40497 19805 40509 19808
rect 40543 19805 40555 19839
rect 40497 19799 40555 19805
rect 40589 19839 40647 19845
rect 40589 19805 40601 19839
rect 40635 19805 40647 19839
rect 40589 19799 40647 19805
rect 40678 19796 40684 19848
rect 40736 19836 40742 19848
rect 40865 19839 40923 19845
rect 40736 19808 40781 19836
rect 40736 19796 40742 19808
rect 40865 19805 40877 19839
rect 40911 19836 40923 19839
rect 41138 19836 41144 19848
rect 40911 19808 41144 19836
rect 40911 19805 40923 19808
rect 40865 19799 40923 19805
rect 41138 19796 41144 19808
rect 41196 19796 41202 19848
rect 58158 19836 58164 19848
rect 58119 19808 58164 19836
rect 58158 19796 58164 19808
rect 58216 19796 58222 19848
rect 41690 19768 41696 19780
rect 38028 19740 41696 19768
rect 37921 19731 37979 19737
rect 41690 19728 41696 19740
rect 41748 19728 41754 19780
rect 2406 19700 2412 19712
rect 2367 19672 2412 19700
rect 2406 19660 2412 19672
rect 2464 19660 2470 19712
rect 5626 19700 5632 19712
rect 5587 19672 5632 19700
rect 5626 19660 5632 19672
rect 5684 19660 5690 19712
rect 5902 19660 5908 19712
rect 5960 19700 5966 19712
rect 6089 19703 6147 19709
rect 6089 19700 6101 19703
rect 5960 19672 6101 19700
rect 5960 19660 5966 19672
rect 6089 19669 6101 19672
rect 6135 19669 6147 19703
rect 8386 19700 8392 19712
rect 8347 19672 8392 19700
rect 6089 19663 6147 19669
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 10502 19660 10508 19712
rect 10560 19700 10566 19712
rect 10781 19703 10839 19709
rect 10781 19700 10793 19703
rect 10560 19672 10793 19700
rect 10560 19660 10566 19672
rect 10781 19669 10793 19672
rect 10827 19669 10839 19703
rect 10781 19663 10839 19669
rect 11330 19660 11336 19712
rect 11388 19700 11394 19712
rect 13906 19700 13912 19712
rect 11388 19672 13912 19700
rect 11388 19660 11394 19672
rect 13906 19660 13912 19672
rect 13964 19660 13970 19712
rect 20346 19700 20352 19712
rect 20307 19672 20352 19700
rect 20346 19660 20352 19672
rect 20404 19660 20410 19712
rect 26145 19703 26203 19709
rect 26145 19669 26157 19703
rect 26191 19700 26203 19703
rect 26602 19700 26608 19712
rect 26191 19672 26608 19700
rect 26191 19669 26203 19672
rect 26145 19663 26203 19669
rect 26602 19660 26608 19672
rect 26660 19700 26666 19712
rect 27246 19700 27252 19712
rect 26660 19672 27252 19700
rect 26660 19660 26666 19672
rect 27246 19660 27252 19672
rect 27304 19660 27310 19712
rect 27890 19700 27896 19712
rect 27851 19672 27896 19700
rect 27890 19660 27896 19672
rect 27948 19660 27954 19712
rect 32214 19660 32220 19712
rect 32272 19700 32278 19712
rect 39209 19703 39267 19709
rect 39209 19700 39221 19703
rect 32272 19672 39221 19700
rect 32272 19660 32278 19672
rect 39209 19669 39221 19672
rect 39255 19700 39267 19703
rect 40034 19700 40040 19712
rect 39255 19672 40040 19700
rect 39255 19669 39267 19672
rect 39209 19663 39267 19669
rect 40034 19660 40040 19672
rect 40092 19660 40098 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 5169 19499 5227 19505
rect 5169 19465 5181 19499
rect 5215 19496 5227 19499
rect 5626 19496 5632 19508
rect 5215 19468 5632 19496
rect 5215 19465 5227 19468
rect 5169 19459 5227 19465
rect 5626 19456 5632 19468
rect 5684 19496 5690 19508
rect 5684 19468 7512 19496
rect 5684 19456 5690 19468
rect 5902 19388 5908 19440
rect 5960 19428 5966 19440
rect 7101 19431 7159 19437
rect 7101 19428 7113 19431
rect 5960 19400 7113 19428
rect 5960 19388 5966 19400
rect 7101 19397 7113 19400
rect 7147 19397 7159 19431
rect 7484 19428 7512 19468
rect 7558 19456 7564 19508
rect 7616 19496 7622 19508
rect 8665 19499 8723 19505
rect 8665 19496 8677 19499
rect 7616 19468 8677 19496
rect 7616 19456 7622 19468
rect 8665 19465 8677 19468
rect 8711 19465 8723 19499
rect 11330 19496 11336 19508
rect 8665 19459 8723 19465
rect 8956 19468 11336 19496
rect 7926 19428 7932 19440
rect 7484 19400 7932 19428
rect 7101 19391 7159 19397
rect 7926 19388 7932 19400
rect 7984 19388 7990 19440
rect 8570 19428 8576 19440
rect 8128 19400 8576 19428
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19360 4399 19363
rect 4614 19360 4620 19372
rect 4387 19332 4620 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 4614 19320 4620 19332
rect 4672 19320 4678 19372
rect 5258 19360 5264 19372
rect 5219 19332 5264 19360
rect 5258 19320 5264 19332
rect 5316 19320 5322 19372
rect 8128 19360 8156 19400
rect 8570 19388 8576 19400
rect 8628 19388 8634 19440
rect 7944 19332 8156 19360
rect 8205 19363 8263 19369
rect 4890 19252 4896 19304
rect 4948 19292 4954 19304
rect 5353 19295 5411 19301
rect 5353 19292 5365 19295
rect 4948 19264 5365 19292
rect 4948 19252 4954 19264
rect 5353 19261 5365 19264
rect 5399 19261 5411 19295
rect 5353 19255 5411 19261
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 7944 19292 7972 19332
rect 8205 19329 8217 19363
rect 8251 19360 8263 19363
rect 8956 19360 8984 19468
rect 11330 19456 11336 19468
rect 11388 19456 11394 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19496 11575 19499
rect 11698 19496 11704 19508
rect 11563 19468 11704 19496
rect 11563 19465 11575 19468
rect 11517 19459 11575 19465
rect 11698 19456 11704 19468
rect 11756 19456 11762 19508
rect 14182 19496 14188 19508
rect 14143 19468 14188 19496
rect 14182 19456 14188 19468
rect 14240 19456 14246 19508
rect 14366 19456 14372 19508
rect 14424 19456 14430 19508
rect 14829 19499 14887 19505
rect 14829 19465 14841 19499
rect 14875 19496 14887 19499
rect 14918 19496 14924 19508
rect 14875 19468 14924 19496
rect 14875 19465 14887 19468
rect 14829 19459 14887 19465
rect 14918 19456 14924 19468
rect 14976 19456 14982 19508
rect 21174 19496 21180 19508
rect 15120 19468 21180 19496
rect 13630 19428 13636 19440
rect 9048 19400 13636 19428
rect 9048 19369 9076 19400
rect 13630 19388 13636 19400
rect 13688 19388 13694 19440
rect 14384 19428 14412 19456
rect 15120 19428 15148 19468
rect 21174 19456 21180 19468
rect 21232 19456 21238 19508
rect 25823 19499 25881 19505
rect 25823 19465 25835 19499
rect 25869 19496 25881 19499
rect 26878 19496 26884 19508
rect 25869 19468 26884 19496
rect 25869 19465 25881 19468
rect 25823 19459 25881 19465
rect 26878 19456 26884 19468
rect 26936 19456 26942 19508
rect 26973 19499 27031 19505
rect 26973 19465 26985 19499
rect 27019 19496 27031 19499
rect 28997 19499 29055 19505
rect 27019 19468 27108 19496
rect 27019 19465 27031 19468
rect 26973 19459 27031 19465
rect 20070 19428 20076 19440
rect 14200 19400 15148 19428
rect 15212 19400 20076 19428
rect 8251 19332 8984 19360
rect 9033 19363 9091 19369
rect 8251 19329 8263 19332
rect 8205 19323 8263 19329
rect 9033 19329 9045 19363
rect 9079 19329 9091 19363
rect 9033 19323 9091 19329
rect 10502 19320 10508 19372
rect 10560 19360 10566 19372
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 10560 19332 11713 19360
rect 10560 19320 10566 19332
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 11885 19363 11943 19369
rect 11885 19329 11897 19363
rect 11931 19360 11943 19363
rect 12526 19360 12532 19372
rect 11931 19332 12532 19360
rect 11931 19329 11943 19332
rect 11885 19323 11943 19329
rect 12526 19320 12532 19332
rect 12584 19360 12590 19372
rect 13354 19360 13360 19372
rect 12584 19332 13360 19360
rect 12584 19320 12590 19332
rect 13354 19320 13360 19332
rect 13412 19320 13418 19372
rect 14200 19369 14228 19400
rect 14185 19363 14243 19369
rect 14185 19329 14197 19363
rect 14231 19329 14243 19363
rect 14185 19323 14243 19329
rect 14274 19320 14280 19372
rect 14332 19360 14338 19372
rect 15212 19369 15240 19400
rect 20070 19388 20076 19400
rect 20128 19388 20134 19440
rect 21910 19388 21916 19440
rect 21968 19428 21974 19440
rect 22005 19431 22063 19437
rect 22005 19428 22017 19431
rect 21968 19400 22017 19428
rect 21968 19388 21974 19400
rect 22005 19397 22017 19400
rect 22051 19397 22063 19431
rect 27080 19428 27108 19468
rect 28997 19465 29009 19499
rect 29043 19496 29055 19499
rect 30374 19496 30380 19508
rect 29043 19468 30380 19496
rect 29043 19465 29055 19468
rect 28997 19459 29055 19465
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 32677 19499 32735 19505
rect 30944 19468 31754 19496
rect 22005 19391 22063 19397
rect 24504 19400 27108 19428
rect 27433 19431 27491 19437
rect 14369 19363 14427 19369
rect 14369 19360 14381 19363
rect 14332 19332 14381 19360
rect 14332 19320 14338 19332
rect 14369 19329 14381 19332
rect 14415 19329 14427 19363
rect 14369 19323 14427 19329
rect 15197 19363 15255 19369
rect 15197 19329 15209 19363
rect 15243 19329 15255 19363
rect 15197 19323 15255 19329
rect 16482 19320 16488 19372
rect 16540 19360 16546 19372
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 16540 19332 16681 19360
rect 16540 19320 16546 19332
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 16758 19320 16764 19372
rect 16816 19360 16822 19372
rect 16925 19363 16983 19369
rect 16925 19360 16937 19363
rect 16816 19332 16937 19360
rect 16816 19320 16822 19332
rect 16925 19329 16937 19332
rect 16971 19329 16983 19363
rect 22186 19360 22192 19372
rect 16925 19323 16983 19329
rect 22066 19332 22192 19360
rect 8110 19292 8116 19304
rect 6871 19264 7972 19292
rect 8071 19264 8116 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 8110 19252 8116 19264
rect 8168 19292 8174 19304
rect 8386 19292 8392 19304
rect 8168 19264 8392 19292
rect 8168 19252 8174 19264
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 8941 19295 8999 19301
rect 8941 19261 8953 19295
rect 8987 19261 8999 19295
rect 8941 19255 8999 19261
rect 15105 19295 15163 19301
rect 15105 19261 15117 19295
rect 15151 19261 15163 19295
rect 15105 19255 15163 19261
rect 2866 19224 2872 19236
rect 2827 19196 2872 19224
rect 2866 19184 2872 19196
rect 2924 19184 2930 19236
rect 7650 19184 7656 19236
rect 7708 19224 7714 19236
rect 8956 19224 8984 19255
rect 9585 19227 9643 19233
rect 9585 19224 9597 19227
rect 7708 19196 8064 19224
rect 8956 19196 9597 19224
rect 7708 19184 7714 19196
rect 4798 19156 4804 19168
rect 4759 19128 4804 19156
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 7466 19116 7472 19168
rect 7524 19156 7530 19168
rect 8036 19165 8064 19196
rect 9585 19193 9597 19196
rect 9631 19224 9643 19227
rect 11698 19224 11704 19236
rect 9631 19196 11704 19224
rect 9631 19193 9643 19196
rect 9585 19187 9643 19193
rect 11698 19184 11704 19196
rect 11756 19184 11762 19236
rect 15120 19224 15148 19255
rect 21450 19252 21456 19304
rect 21508 19292 21514 19304
rect 22066 19292 22094 19332
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 21508 19264 22094 19292
rect 21508 19252 21514 19264
rect 24504 19224 24532 19400
rect 27433 19397 27445 19431
rect 27479 19428 27491 19431
rect 27522 19428 27528 19440
rect 27479 19400 27528 19428
rect 27479 19397 27491 19400
rect 27433 19391 27491 19397
rect 27522 19388 27528 19400
rect 27580 19388 27586 19440
rect 28721 19431 28779 19437
rect 28721 19397 28733 19431
rect 28767 19428 28779 19431
rect 30944 19428 30972 19468
rect 28767 19400 30972 19428
rect 31726 19428 31754 19468
rect 32677 19465 32689 19499
rect 32723 19465 32735 19499
rect 32677 19459 32735 19465
rect 32398 19428 32404 19440
rect 31726 19400 32404 19428
rect 28767 19397 28779 19400
rect 28721 19391 28779 19397
rect 32398 19388 32404 19400
rect 32456 19428 32462 19440
rect 32692 19428 32720 19459
rect 33778 19456 33784 19508
rect 33836 19496 33842 19508
rect 35989 19499 36047 19505
rect 35989 19496 36001 19499
rect 33836 19468 36001 19496
rect 33836 19456 33842 19468
rect 35989 19465 36001 19468
rect 36035 19465 36047 19499
rect 35989 19459 36047 19465
rect 36262 19456 36268 19508
rect 36320 19496 36326 19508
rect 39666 19496 39672 19508
rect 36320 19468 36400 19496
rect 36320 19456 36326 19468
rect 36372 19437 36400 19468
rect 36464 19468 39672 19496
rect 32456 19400 32720 19428
rect 36357 19431 36415 19437
rect 32456 19388 32462 19400
rect 36357 19397 36369 19431
rect 36403 19397 36415 19431
rect 36357 19391 36415 19397
rect 27154 19360 27160 19372
rect 27115 19332 27160 19360
rect 27154 19320 27160 19332
rect 27212 19320 27218 19372
rect 27338 19320 27344 19372
rect 27396 19360 27402 19372
rect 28445 19363 28503 19369
rect 28445 19360 28457 19363
rect 27396 19332 28457 19360
rect 27396 19320 27402 19332
rect 28445 19329 28457 19332
rect 28491 19329 28503 19363
rect 28629 19363 28687 19369
rect 28629 19360 28641 19363
rect 28445 19323 28503 19329
rect 28552 19332 28641 19360
rect 24670 19252 24676 19304
rect 24728 19292 24734 19304
rect 25593 19295 25651 19301
rect 25593 19292 25605 19295
rect 24728 19264 25605 19292
rect 24728 19252 24734 19264
rect 25593 19261 25605 19264
rect 25639 19261 25651 19295
rect 25593 19255 25651 19261
rect 26694 19252 26700 19304
rect 26752 19292 26758 19304
rect 27249 19295 27307 19301
rect 27249 19292 27261 19295
rect 26752 19264 27261 19292
rect 26752 19252 26758 19264
rect 27249 19261 27261 19264
rect 27295 19261 27307 19295
rect 27249 19255 27307 19261
rect 28350 19252 28356 19304
rect 28408 19292 28414 19304
rect 28552 19292 28580 19332
rect 28629 19329 28641 19332
rect 28675 19329 28687 19363
rect 28810 19360 28816 19372
rect 28771 19332 28816 19360
rect 28629 19323 28687 19329
rect 28810 19320 28816 19332
rect 28868 19320 28874 19372
rect 29457 19363 29515 19369
rect 29457 19329 29469 19363
rect 29503 19329 29515 19363
rect 29457 19323 29515 19329
rect 29362 19292 29368 19304
rect 28408 19264 29368 19292
rect 28408 19252 28414 19264
rect 29362 19252 29368 19264
rect 29420 19292 29426 19304
rect 29472 19292 29500 19323
rect 30834 19320 30840 19372
rect 30892 19369 30898 19372
rect 30892 19363 30941 19369
rect 30892 19329 30895 19363
rect 30929 19329 30941 19363
rect 30892 19323 30941 19329
rect 31021 19363 31079 19369
rect 31021 19329 31033 19363
rect 31067 19329 31079 19363
rect 31021 19323 31079 19329
rect 31113 19363 31171 19369
rect 31113 19329 31125 19363
rect 31159 19329 31171 19363
rect 31113 19323 31171 19329
rect 30892 19320 30898 19323
rect 29730 19292 29736 19304
rect 29420 19264 29500 19292
rect 29643 19264 29736 19292
rect 29420 19252 29426 19264
rect 29730 19252 29736 19264
rect 29788 19292 29794 19304
rect 30742 19292 30748 19304
rect 29788 19264 30748 19292
rect 29788 19252 29794 19264
rect 30742 19252 30748 19264
rect 30800 19252 30806 19304
rect 15120 19196 16712 19224
rect 7837 19159 7895 19165
rect 7837 19156 7849 19159
rect 7524 19128 7849 19156
rect 7524 19116 7530 19128
rect 7837 19125 7849 19128
rect 7883 19125 7895 19159
rect 7837 19119 7895 19125
rect 8021 19159 8079 19165
rect 8021 19125 8033 19159
rect 8067 19125 8079 19159
rect 8846 19156 8852 19168
rect 8807 19128 8852 19156
rect 8021 19119 8079 19125
rect 8846 19116 8852 19128
rect 8904 19116 8910 19168
rect 10965 19159 11023 19165
rect 10965 19125 10977 19159
rect 11011 19156 11023 19159
rect 11238 19156 11244 19168
rect 11011 19128 11244 19156
rect 11011 19125 11023 19128
rect 10965 19119 11023 19125
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 12621 19159 12679 19165
rect 12621 19125 12633 19159
rect 12667 19156 12679 19159
rect 12710 19156 12716 19168
rect 12667 19128 12716 19156
rect 12667 19125 12679 19128
rect 12621 19119 12679 19125
rect 12710 19116 12716 19128
rect 12768 19116 12774 19168
rect 15010 19156 15016 19168
rect 14971 19128 15016 19156
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 15749 19159 15807 19165
rect 15749 19125 15761 19159
rect 15795 19156 15807 19159
rect 15838 19156 15844 19168
rect 15795 19128 15844 19156
rect 15795 19125 15807 19128
rect 15749 19119 15807 19125
rect 15838 19116 15844 19128
rect 15896 19116 15902 19168
rect 16684 19156 16712 19196
rect 17972 19196 24532 19224
rect 17972 19156 18000 19196
rect 26234 19184 26240 19236
rect 26292 19224 26298 19236
rect 27430 19224 27436 19236
rect 26292 19196 27436 19224
rect 26292 19184 26298 19196
rect 27430 19184 27436 19196
rect 27488 19224 27494 19236
rect 27893 19227 27951 19233
rect 27893 19224 27905 19227
rect 27488 19196 27905 19224
rect 27488 19184 27494 19196
rect 27893 19193 27905 19196
rect 27939 19193 27951 19227
rect 27893 19187 27951 19193
rect 29546 19184 29552 19236
rect 29604 19224 29610 19236
rect 31036 19224 31064 19323
rect 29604 19196 31064 19224
rect 31128 19292 31156 19323
rect 31294 19320 31300 19372
rect 31352 19360 31358 19372
rect 32122 19360 32128 19372
rect 31352 19332 31397 19360
rect 31726 19332 32128 19360
rect 31352 19320 31358 19332
rect 31726 19292 31754 19332
rect 32122 19320 32128 19332
rect 32180 19320 32186 19372
rect 33226 19320 33232 19372
rect 33284 19360 33290 19372
rect 33790 19363 33848 19369
rect 33790 19360 33802 19363
rect 33284 19332 33802 19360
rect 33284 19320 33290 19332
rect 33790 19329 33802 19332
rect 33836 19329 33848 19363
rect 33790 19323 33848 19329
rect 34057 19363 34115 19369
rect 34057 19329 34069 19363
rect 34103 19360 34115 19363
rect 34238 19360 34244 19372
rect 34103 19332 34244 19360
rect 34103 19329 34115 19332
rect 34057 19323 34115 19329
rect 34238 19320 34244 19332
rect 34296 19320 34302 19372
rect 35986 19320 35992 19372
rect 36044 19360 36050 19372
rect 36173 19363 36231 19369
rect 36173 19360 36185 19363
rect 36044 19332 36185 19360
rect 36044 19320 36050 19332
rect 36173 19329 36185 19332
rect 36219 19329 36231 19363
rect 36173 19323 36231 19329
rect 36265 19363 36323 19369
rect 36265 19329 36277 19363
rect 36311 19360 36323 19363
rect 36464 19360 36492 19468
rect 39666 19456 39672 19468
rect 39724 19456 39730 19508
rect 41690 19496 41696 19508
rect 41651 19468 41696 19496
rect 41690 19456 41696 19468
rect 41748 19456 41754 19508
rect 36311 19332 36492 19360
rect 36541 19363 36599 19369
rect 36311 19329 36323 19332
rect 36265 19323 36323 19329
rect 36541 19329 36553 19363
rect 36587 19360 36599 19363
rect 37274 19360 37280 19372
rect 36587 19332 37280 19360
rect 36587 19329 36599 19332
rect 36541 19323 36599 19329
rect 37274 19320 37280 19332
rect 37332 19320 37338 19372
rect 37645 19363 37703 19369
rect 37645 19329 37657 19363
rect 37691 19360 37703 19363
rect 38105 19363 38163 19369
rect 38105 19360 38117 19363
rect 37691 19332 38117 19360
rect 37691 19329 37703 19332
rect 37645 19323 37703 19329
rect 38105 19329 38117 19332
rect 38151 19329 38163 19363
rect 38105 19323 38163 19329
rect 31128 19264 31754 19292
rect 29604 19184 29610 19196
rect 16684 19128 18000 19156
rect 18046 19116 18052 19168
rect 18104 19156 18110 19168
rect 21818 19156 21824 19168
rect 18104 19128 18149 19156
rect 21779 19128 21824 19156
rect 18104 19116 18110 19128
rect 21818 19116 21824 19128
rect 21876 19116 21882 19168
rect 25774 19116 25780 19168
rect 25832 19156 25838 19168
rect 27157 19159 27215 19165
rect 27157 19156 27169 19159
rect 25832 19128 27169 19156
rect 25832 19116 25838 19128
rect 27157 19125 27169 19128
rect 27203 19125 27215 19159
rect 30742 19156 30748 19168
rect 30703 19128 30748 19156
rect 27157 19119 27215 19125
rect 30742 19116 30748 19128
rect 30800 19116 30806 19168
rect 30834 19116 30840 19168
rect 30892 19156 30898 19168
rect 31128 19156 31156 19264
rect 36906 19252 36912 19304
rect 36964 19292 36970 19304
rect 37660 19292 37688 19323
rect 40402 19320 40408 19372
rect 40460 19360 40466 19372
rect 40569 19363 40627 19369
rect 40569 19360 40581 19363
rect 40460 19332 40581 19360
rect 40460 19320 40466 19332
rect 40569 19329 40581 19332
rect 40615 19329 40627 19363
rect 40569 19323 40627 19329
rect 36964 19264 37688 19292
rect 39853 19295 39911 19301
rect 36964 19252 36970 19264
rect 39853 19261 39865 19295
rect 39899 19292 39911 19295
rect 39942 19292 39948 19304
rect 39899 19264 39948 19292
rect 39899 19261 39911 19264
rect 39853 19255 39911 19261
rect 39942 19252 39948 19264
rect 40000 19292 40006 19304
rect 40313 19295 40371 19301
rect 40313 19292 40325 19295
rect 40000 19264 40325 19292
rect 40000 19252 40006 19264
rect 40313 19261 40325 19264
rect 40359 19261 40371 19295
rect 40313 19255 40371 19261
rect 30892 19128 31156 19156
rect 30892 19116 30898 19128
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 3237 18955 3295 18961
rect 3237 18921 3249 18955
rect 3283 18952 3295 18955
rect 5258 18952 5264 18964
rect 3283 18924 5264 18952
rect 3283 18921 3295 18924
rect 3237 18915 3295 18921
rect 5258 18912 5264 18924
rect 5316 18912 5322 18964
rect 6273 18955 6331 18961
rect 6273 18921 6285 18955
rect 6319 18952 6331 18955
rect 6638 18952 6644 18964
rect 6319 18924 6644 18952
rect 6319 18921 6331 18924
rect 6273 18915 6331 18921
rect 6638 18912 6644 18924
rect 6696 18952 6702 18964
rect 6696 18924 12112 18952
rect 6696 18912 6702 18924
rect 3786 18844 3792 18896
rect 3844 18884 3850 18896
rect 5629 18887 5687 18893
rect 5629 18884 5641 18887
rect 3844 18856 5641 18884
rect 3844 18844 3850 18856
rect 5629 18853 5641 18856
rect 5675 18884 5687 18887
rect 12084 18884 12112 18924
rect 12158 18912 12164 18964
rect 12216 18952 12222 18964
rect 12897 18955 12955 18961
rect 12897 18952 12909 18955
rect 12216 18924 12909 18952
rect 12216 18912 12222 18924
rect 12897 18921 12909 18924
rect 12943 18921 12955 18955
rect 12897 18915 12955 18921
rect 14366 18912 14372 18964
rect 14424 18952 14430 18964
rect 14461 18955 14519 18961
rect 14461 18952 14473 18955
rect 14424 18924 14473 18952
rect 14424 18912 14430 18924
rect 14461 18921 14473 18924
rect 14507 18921 14519 18955
rect 14461 18915 14519 18921
rect 16301 18955 16359 18961
rect 16301 18921 16313 18955
rect 16347 18952 16359 18955
rect 16758 18952 16764 18964
rect 16347 18924 16764 18952
rect 16347 18921 16359 18924
rect 16301 18915 16359 18921
rect 16758 18912 16764 18924
rect 16816 18912 16822 18964
rect 21683 18955 21741 18961
rect 21683 18952 21695 18955
rect 17972 18924 21695 18952
rect 12710 18884 12716 18896
rect 5675 18856 6914 18884
rect 12084 18856 12716 18884
rect 5675 18853 5687 18856
rect 5629 18847 5687 18853
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 4890 18816 4896 18828
rect 4479 18788 4896 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 1857 18751 1915 18757
rect 1857 18717 1869 18751
rect 1903 18748 1915 18751
rect 2866 18748 2872 18760
rect 1903 18720 2872 18748
rect 1903 18717 1915 18720
rect 1857 18711 1915 18717
rect 2866 18708 2872 18720
rect 2924 18708 2930 18760
rect 4157 18751 4215 18757
rect 4157 18717 4169 18751
rect 4203 18748 4215 18751
rect 4706 18748 4712 18760
rect 4203 18720 4712 18748
rect 4203 18717 4215 18720
rect 4157 18711 4215 18717
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 6886 18748 6914 18856
rect 12710 18844 12716 18856
rect 12768 18884 12774 18896
rect 12768 18856 13768 18884
rect 12768 18844 12774 18856
rect 8205 18819 8263 18825
rect 8205 18785 8217 18819
rect 8251 18816 8263 18819
rect 8294 18816 8300 18828
rect 8251 18788 8300 18816
rect 8251 18785 8263 18788
rect 8205 18779 8263 18785
rect 8294 18776 8300 18788
rect 8352 18816 8358 18828
rect 8662 18816 8668 18828
rect 8352 18788 8668 18816
rect 8352 18776 8358 18788
rect 8662 18776 8668 18788
rect 8720 18816 8726 18828
rect 9582 18816 9588 18828
rect 8720 18788 9588 18816
rect 8720 18776 8726 18788
rect 9582 18776 9588 18788
rect 9640 18816 9646 18828
rect 10229 18819 10287 18825
rect 10229 18816 10241 18819
rect 9640 18788 10241 18816
rect 9640 18776 9646 18788
rect 10229 18785 10241 18788
rect 10275 18785 10287 18819
rect 10229 18779 10287 18785
rect 11238 18748 11244 18760
rect 6886 18720 11244 18748
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 12437 18751 12495 18757
rect 12437 18717 12449 18751
rect 12483 18748 12495 18751
rect 12526 18748 12532 18760
rect 12483 18720 12532 18748
rect 12483 18717 12495 18720
rect 12437 18711 12495 18717
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 2124 18683 2182 18689
rect 2124 18649 2136 18683
rect 2170 18680 2182 18683
rect 2406 18680 2412 18692
rect 2170 18652 2412 18680
rect 2170 18649 2182 18652
rect 2124 18643 2182 18649
rect 2406 18640 2412 18652
rect 2464 18640 2470 18692
rect 5350 18640 5356 18692
rect 5408 18680 5414 18692
rect 5445 18683 5503 18689
rect 5445 18680 5457 18683
rect 5408 18652 5457 18680
rect 5408 18640 5414 18652
rect 5445 18649 5457 18652
rect 5491 18680 5503 18683
rect 5994 18680 6000 18692
rect 5491 18652 6000 18680
rect 5491 18649 5503 18652
rect 5445 18643 5503 18649
rect 5994 18640 6000 18652
rect 6052 18640 6058 18692
rect 6178 18680 6184 18692
rect 6139 18652 6184 18680
rect 6178 18640 6184 18652
rect 6236 18640 6242 18692
rect 6914 18640 6920 18692
rect 6972 18680 6978 18692
rect 7938 18683 7996 18689
rect 7938 18680 7950 18683
rect 6972 18652 7950 18680
rect 6972 18640 6978 18652
rect 7938 18649 7950 18652
rect 7984 18649 7996 18683
rect 7938 18643 7996 18649
rect 10496 18683 10554 18689
rect 10496 18649 10508 18683
rect 10542 18680 10554 18683
rect 11514 18680 11520 18692
rect 10542 18652 11520 18680
rect 10542 18649 10554 18652
rect 10496 18643 10554 18649
rect 11514 18640 11520 18652
rect 11572 18640 11578 18692
rect 12253 18683 12311 18689
rect 12253 18680 12265 18683
rect 11624 18652 12265 18680
rect 11624 18624 11652 18652
rect 12253 18649 12265 18652
rect 12299 18649 12311 18683
rect 13740 18680 13768 18856
rect 17770 18816 17776 18828
rect 16684 18788 17776 18816
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 16684 18757 16712 18788
rect 17770 18776 17776 18788
rect 17828 18816 17834 18828
rect 17972 18816 18000 18924
rect 21683 18921 21695 18924
rect 21729 18921 21741 18955
rect 25774 18952 25780 18964
rect 25735 18924 25780 18952
rect 21683 18915 21741 18921
rect 25774 18912 25780 18924
rect 25832 18912 25838 18964
rect 26142 18912 26148 18964
rect 26200 18952 26206 18964
rect 28350 18952 28356 18964
rect 26200 18924 28356 18952
rect 26200 18912 26206 18924
rect 28350 18912 28356 18924
rect 28408 18912 28414 18964
rect 30101 18955 30159 18961
rect 30101 18921 30113 18955
rect 30147 18952 30159 18955
rect 30745 18955 30803 18961
rect 30745 18952 30757 18955
rect 30147 18924 30757 18952
rect 30147 18921 30159 18924
rect 30101 18915 30159 18921
rect 30745 18921 30757 18924
rect 30791 18921 30803 18955
rect 30745 18915 30803 18921
rect 32953 18955 33011 18961
rect 32953 18921 32965 18955
rect 32999 18952 33011 18955
rect 33226 18952 33232 18964
rect 32999 18924 33232 18952
rect 32999 18921 33011 18924
rect 32953 18915 33011 18921
rect 33226 18912 33232 18924
rect 33284 18912 33290 18964
rect 40402 18952 40408 18964
rect 40363 18924 40408 18952
rect 40402 18912 40408 18924
rect 40460 18912 40466 18964
rect 31294 18884 31300 18896
rect 17828 18788 18000 18816
rect 17828 18776 17834 18788
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 13872 18720 15853 18748
rect 13872 18708 13878 18720
rect 15841 18717 15853 18720
rect 15887 18748 15899 18751
rect 16577 18751 16635 18757
rect 16577 18748 16589 18751
rect 15887 18720 16589 18748
rect 15887 18717 15899 18720
rect 15841 18711 15899 18717
rect 16577 18717 16589 18720
rect 16623 18717 16635 18751
rect 16577 18711 16635 18717
rect 16669 18751 16727 18757
rect 16669 18717 16681 18751
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 16758 18708 16764 18760
rect 16816 18748 16822 18760
rect 16945 18751 17003 18757
rect 16816 18720 16861 18748
rect 16816 18708 16822 18720
rect 16945 18717 16957 18751
rect 16991 18748 17003 18751
rect 17034 18748 17040 18760
rect 16991 18720 17040 18748
rect 16991 18717 17003 18720
rect 16945 18711 17003 18717
rect 17034 18708 17040 18720
rect 17092 18748 17098 18760
rect 17681 18751 17739 18757
rect 17681 18748 17693 18751
rect 17092 18720 17693 18748
rect 17092 18708 17098 18720
rect 17681 18717 17693 18720
rect 17727 18717 17739 18751
rect 17862 18748 17868 18760
rect 17823 18720 17868 18748
rect 17681 18711 17739 18717
rect 17862 18708 17868 18720
rect 17920 18708 17926 18760
rect 17972 18757 18000 18788
rect 20640 18856 31300 18884
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18748 18107 18751
rect 18138 18748 18144 18760
rect 18095 18720 18144 18748
rect 18095 18717 18107 18720
rect 18049 18711 18107 18717
rect 18064 18680 18092 18711
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 19242 18748 19248 18760
rect 19203 18720 19248 18748
rect 19242 18708 19248 18720
rect 19300 18708 19306 18760
rect 13740 18652 18092 18680
rect 18325 18683 18383 18689
rect 12253 18643 12311 18649
rect 18325 18649 18337 18683
rect 18371 18680 18383 18683
rect 19490 18683 19548 18689
rect 19490 18680 19502 18683
rect 18371 18652 19502 18680
rect 18371 18649 18383 18652
rect 18325 18643 18383 18649
rect 19490 18649 19502 18652
rect 19536 18649 19548 18683
rect 19490 18643 19548 18649
rect 3786 18612 3792 18624
rect 3747 18584 3792 18612
rect 3786 18572 3792 18584
rect 3844 18572 3850 18624
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 4522 18612 4528 18624
rect 4295 18584 4528 18612
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 4522 18572 4528 18584
rect 4580 18572 4586 18624
rect 6730 18572 6736 18624
rect 6788 18612 6794 18624
rect 6825 18615 6883 18621
rect 6825 18612 6837 18615
rect 6788 18584 6837 18612
rect 6788 18572 6794 18584
rect 6825 18581 6837 18584
rect 6871 18581 6883 18615
rect 11606 18612 11612 18624
rect 11567 18584 11612 18612
rect 6825 18575 6883 18581
rect 11606 18572 11612 18584
rect 11664 18572 11670 18624
rect 11974 18572 11980 18624
rect 12032 18612 12038 18624
rect 12069 18615 12127 18621
rect 12069 18612 12081 18615
rect 12032 18584 12081 18612
rect 12032 18572 12038 18584
rect 12069 18581 12081 18584
rect 12115 18581 12127 18615
rect 12069 18575 12127 18581
rect 18782 18572 18788 18624
rect 18840 18612 18846 18624
rect 20640 18621 20668 18856
rect 31294 18844 31300 18856
rect 31352 18844 31358 18896
rect 31849 18887 31907 18893
rect 31849 18853 31861 18887
rect 31895 18884 31907 18887
rect 36078 18884 36084 18896
rect 31895 18856 32858 18884
rect 36039 18856 36084 18884
rect 31895 18853 31907 18856
rect 31849 18847 31907 18853
rect 21913 18819 21971 18825
rect 21913 18785 21925 18819
rect 21959 18816 21971 18819
rect 22094 18816 22100 18828
rect 21959 18788 22100 18816
rect 21959 18785 21971 18788
rect 21913 18779 21971 18785
rect 22094 18776 22100 18788
rect 22152 18776 22158 18828
rect 22186 18776 22192 18828
rect 22244 18816 22250 18828
rect 23017 18819 23075 18825
rect 23017 18816 23029 18819
rect 22244 18788 23029 18816
rect 22244 18776 22250 18788
rect 23017 18785 23029 18788
rect 23063 18785 23075 18819
rect 23017 18779 23075 18785
rect 23293 18819 23351 18825
rect 23293 18785 23305 18819
rect 23339 18816 23351 18819
rect 23842 18816 23848 18828
rect 23339 18788 23848 18816
rect 23339 18785 23351 18788
rect 23293 18779 23351 18785
rect 23842 18776 23848 18788
rect 23900 18776 23906 18828
rect 23934 18776 23940 18828
rect 23992 18816 23998 18828
rect 24489 18819 24547 18825
rect 24489 18816 24501 18819
rect 23992 18788 24501 18816
rect 23992 18776 23998 18788
rect 24489 18785 24501 18788
rect 24535 18816 24547 18819
rect 26234 18816 26240 18828
rect 24535 18788 26240 18816
rect 24535 18785 24547 18788
rect 24489 18779 24547 18785
rect 26234 18776 26240 18788
rect 26292 18776 26298 18828
rect 30926 18816 30932 18828
rect 30760 18788 30932 18816
rect 24578 18708 24584 18760
rect 24636 18748 24642 18760
rect 25225 18751 25283 18757
rect 25225 18748 25237 18751
rect 24636 18720 25237 18748
rect 24636 18708 24642 18720
rect 25225 18717 25237 18720
rect 25271 18717 25283 18751
rect 25406 18748 25412 18760
rect 25367 18720 25412 18748
rect 25225 18711 25283 18717
rect 25406 18708 25412 18720
rect 25464 18708 25470 18760
rect 25590 18748 25596 18760
rect 25551 18720 25596 18748
rect 25590 18708 25596 18720
rect 25648 18708 25654 18760
rect 26326 18708 26332 18760
rect 26384 18748 26390 18760
rect 29549 18751 29607 18757
rect 29549 18748 29561 18751
rect 26384 18720 29561 18748
rect 26384 18708 26390 18720
rect 29549 18717 29561 18720
rect 29595 18717 29607 18751
rect 29730 18748 29736 18760
rect 29691 18720 29736 18748
rect 29549 18711 29607 18717
rect 29730 18708 29736 18720
rect 29788 18708 29794 18760
rect 29914 18748 29920 18760
rect 29875 18720 29920 18748
rect 29914 18708 29920 18720
rect 29972 18708 29978 18760
rect 30760 18757 30788 18788
rect 30926 18776 30932 18788
rect 30984 18776 30990 18828
rect 30745 18751 30803 18757
rect 30745 18717 30757 18751
rect 30791 18717 30803 18751
rect 30745 18711 30803 18717
rect 30834 18708 30840 18760
rect 30892 18748 30898 18760
rect 31018 18748 31024 18760
rect 30892 18720 30937 18748
rect 30979 18720 31024 18748
rect 30892 18708 30898 18720
rect 31018 18708 31024 18720
rect 31076 18708 31082 18760
rect 25498 18640 25504 18692
rect 25556 18680 25562 18692
rect 26605 18683 26663 18689
rect 25556 18652 25601 18680
rect 25556 18640 25562 18652
rect 26605 18649 26617 18683
rect 26651 18680 26663 18683
rect 26786 18680 26792 18692
rect 26651 18652 26792 18680
rect 26651 18649 26663 18652
rect 26605 18643 26663 18649
rect 26786 18640 26792 18652
rect 26844 18680 26850 18692
rect 27157 18683 27215 18689
rect 27157 18680 27169 18683
rect 26844 18652 27169 18680
rect 26844 18640 26850 18652
rect 27157 18649 27169 18652
rect 27203 18680 27215 18683
rect 27430 18680 27436 18692
rect 27203 18652 27436 18680
rect 27203 18649 27215 18652
rect 27157 18643 27215 18649
rect 27430 18640 27436 18652
rect 27488 18640 27494 18692
rect 29822 18640 29828 18692
rect 29880 18680 29886 18692
rect 31864 18680 31892 18847
rect 32830 18816 32858 18856
rect 36078 18844 36084 18856
rect 36136 18844 36142 18896
rect 41877 18819 41935 18825
rect 41877 18816 41889 18819
rect 32830 18788 39988 18816
rect 32306 18748 32312 18760
rect 32267 18720 32312 18748
rect 32306 18708 32312 18720
rect 32364 18708 32370 18760
rect 32488 18745 32546 18751
rect 32488 18711 32500 18745
rect 32534 18711 32546 18745
rect 32488 18705 32546 18711
rect 32588 18748 32646 18754
rect 32588 18714 32600 18748
rect 32634 18714 32646 18748
rect 32588 18708 32646 18714
rect 32677 18751 32735 18757
rect 32677 18717 32689 18751
rect 32723 18745 32735 18751
rect 32830 18745 32858 18788
rect 32723 18717 32858 18745
rect 32677 18711 32735 18717
rect 35986 18708 35992 18760
rect 36044 18748 36050 18760
rect 36265 18751 36323 18757
rect 36265 18748 36277 18751
rect 36044 18720 36277 18748
rect 36044 18708 36050 18720
rect 36265 18717 36277 18720
rect 36311 18717 36323 18751
rect 36446 18748 36452 18760
rect 36407 18720 36452 18748
rect 36265 18711 36323 18717
rect 36446 18708 36452 18720
rect 36504 18708 36510 18760
rect 36630 18748 36636 18760
rect 36591 18720 36636 18748
rect 36630 18708 36636 18720
rect 36688 18708 36694 18760
rect 39960 18757 39988 18788
rect 40880 18788 41889 18816
rect 39945 18751 40003 18757
rect 39945 18717 39957 18751
rect 39991 18748 40003 18751
rect 40494 18748 40500 18760
rect 39991 18720 40500 18748
rect 39991 18717 40003 18720
rect 39945 18711 40003 18717
rect 40494 18708 40500 18720
rect 40552 18748 40558 18760
rect 40635 18751 40693 18757
rect 40635 18748 40647 18751
rect 40552 18720 40647 18748
rect 40552 18708 40558 18720
rect 40635 18717 40647 18720
rect 40681 18717 40693 18751
rect 40770 18748 40776 18760
rect 40731 18720 40776 18748
rect 40635 18711 40693 18717
rect 40770 18708 40776 18720
rect 40828 18708 40834 18760
rect 40880 18757 40908 18788
rect 41877 18785 41889 18788
rect 41923 18785 41935 18819
rect 41877 18779 41935 18785
rect 40865 18751 40923 18757
rect 40865 18717 40877 18751
rect 40911 18717 40923 18751
rect 40865 18711 40923 18717
rect 41049 18751 41107 18757
rect 41049 18717 41061 18751
rect 41095 18748 41107 18751
rect 41138 18748 41144 18760
rect 41095 18720 41144 18748
rect 41095 18717 41107 18720
rect 41049 18711 41107 18717
rect 41138 18708 41144 18720
rect 41196 18708 41202 18760
rect 41690 18748 41696 18760
rect 41651 18720 41696 18748
rect 41690 18708 41696 18720
rect 41748 18708 41754 18760
rect 58158 18748 58164 18760
rect 58119 18720 58164 18748
rect 58158 18708 58164 18720
rect 58216 18708 58222 18760
rect 29880 18652 29925 18680
rect 30346 18652 31892 18680
rect 29880 18640 29886 18652
rect 20625 18615 20683 18621
rect 20625 18612 20637 18615
rect 18840 18584 20637 18612
rect 18840 18572 18846 18584
rect 20625 18581 20637 18584
rect 20671 18581 20683 18615
rect 20625 18575 20683 18581
rect 25406 18572 25412 18624
rect 25464 18612 25470 18624
rect 26142 18612 26148 18624
rect 25464 18584 26148 18612
rect 25464 18572 25470 18584
rect 26142 18572 26148 18584
rect 26200 18572 26206 18624
rect 27062 18572 27068 18624
rect 27120 18612 27126 18624
rect 27249 18615 27307 18621
rect 27249 18612 27261 18615
rect 27120 18584 27261 18612
rect 27120 18572 27126 18584
rect 27249 18581 27261 18584
rect 27295 18612 27307 18615
rect 29270 18612 29276 18624
rect 27295 18584 29276 18612
rect 27295 18581 27307 18584
rect 27249 18575 27307 18581
rect 29270 18572 29276 18584
rect 29328 18612 29334 18624
rect 30346 18612 30374 18652
rect 30558 18612 30564 18624
rect 29328 18584 30374 18612
rect 30519 18584 30564 18612
rect 29328 18572 29334 18584
rect 30558 18572 30564 18584
rect 30616 18572 30622 18624
rect 32508 18612 32536 18705
rect 32600 18680 32628 18708
rect 36354 18680 36360 18692
rect 32600 18652 32720 18680
rect 36315 18652 36360 18680
rect 32692 18624 32720 18652
rect 36354 18640 36360 18652
rect 36412 18640 36418 18692
rect 39758 18640 39764 18692
rect 39816 18680 39822 18692
rect 41509 18683 41567 18689
rect 41509 18680 41521 18683
rect 39816 18652 41521 18680
rect 39816 18640 39822 18652
rect 41509 18649 41521 18652
rect 41555 18649 41567 18683
rect 41509 18643 41567 18649
rect 32582 18612 32588 18624
rect 32508 18584 32588 18612
rect 32582 18572 32588 18584
rect 32640 18572 32646 18624
rect 32674 18572 32680 18624
rect 32732 18572 32738 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 2409 18411 2467 18417
rect 2409 18377 2421 18411
rect 2455 18408 2467 18411
rect 2590 18408 2596 18420
rect 2455 18380 2596 18408
rect 2455 18377 2467 18380
rect 2409 18371 2467 18377
rect 2590 18368 2596 18380
rect 2648 18368 2654 18420
rect 4525 18411 4583 18417
rect 4525 18377 4537 18411
rect 4571 18408 4583 18411
rect 4614 18408 4620 18420
rect 4571 18380 4620 18408
rect 4571 18377 4583 18380
rect 4525 18371 4583 18377
rect 4614 18368 4620 18380
rect 4672 18408 4678 18420
rect 9030 18408 9036 18420
rect 4672 18380 9036 18408
rect 4672 18368 4678 18380
rect 9030 18368 9036 18380
rect 9088 18408 9094 18420
rect 9088 18380 9260 18408
rect 9088 18368 9094 18380
rect 3786 18340 3792 18352
rect 3068 18312 3792 18340
rect 3068 18281 3096 18312
rect 3786 18300 3792 18312
rect 3844 18300 3850 18352
rect 6914 18300 6920 18352
rect 6972 18340 6978 18352
rect 8389 18343 8447 18349
rect 6972 18312 7017 18340
rect 6972 18300 6978 18312
rect 8389 18309 8401 18343
rect 8435 18340 8447 18343
rect 8478 18340 8484 18352
rect 8435 18312 8484 18340
rect 8435 18309 8447 18312
rect 8389 18303 8447 18309
rect 8478 18300 8484 18312
rect 8536 18300 8542 18352
rect 9232 18349 9260 18380
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 10505 18411 10563 18417
rect 10505 18408 10517 18411
rect 9640 18380 10517 18408
rect 9640 18368 9646 18380
rect 10505 18377 10517 18380
rect 10551 18408 10563 18411
rect 11054 18408 11060 18420
rect 10551 18380 11060 18408
rect 10551 18377 10563 18380
rect 10505 18371 10563 18377
rect 11054 18368 11060 18380
rect 11112 18368 11118 18420
rect 11514 18408 11520 18420
rect 11475 18380 11520 18408
rect 11514 18368 11520 18380
rect 11572 18368 11578 18420
rect 11698 18368 11704 18420
rect 11756 18408 11762 18420
rect 11756 18380 25452 18408
rect 11756 18368 11762 18380
rect 9217 18343 9275 18349
rect 9217 18309 9229 18343
rect 9263 18309 9275 18343
rect 12066 18340 12072 18352
rect 9217 18303 9275 18309
rect 11900 18312 12072 18340
rect 7665 18285 7723 18291
rect 2225 18275 2283 18281
rect 2225 18241 2237 18275
rect 2271 18272 2283 18275
rect 3053 18275 3111 18281
rect 2271 18244 3004 18272
rect 2271 18241 2283 18244
rect 2225 18235 2283 18241
rect 2041 18207 2099 18213
rect 2041 18173 2053 18207
rect 2087 18204 2099 18207
rect 2869 18207 2927 18213
rect 2869 18204 2881 18207
rect 2087 18176 2881 18204
rect 2087 18173 2099 18176
rect 2041 18167 2099 18173
rect 2240 18148 2268 18176
rect 2869 18173 2881 18176
rect 2915 18173 2927 18207
rect 2976 18204 3004 18244
rect 3053 18241 3065 18275
rect 3099 18241 3111 18275
rect 3053 18235 3111 18241
rect 3237 18275 3295 18281
rect 3237 18241 3249 18275
rect 3283 18272 3295 18275
rect 3881 18275 3939 18281
rect 3881 18272 3893 18275
rect 3283 18244 3893 18272
rect 3283 18241 3295 18244
rect 3237 18235 3295 18241
rect 3881 18241 3893 18244
rect 3927 18241 3939 18275
rect 3881 18235 3939 18241
rect 4985 18275 5043 18281
rect 4985 18241 4997 18275
rect 5031 18272 5043 18275
rect 5902 18272 5908 18284
rect 5031 18244 5908 18272
rect 5031 18241 5043 18244
rect 4985 18235 5043 18241
rect 5902 18232 5908 18244
rect 5960 18232 5966 18284
rect 6730 18232 6736 18284
rect 6788 18272 6794 18284
rect 7101 18275 7159 18281
rect 7101 18272 7113 18275
rect 6788 18244 7113 18272
rect 6788 18232 6794 18244
rect 7101 18241 7113 18244
rect 7147 18241 7159 18275
rect 7101 18235 7159 18241
rect 7190 18232 7196 18284
rect 7248 18281 7254 18284
rect 7248 18275 7297 18281
rect 7248 18241 7251 18275
rect 7285 18241 7297 18275
rect 7248 18235 7297 18241
rect 7248 18232 7254 18235
rect 7475 18232 7481 18284
rect 7533 18270 7539 18284
rect 7533 18242 7576 18270
rect 7665 18251 7677 18285
rect 7711 18272 7723 18285
rect 7711 18251 7788 18272
rect 7665 18245 7788 18251
rect 7668 18244 7788 18245
rect 7533 18232 7539 18242
rect 7760 18216 7788 18244
rect 7926 18232 7932 18284
rect 7984 18272 7990 18284
rect 8205 18275 8263 18281
rect 8205 18272 8217 18275
rect 7984 18244 8217 18272
rect 7984 18232 7990 18244
rect 8205 18241 8217 18244
rect 8251 18241 8263 18275
rect 11514 18272 11520 18284
rect 8205 18235 8263 18241
rect 8312 18244 11520 18272
rect 4798 18204 4804 18216
rect 2976 18176 4804 18204
rect 2869 18167 2927 18173
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 5442 18164 5448 18216
rect 5500 18204 5506 18216
rect 7353 18207 7411 18213
rect 7353 18204 7365 18207
rect 5500 18176 7365 18204
rect 5500 18164 5506 18176
rect 7353 18173 7365 18176
rect 7399 18173 7411 18207
rect 7353 18167 7411 18173
rect 7742 18164 7748 18216
rect 7800 18164 7806 18216
rect 2222 18096 2228 18148
rect 2280 18096 2286 18148
rect 5074 18096 5080 18148
rect 5132 18136 5138 18148
rect 5169 18139 5227 18145
rect 5169 18136 5181 18139
rect 5132 18108 5181 18136
rect 5132 18096 5138 18108
rect 5169 18105 5181 18108
rect 5215 18136 5227 18139
rect 8312 18136 8340 18244
rect 11514 18232 11520 18244
rect 11572 18272 11578 18284
rect 11900 18281 11928 18312
rect 12066 18300 12072 18312
rect 12124 18340 12130 18352
rect 12434 18340 12440 18352
rect 12124 18312 12440 18340
rect 12124 18300 12130 18312
rect 12434 18300 12440 18312
rect 12492 18300 12498 18352
rect 12989 18343 13047 18349
rect 12989 18309 13001 18343
rect 13035 18340 13047 18343
rect 13035 18312 13860 18340
rect 13035 18309 13047 18312
rect 12989 18303 13047 18309
rect 11793 18275 11851 18281
rect 11793 18272 11805 18275
rect 11572 18244 11805 18272
rect 11572 18232 11578 18244
rect 11793 18241 11805 18244
rect 11839 18241 11851 18275
rect 11793 18235 11851 18241
rect 11885 18275 11943 18281
rect 11885 18241 11897 18275
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 11974 18232 11980 18284
rect 12032 18272 12038 18284
rect 12158 18272 12164 18284
rect 12032 18244 12077 18272
rect 12119 18244 12164 18272
rect 12032 18232 12038 18244
rect 12158 18232 12164 18244
rect 12216 18232 12222 18284
rect 8478 18164 8484 18216
rect 8536 18204 8542 18216
rect 13004 18204 13032 18303
rect 13832 18284 13860 18312
rect 16758 18300 16764 18352
rect 16816 18340 16822 18352
rect 17129 18343 17187 18349
rect 17129 18340 17141 18343
rect 16816 18312 17141 18340
rect 16816 18300 16822 18312
rect 17129 18309 17141 18312
rect 17175 18309 17187 18343
rect 17129 18303 17187 18309
rect 17862 18300 17868 18352
rect 17920 18340 17926 18352
rect 18601 18343 18659 18349
rect 18601 18340 18613 18343
rect 17920 18312 18613 18340
rect 17920 18300 17926 18312
rect 18601 18309 18613 18312
rect 18647 18309 18659 18343
rect 18782 18340 18788 18352
rect 18743 18312 18788 18340
rect 18601 18303 18659 18309
rect 18782 18300 18788 18312
rect 18840 18300 18846 18352
rect 19242 18300 19248 18352
rect 19300 18340 19306 18352
rect 23934 18340 23940 18352
rect 19300 18312 22692 18340
rect 23895 18312 23940 18340
rect 19300 18300 19306 18312
rect 13446 18272 13452 18284
rect 13407 18244 13452 18272
rect 13446 18232 13452 18244
rect 13504 18232 13510 18284
rect 13630 18272 13636 18284
rect 13591 18244 13636 18272
rect 13630 18232 13636 18244
rect 13688 18232 13694 18284
rect 13725 18275 13783 18281
rect 13725 18241 13737 18275
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 8536 18176 13032 18204
rect 8536 18164 8542 18176
rect 10962 18136 10968 18148
rect 5215 18108 8340 18136
rect 8404 18108 10968 18136
rect 5215 18105 5227 18108
rect 5169 18099 5227 18105
rect 3694 18068 3700 18080
rect 3655 18040 3700 18068
rect 3694 18028 3700 18040
rect 3752 18028 3758 18080
rect 5350 18028 5356 18080
rect 5408 18068 5414 18080
rect 5721 18071 5779 18077
rect 5721 18068 5733 18071
rect 5408 18040 5733 18068
rect 5408 18028 5414 18040
rect 5721 18037 5733 18040
rect 5767 18037 5779 18071
rect 5721 18031 5779 18037
rect 6178 18028 6184 18080
rect 6236 18068 6242 18080
rect 6365 18071 6423 18077
rect 6365 18068 6377 18071
rect 6236 18040 6377 18068
rect 6236 18028 6242 18040
rect 6365 18037 6377 18040
rect 6411 18068 6423 18071
rect 8404 18068 8432 18108
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 11238 18096 11244 18148
rect 11296 18136 11302 18148
rect 11296 18108 12434 18136
rect 11296 18096 11302 18108
rect 6411 18040 8432 18068
rect 12406 18068 12434 18108
rect 12526 18096 12532 18148
rect 12584 18136 12590 18148
rect 13740 18136 13768 18235
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 17313 18275 17371 18281
rect 13872 18244 13917 18272
rect 13872 18232 13878 18244
rect 17313 18241 17325 18275
rect 17359 18241 17371 18275
rect 17313 18235 17371 18241
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18272 17555 18275
rect 18969 18275 19027 18281
rect 18969 18272 18981 18275
rect 17543 18244 18981 18272
rect 17543 18241 17555 18244
rect 17497 18235 17555 18241
rect 18969 18241 18981 18244
rect 19015 18272 19027 18275
rect 19334 18272 19340 18284
rect 19015 18244 19340 18272
rect 19015 18241 19027 18244
rect 18969 18235 19027 18241
rect 17328 18204 17356 18235
rect 19334 18232 19340 18244
rect 19392 18272 19398 18284
rect 20441 18275 20499 18281
rect 19392 18244 20300 18272
rect 19392 18232 19398 18244
rect 17954 18204 17960 18216
rect 17328 18176 17960 18204
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18204 18107 18207
rect 18138 18204 18144 18216
rect 18095 18176 18144 18204
rect 18095 18173 18107 18176
rect 18049 18167 18107 18173
rect 18138 18164 18144 18176
rect 18196 18164 18202 18216
rect 17862 18136 17868 18148
rect 12584 18108 13768 18136
rect 14016 18108 17868 18136
rect 12584 18096 12590 18108
rect 14016 18068 14044 18108
rect 17862 18096 17868 18108
rect 17920 18096 17926 18148
rect 20272 18145 20300 18244
rect 20441 18241 20453 18275
rect 20487 18272 20499 18275
rect 21085 18275 21143 18281
rect 20487 18244 21036 18272
rect 20487 18241 20499 18244
rect 20441 18235 20499 18241
rect 20901 18207 20959 18213
rect 20901 18204 20913 18207
rect 20456 18176 20913 18204
rect 20257 18139 20315 18145
rect 20257 18105 20269 18139
rect 20303 18105 20315 18139
rect 20257 18099 20315 18105
rect 20456 18080 20484 18176
rect 20901 18173 20913 18176
rect 20947 18173 20959 18207
rect 21008 18204 21036 18244
rect 21085 18241 21097 18275
rect 21131 18272 21143 18275
rect 22370 18272 22376 18284
rect 21131 18244 22376 18272
rect 21131 18241 21143 18244
rect 21085 18235 21143 18241
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 21266 18204 21272 18216
rect 21008 18176 21272 18204
rect 20901 18167 20959 18173
rect 21266 18164 21272 18176
rect 21324 18164 21330 18216
rect 22664 18204 22692 18312
rect 23934 18300 23940 18312
rect 23992 18300 23998 18352
rect 25424 18340 25452 18380
rect 25498 18368 25504 18420
rect 25556 18408 25562 18420
rect 25958 18408 25964 18420
rect 25556 18380 25964 18408
rect 25556 18368 25562 18380
rect 25958 18368 25964 18380
rect 26016 18408 26022 18420
rect 26237 18411 26295 18417
rect 26237 18408 26249 18411
rect 26016 18380 26249 18408
rect 26016 18368 26022 18380
rect 26237 18377 26249 18380
rect 26283 18377 26295 18411
rect 26237 18371 26295 18377
rect 26326 18368 26332 18420
rect 26384 18408 26390 18420
rect 28534 18408 28540 18420
rect 26384 18380 28540 18408
rect 26384 18368 26390 18380
rect 28534 18368 28540 18380
rect 28592 18368 28598 18420
rect 29641 18411 29699 18417
rect 29641 18377 29653 18411
rect 29687 18377 29699 18411
rect 32582 18408 32588 18420
rect 32543 18380 32588 18408
rect 29641 18371 29699 18377
rect 29656 18340 29684 18371
rect 32582 18368 32588 18380
rect 32640 18368 32646 18420
rect 33870 18408 33876 18420
rect 33244 18380 33876 18408
rect 25424 18312 29684 18340
rect 30101 18343 30159 18349
rect 30101 18309 30113 18343
rect 30147 18340 30159 18343
rect 30190 18340 30196 18352
rect 30147 18312 30196 18340
rect 30147 18309 30159 18312
rect 30101 18303 30159 18309
rect 30190 18300 30196 18312
rect 30248 18300 30254 18352
rect 31938 18300 31944 18352
rect 31996 18340 32002 18352
rect 32217 18343 32275 18349
rect 32217 18340 32229 18343
rect 31996 18312 32229 18340
rect 31996 18300 32002 18312
rect 32217 18309 32229 18312
rect 32263 18309 32275 18343
rect 32398 18340 32404 18352
rect 32359 18312 32404 18340
rect 32217 18303 32275 18309
rect 25124 18275 25182 18281
rect 25124 18241 25136 18275
rect 25170 18272 25182 18275
rect 25682 18272 25688 18284
rect 25170 18244 25688 18272
rect 25170 18241 25182 18244
rect 25124 18235 25182 18241
rect 25682 18232 25688 18244
rect 25740 18232 25746 18284
rect 29825 18275 29883 18281
rect 29825 18241 29837 18275
rect 29871 18272 29883 18275
rect 32232 18272 32260 18303
rect 32398 18300 32404 18312
rect 32456 18300 32462 18352
rect 33244 18349 33272 18380
rect 33870 18368 33876 18380
rect 33928 18368 33934 18420
rect 38746 18408 38752 18420
rect 38707 18380 38752 18408
rect 38746 18368 38752 18380
rect 38804 18368 38810 18420
rect 33229 18343 33287 18349
rect 33229 18309 33241 18343
rect 33275 18309 33287 18343
rect 33229 18303 33287 18309
rect 34057 18343 34115 18349
rect 34057 18309 34069 18343
rect 34103 18340 34115 18343
rect 34146 18340 34152 18352
rect 34103 18312 34152 18340
rect 34103 18309 34115 18312
rect 34057 18303 34115 18309
rect 34146 18300 34152 18312
rect 34204 18300 34210 18352
rect 39884 18343 39942 18349
rect 39884 18309 39896 18343
rect 39930 18340 39942 18343
rect 40589 18343 40647 18349
rect 40589 18340 40601 18343
rect 39930 18312 40601 18340
rect 39930 18309 39942 18312
rect 39884 18303 39942 18309
rect 40589 18309 40601 18312
rect 40635 18309 40647 18343
rect 40589 18303 40647 18309
rect 33413 18275 33471 18281
rect 33413 18272 33425 18275
rect 29871 18244 30052 18272
rect 32232 18244 33425 18272
rect 29871 18241 29883 18244
rect 29825 18235 29883 18241
rect 23198 18204 23204 18216
rect 22664 18176 23204 18204
rect 22664 18145 22692 18176
rect 23198 18164 23204 18176
rect 23256 18204 23262 18216
rect 24857 18207 24915 18213
rect 24857 18204 24869 18207
rect 23256 18176 24869 18204
rect 23256 18164 23262 18176
rect 24857 18173 24869 18176
rect 24903 18173 24915 18207
rect 24857 18167 24915 18173
rect 28534 18164 28540 18216
rect 28592 18204 28598 18216
rect 29917 18207 29975 18213
rect 29917 18204 29929 18207
rect 28592 18176 29929 18204
rect 28592 18164 28598 18176
rect 29917 18173 29929 18176
rect 29963 18173 29975 18207
rect 30024 18204 30052 18244
rect 33413 18241 33425 18244
rect 33459 18272 33471 18275
rect 33873 18275 33931 18281
rect 33873 18272 33885 18275
rect 33459 18244 33885 18272
rect 33459 18241 33471 18244
rect 33413 18235 33471 18241
rect 33873 18241 33885 18244
rect 33919 18241 33931 18275
rect 33873 18235 33931 18241
rect 37553 18275 37611 18281
rect 37553 18241 37565 18275
rect 37599 18272 37611 18275
rect 38470 18272 38476 18284
rect 37599 18244 38476 18272
rect 37599 18241 37611 18244
rect 37553 18235 37611 18241
rect 38470 18232 38476 18244
rect 38528 18232 38534 18284
rect 38930 18232 38936 18284
rect 38988 18272 38994 18284
rect 38988 18244 40448 18272
rect 38988 18232 38994 18244
rect 33778 18204 33784 18216
rect 30024 18176 33784 18204
rect 29917 18167 29975 18173
rect 33778 18164 33784 18176
rect 33836 18164 33842 18216
rect 37277 18207 37335 18213
rect 37277 18173 37289 18207
rect 37323 18204 37335 18207
rect 37642 18204 37648 18216
rect 37323 18176 37648 18204
rect 37323 18173 37335 18176
rect 37277 18167 37335 18173
rect 37642 18164 37648 18176
rect 37700 18164 37706 18216
rect 40129 18207 40187 18213
rect 40129 18173 40141 18207
rect 40175 18173 40187 18207
rect 40420 18204 40448 18244
rect 40494 18232 40500 18284
rect 40552 18272 40558 18284
rect 40819 18275 40877 18281
rect 40819 18272 40831 18275
rect 40552 18244 40831 18272
rect 40552 18232 40558 18244
rect 40819 18241 40831 18244
rect 40865 18241 40877 18275
rect 40954 18272 40960 18284
rect 40915 18244 40960 18272
rect 40819 18235 40877 18241
rect 40954 18232 40960 18244
rect 41012 18232 41018 18284
rect 41046 18232 41052 18284
rect 41104 18272 41110 18284
rect 41233 18275 41291 18281
rect 41104 18244 41149 18272
rect 41104 18232 41110 18244
rect 41233 18241 41245 18275
rect 41279 18272 41291 18275
rect 41693 18275 41751 18281
rect 41693 18272 41705 18275
rect 41279 18244 41705 18272
rect 41279 18241 41291 18244
rect 41233 18235 41291 18241
rect 41693 18241 41705 18244
rect 41739 18241 41751 18275
rect 41693 18235 41751 18241
rect 41248 18204 41276 18235
rect 40420 18176 41276 18204
rect 40129 18167 40187 18173
rect 22649 18139 22707 18145
rect 22649 18105 22661 18139
rect 22695 18105 22707 18139
rect 22649 18099 22707 18105
rect 32950 18096 32956 18148
rect 33008 18136 33014 18148
rect 34241 18139 34299 18145
rect 34241 18136 34253 18139
rect 33008 18108 34253 18136
rect 33008 18096 33014 18108
rect 34241 18105 34253 18108
rect 34287 18105 34299 18139
rect 34241 18099 34299 18105
rect 12406 18040 14044 18068
rect 14093 18071 14151 18077
rect 6411 18037 6423 18040
rect 6365 18031 6423 18037
rect 14093 18037 14105 18071
rect 14139 18068 14151 18071
rect 15194 18068 15200 18080
rect 14139 18040 15200 18068
rect 14139 18037 14151 18040
rect 14093 18031 14151 18037
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 15838 18028 15844 18080
rect 15896 18068 15902 18080
rect 19797 18071 19855 18077
rect 19797 18068 19809 18071
rect 15896 18040 19809 18068
rect 15896 18028 15902 18040
rect 19797 18037 19809 18040
rect 19843 18068 19855 18071
rect 20438 18068 20444 18080
rect 19843 18040 20444 18068
rect 19843 18037 19855 18040
rect 19797 18031 19855 18037
rect 20438 18028 20444 18040
rect 20496 18028 20502 18080
rect 20898 18028 20904 18080
rect 20956 18068 20962 18080
rect 24670 18068 24676 18080
rect 20956 18040 24676 18068
rect 20956 18028 20962 18040
rect 24670 18028 24676 18040
rect 24728 18028 24734 18080
rect 30101 18071 30159 18077
rect 30101 18037 30113 18071
rect 30147 18068 30159 18071
rect 30742 18068 30748 18080
rect 30147 18040 30748 18068
rect 30147 18037 30159 18040
rect 30101 18031 30159 18037
rect 30742 18028 30748 18040
rect 30800 18028 30806 18080
rect 33042 18068 33048 18080
rect 33003 18040 33048 18068
rect 33042 18028 33048 18040
rect 33100 18028 33106 18080
rect 35618 18028 35624 18080
rect 35676 18068 35682 18080
rect 36357 18071 36415 18077
rect 36357 18068 36369 18071
rect 35676 18040 36369 18068
rect 35676 18028 35682 18040
rect 36357 18037 36369 18040
rect 36403 18068 36415 18071
rect 38930 18068 38936 18080
rect 36403 18040 38936 18068
rect 36403 18037 36415 18040
rect 36357 18031 36415 18037
rect 38930 18028 38936 18040
rect 38988 18028 38994 18080
rect 39942 18028 39948 18080
rect 40000 18068 40006 18080
rect 40144 18068 40172 18167
rect 40880 18148 40908 18176
rect 40862 18096 40868 18148
rect 40920 18096 40926 18148
rect 40000 18040 40172 18068
rect 40000 18028 40006 18040
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4120 17836 5396 17864
rect 4120 17824 4126 17836
rect 4341 17799 4399 17805
rect 4341 17765 4353 17799
rect 4387 17796 4399 17799
rect 4706 17796 4712 17808
rect 4387 17768 4712 17796
rect 4387 17765 4399 17768
rect 4341 17759 4399 17765
rect 4706 17756 4712 17768
rect 4764 17796 4770 17808
rect 4982 17796 4988 17808
rect 4764 17768 4988 17796
rect 4764 17756 4770 17768
rect 4982 17756 4988 17768
rect 5040 17756 5046 17808
rect 5258 17796 5264 17808
rect 5184 17768 5264 17796
rect 5184 17737 5212 17768
rect 5258 17756 5264 17768
rect 5316 17756 5322 17808
rect 5368 17796 5396 17836
rect 5442 17824 5448 17876
rect 5500 17864 5506 17876
rect 9030 17864 9036 17876
rect 5500 17836 5545 17864
rect 8991 17836 9036 17864
rect 5500 17824 5506 17836
rect 9030 17824 9036 17836
rect 9088 17824 9094 17876
rect 9398 17824 9404 17876
rect 9456 17864 9462 17876
rect 10781 17867 10839 17873
rect 10781 17864 10793 17867
rect 9456 17836 10793 17864
rect 9456 17824 9462 17836
rect 10781 17833 10793 17836
rect 10827 17833 10839 17867
rect 10781 17827 10839 17833
rect 5368 17768 6914 17796
rect 5169 17731 5227 17737
rect 5169 17697 5181 17731
rect 5215 17697 5227 17731
rect 6886 17728 6914 17768
rect 6886 17700 8294 17728
rect 5169 17691 5227 17697
rect 5261 17663 5319 17669
rect 5261 17629 5273 17663
rect 5307 17660 5319 17663
rect 5626 17660 5632 17672
rect 5307 17632 5632 17660
rect 5307 17629 5319 17632
rect 5261 17623 5319 17629
rect 5626 17620 5632 17632
rect 5684 17620 5690 17672
rect 8266 17592 8294 17700
rect 10796 17660 10824 17827
rect 10870 17824 10876 17876
rect 10928 17864 10934 17876
rect 11146 17864 11152 17876
rect 10928 17836 11152 17864
rect 10928 17824 10934 17836
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 13541 17867 13599 17873
rect 13541 17833 13553 17867
rect 13587 17864 13599 17867
rect 13630 17864 13636 17876
rect 13587 17836 13636 17864
rect 13587 17833 13599 17836
rect 13541 17827 13599 17833
rect 13630 17824 13636 17836
rect 13688 17824 13694 17876
rect 21821 17867 21879 17873
rect 21821 17833 21833 17867
rect 21867 17864 21879 17867
rect 21910 17864 21916 17876
rect 21867 17836 21916 17864
rect 21867 17833 21879 17836
rect 21821 17827 21879 17833
rect 21910 17824 21916 17836
rect 21968 17824 21974 17876
rect 25682 17864 25688 17876
rect 25643 17836 25688 17864
rect 25682 17824 25688 17836
rect 25740 17824 25746 17876
rect 30745 17867 30803 17873
rect 30745 17833 30757 17867
rect 30791 17864 30803 17867
rect 31938 17864 31944 17876
rect 30791 17836 31944 17864
rect 30791 17833 30803 17836
rect 30745 17827 30803 17833
rect 31938 17824 31944 17836
rect 31996 17824 32002 17876
rect 36722 17864 36728 17876
rect 32600 17836 36584 17864
rect 36683 17836 36728 17864
rect 24949 17799 25007 17805
rect 24949 17765 24961 17799
rect 24995 17796 25007 17799
rect 25130 17796 25136 17808
rect 24995 17768 25136 17796
rect 24995 17765 25007 17768
rect 24949 17759 25007 17765
rect 25130 17756 25136 17768
rect 25188 17756 25194 17808
rect 26970 17756 26976 17808
rect 27028 17796 27034 17808
rect 32600 17796 32628 17836
rect 27028 17768 32628 17796
rect 27028 17756 27034 17768
rect 34606 17756 34612 17808
rect 34664 17796 34670 17808
rect 35802 17796 35808 17808
rect 34664 17768 35808 17796
rect 34664 17756 34670 17768
rect 35802 17756 35808 17768
rect 35860 17756 35866 17808
rect 36556 17796 36584 17836
rect 36722 17824 36728 17836
rect 36780 17824 36786 17876
rect 40405 17867 40463 17873
rect 40405 17833 40417 17867
rect 40451 17864 40463 17867
rect 41046 17864 41052 17876
rect 40451 17836 41052 17864
rect 40451 17833 40463 17836
rect 40405 17827 40463 17833
rect 41046 17824 41052 17836
rect 41104 17824 41110 17876
rect 37366 17796 37372 17808
rect 36556 17768 37372 17796
rect 37366 17756 37372 17768
rect 37424 17756 37430 17808
rect 38013 17799 38071 17805
rect 38013 17765 38025 17799
rect 38059 17796 38071 17799
rect 40954 17796 40960 17808
rect 38059 17768 40960 17796
rect 38059 17765 38071 17768
rect 38013 17759 38071 17765
rect 40954 17756 40960 17768
rect 41012 17756 41018 17808
rect 15473 17731 15531 17737
rect 15473 17697 15485 17731
rect 15519 17728 15531 17731
rect 16482 17728 16488 17740
rect 15519 17700 16488 17728
rect 15519 17697 15531 17700
rect 15473 17691 15531 17697
rect 16482 17688 16488 17700
rect 16540 17688 16546 17740
rect 20898 17688 20904 17740
rect 20956 17728 20962 17740
rect 21818 17728 21824 17740
rect 20956 17700 21128 17728
rect 20956 17688 20962 17700
rect 12158 17660 12164 17672
rect 10796 17632 12164 17660
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17629 12311 17663
rect 12253 17623 12311 17629
rect 8266 17564 12020 17592
rect 4706 17484 4712 17536
rect 4764 17524 4770 17536
rect 4801 17527 4859 17533
rect 4801 17524 4813 17527
rect 4764 17496 4813 17524
rect 4764 17484 4770 17496
rect 4801 17493 4813 17496
rect 4847 17493 4859 17527
rect 5902 17524 5908 17536
rect 5863 17496 5908 17524
rect 4801 17487 4859 17493
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 7926 17524 7932 17536
rect 7887 17496 7932 17524
rect 7926 17484 7932 17496
rect 7984 17484 7990 17536
rect 11425 17527 11483 17533
rect 11425 17493 11437 17527
rect 11471 17524 11483 17527
rect 11514 17524 11520 17536
rect 11471 17496 11520 17524
rect 11471 17493 11483 17496
rect 11425 17487 11483 17493
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 11882 17524 11888 17536
rect 11843 17496 11888 17524
rect 11882 17484 11888 17496
rect 11940 17484 11946 17536
rect 11992 17524 12020 17564
rect 12066 17552 12072 17604
rect 12124 17592 12130 17604
rect 12268 17592 12296 17623
rect 12342 17620 12348 17672
rect 12400 17660 12406 17672
rect 12529 17663 12587 17669
rect 12400 17632 12445 17660
rect 12400 17620 12406 17632
rect 12529 17629 12541 17663
rect 12575 17629 12587 17663
rect 12529 17623 12587 17629
rect 12124 17564 12296 17592
rect 12544 17592 12572 17623
rect 12618 17620 12624 17672
rect 12676 17660 12682 17672
rect 13173 17663 13231 17669
rect 13173 17660 13185 17663
rect 12676 17632 13185 17660
rect 12676 17620 12682 17632
rect 13173 17629 13185 17632
rect 13219 17629 13231 17663
rect 13446 17660 13452 17672
rect 13173 17623 13231 17629
rect 13280 17632 13452 17660
rect 13280 17592 13308 17632
rect 13446 17620 13452 17632
rect 13504 17620 13510 17672
rect 15194 17620 15200 17672
rect 15252 17669 15258 17672
rect 21100 17669 21128 17700
rect 21284 17700 21824 17728
rect 15252 17660 15264 17669
rect 20993 17663 21051 17669
rect 15252 17632 15297 17660
rect 15252 17623 15264 17632
rect 20993 17629 21005 17663
rect 21039 17629 21051 17663
rect 20993 17623 21051 17629
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 21198 17663 21256 17669
rect 21198 17629 21210 17663
rect 21244 17660 21256 17663
rect 21284 17660 21312 17700
rect 21818 17688 21824 17700
rect 21876 17688 21882 17740
rect 23198 17728 23204 17740
rect 23159 17700 23204 17728
rect 23198 17688 23204 17700
rect 23256 17688 23262 17740
rect 25406 17728 25412 17740
rect 24596 17700 25412 17728
rect 21244 17632 21312 17660
rect 21244 17629 21256 17632
rect 21198 17623 21256 17629
rect 15252 17620 15258 17623
rect 12544 17564 13308 17592
rect 13357 17595 13415 17601
rect 12124 17552 12130 17564
rect 13357 17561 13369 17595
rect 13403 17592 13415 17595
rect 20717 17595 20775 17601
rect 13403 17564 14136 17592
rect 13403 17561 13415 17564
rect 13357 17555 13415 17561
rect 13078 17524 13084 17536
rect 11992 17496 13084 17524
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 14108 17533 14136 17564
rect 20717 17561 20729 17595
rect 20763 17592 20775 17595
rect 20806 17592 20812 17604
rect 20763 17564 20812 17592
rect 20763 17561 20775 17564
rect 20717 17555 20775 17561
rect 20806 17552 20812 17564
rect 20864 17552 20870 17604
rect 14093 17527 14151 17533
rect 14093 17493 14105 17527
rect 14139 17524 14151 17527
rect 14274 17524 14280 17536
rect 14139 17496 14280 17524
rect 14139 17493 14151 17496
rect 14093 17487 14151 17493
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 20257 17527 20315 17533
rect 20257 17493 20269 17527
rect 20303 17524 20315 17527
rect 21008 17524 21036 17623
rect 21358 17620 21364 17672
rect 21416 17660 21422 17672
rect 21416 17632 21461 17660
rect 21416 17620 21422 17632
rect 22922 17620 22928 17672
rect 22980 17669 22986 17672
rect 22980 17660 22992 17669
rect 24394 17660 24400 17672
rect 22980 17632 23025 17660
rect 24355 17632 24400 17660
rect 22980 17623 22992 17632
rect 22980 17620 22986 17623
rect 24394 17620 24400 17632
rect 24452 17620 24458 17672
rect 23290 17552 23296 17604
rect 23348 17592 23354 17604
rect 24596 17601 24624 17700
rect 25406 17688 25412 17700
rect 25464 17688 25470 17740
rect 33042 17728 33048 17740
rect 32692 17700 33048 17728
rect 24762 17660 24768 17672
rect 24723 17632 24768 17660
rect 24762 17620 24768 17632
rect 24820 17660 24826 17672
rect 25590 17660 25596 17672
rect 24820 17632 25596 17660
rect 24820 17620 24826 17632
rect 25590 17620 25596 17632
rect 25648 17620 25654 17672
rect 25961 17663 26019 17669
rect 25961 17629 25973 17663
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 26053 17663 26111 17669
rect 26053 17629 26065 17663
rect 26099 17629 26111 17663
rect 26053 17623 26111 17629
rect 24581 17595 24639 17601
rect 24581 17592 24593 17595
rect 23348 17564 24593 17592
rect 23348 17552 23354 17564
rect 24581 17561 24593 17564
rect 24627 17561 24639 17595
rect 24581 17555 24639 17561
rect 24673 17595 24731 17601
rect 24673 17561 24685 17595
rect 24719 17592 24731 17595
rect 25866 17592 25872 17604
rect 24719 17564 25872 17592
rect 24719 17561 24731 17564
rect 24673 17555 24731 17561
rect 25866 17552 25872 17564
rect 25924 17552 25930 17604
rect 21082 17524 21088 17536
rect 20303 17496 21088 17524
rect 20303 17493 20315 17496
rect 20257 17487 20315 17493
rect 21082 17484 21088 17496
rect 21140 17524 21146 17536
rect 25976 17524 26004 17623
rect 26068 17592 26096 17623
rect 26142 17620 26148 17672
rect 26200 17660 26206 17672
rect 26329 17663 26387 17669
rect 26200 17632 26245 17660
rect 26200 17620 26206 17632
rect 26329 17629 26341 17663
rect 26375 17660 26387 17663
rect 26602 17660 26608 17672
rect 26375 17632 26608 17660
rect 26375 17629 26387 17632
rect 26329 17623 26387 17629
rect 26602 17620 26608 17632
rect 26660 17660 26666 17672
rect 28350 17660 28356 17672
rect 26660 17632 28356 17660
rect 26660 17620 26666 17632
rect 28350 17620 28356 17632
rect 28408 17620 28414 17672
rect 30561 17663 30619 17669
rect 30561 17629 30573 17663
rect 30607 17660 30619 17663
rect 31386 17660 31392 17672
rect 30607 17632 31392 17660
rect 30607 17629 30619 17632
rect 30561 17623 30619 17629
rect 31386 17620 31392 17632
rect 31444 17620 31450 17672
rect 32490 17660 32496 17672
rect 32451 17632 32496 17660
rect 32490 17620 32496 17632
rect 32548 17620 32554 17672
rect 32692 17669 32720 17700
rect 33042 17688 33048 17700
rect 33100 17688 33106 17740
rect 40494 17688 40500 17740
rect 40552 17728 40558 17740
rect 40865 17731 40923 17737
rect 40865 17728 40877 17731
rect 40552 17700 40877 17728
rect 40552 17688 40558 17700
rect 40865 17697 40877 17700
rect 40911 17697 40923 17731
rect 40865 17691 40923 17697
rect 32672 17663 32730 17669
rect 32672 17629 32684 17663
rect 32718 17629 32730 17663
rect 32769 17663 32827 17669
rect 32769 17648 32781 17663
rect 32815 17648 32827 17663
rect 32881 17663 32939 17669
rect 32672 17623 32730 17629
rect 27062 17592 27068 17604
rect 26068 17564 27068 17592
rect 27062 17552 27068 17564
rect 27120 17552 27126 17604
rect 28258 17552 28264 17604
rect 28316 17592 28322 17604
rect 32582 17592 32588 17604
rect 28316 17564 32588 17592
rect 28316 17552 28322 17564
rect 32582 17552 32588 17564
rect 32640 17552 32646 17604
rect 32766 17596 32772 17648
rect 32824 17596 32830 17648
rect 32881 17629 32893 17663
rect 32927 17660 32939 17663
rect 35618 17660 35624 17672
rect 32927 17632 32996 17660
rect 35579 17632 35624 17660
rect 32927 17629 32939 17632
rect 32881 17623 32939 17629
rect 26878 17524 26884 17536
rect 21140 17496 26884 17524
rect 21140 17484 21146 17496
rect 26878 17484 26884 17496
rect 26936 17484 26942 17536
rect 31938 17524 31944 17536
rect 31899 17496 31944 17524
rect 31938 17484 31944 17496
rect 31996 17524 32002 17536
rect 32968 17524 32996 17632
rect 35618 17620 35624 17632
rect 35676 17620 35682 17672
rect 35802 17660 35808 17672
rect 35763 17632 35808 17660
rect 35802 17620 35808 17632
rect 35860 17620 35866 17672
rect 35897 17663 35955 17669
rect 35897 17629 35909 17663
rect 35943 17629 35955 17663
rect 35897 17623 35955 17629
rect 35912 17592 35940 17623
rect 35986 17620 35992 17672
rect 36044 17660 36050 17672
rect 36909 17663 36967 17669
rect 36044 17632 36089 17660
rect 36044 17620 36050 17632
rect 36909 17629 36921 17663
rect 36955 17660 36967 17663
rect 37182 17660 37188 17672
rect 36955 17632 37188 17660
rect 36955 17629 36967 17632
rect 36909 17623 36967 17629
rect 37182 17620 37188 17632
rect 37240 17620 37246 17672
rect 37277 17663 37335 17669
rect 37277 17629 37289 17663
rect 37323 17660 37335 17663
rect 37458 17660 37464 17672
rect 37323 17632 37464 17660
rect 37323 17629 37335 17632
rect 37277 17623 37335 17629
rect 37458 17620 37464 17632
rect 37516 17620 37522 17672
rect 38746 17620 38752 17672
rect 38804 17660 38810 17672
rect 40221 17663 40279 17669
rect 40221 17660 40233 17663
rect 38804 17632 40233 17660
rect 38804 17620 38810 17632
rect 40221 17629 40233 17632
rect 40267 17629 40279 17663
rect 40221 17623 40279 17629
rect 35912 17564 36492 17592
rect 33134 17524 33140 17536
rect 31996 17496 32996 17524
rect 33095 17496 33140 17524
rect 31996 17484 32002 17496
rect 33134 17484 33140 17496
rect 33192 17484 33198 17536
rect 35066 17524 35072 17536
rect 35027 17496 35072 17524
rect 35066 17484 35072 17496
rect 35124 17524 35130 17536
rect 35526 17524 35532 17536
rect 35124 17496 35532 17524
rect 35124 17484 35130 17496
rect 35526 17484 35532 17496
rect 35584 17524 35590 17536
rect 35986 17524 35992 17536
rect 35584 17496 35992 17524
rect 35584 17484 35590 17496
rect 35986 17484 35992 17496
rect 36044 17484 36050 17536
rect 36262 17524 36268 17536
rect 36223 17496 36268 17524
rect 36262 17484 36268 17496
rect 36320 17484 36326 17536
rect 36464 17524 36492 17564
rect 36538 17552 36544 17604
rect 36596 17592 36602 17604
rect 37001 17595 37059 17601
rect 37001 17592 37013 17595
rect 36596 17564 37013 17592
rect 36596 17552 36602 17564
rect 37001 17561 37013 17564
rect 37047 17561 37059 17595
rect 37001 17555 37059 17561
rect 37090 17552 37096 17604
rect 37148 17592 37154 17604
rect 37826 17592 37832 17604
rect 37148 17564 37193 17592
rect 37787 17564 37832 17592
rect 37148 17552 37154 17564
rect 37826 17552 37832 17564
rect 37884 17552 37890 17604
rect 38470 17552 38476 17604
rect 38528 17592 38534 17604
rect 40037 17595 40095 17601
rect 40037 17592 40049 17595
rect 38528 17564 40049 17592
rect 38528 17552 38534 17564
rect 40037 17561 40049 17564
rect 40083 17561 40095 17595
rect 40037 17555 40095 17561
rect 37844 17524 37872 17552
rect 36464 17496 37872 17524
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 4157 17323 4215 17329
rect 4157 17289 4169 17323
rect 4203 17320 4215 17323
rect 4614 17320 4620 17332
rect 4203 17292 4620 17320
rect 4203 17289 4215 17292
rect 4157 17283 4215 17289
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 12253 17323 12311 17329
rect 12253 17289 12265 17323
rect 12299 17320 12311 17323
rect 12342 17320 12348 17332
rect 12299 17292 12348 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 13817 17323 13875 17329
rect 13817 17289 13829 17323
rect 13863 17320 13875 17323
rect 13906 17320 13912 17332
rect 13863 17292 13912 17320
rect 13863 17289 13875 17292
rect 13817 17283 13875 17289
rect 13906 17280 13912 17292
rect 13964 17280 13970 17332
rect 19705 17323 19763 17329
rect 19705 17320 19717 17323
rect 14016 17292 19717 17320
rect 3044 17255 3102 17261
rect 3044 17221 3056 17255
rect 3090 17252 3102 17255
rect 3694 17252 3700 17264
rect 3090 17224 3700 17252
rect 3090 17221 3102 17224
rect 3044 17215 3102 17221
rect 3694 17212 3700 17224
rect 3752 17212 3758 17264
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17184 2835 17187
rect 2866 17184 2872 17196
rect 2823 17156 2872 17184
rect 2823 17153 2835 17156
rect 2777 17147 2835 17153
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 4632 17184 4660 17280
rect 11885 17255 11943 17261
rect 11885 17221 11897 17255
rect 11931 17252 11943 17255
rect 12618 17252 12624 17264
rect 11931 17224 12624 17252
rect 11931 17221 11943 17224
rect 11885 17215 11943 17221
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 13078 17212 13084 17264
rect 13136 17252 13142 17264
rect 14016 17252 14044 17292
rect 19705 17289 19717 17292
rect 19751 17289 19763 17323
rect 25682 17320 25688 17332
rect 19705 17283 19763 17289
rect 24872 17292 25688 17320
rect 14182 17252 14188 17264
rect 13136 17224 14044 17252
rect 14143 17224 14188 17252
rect 13136 17212 13142 17224
rect 14182 17212 14188 17224
rect 14240 17252 14246 17264
rect 14550 17252 14556 17264
rect 14240 17224 14556 17252
rect 14240 17212 14246 17224
rect 14550 17212 14556 17224
rect 14608 17212 14614 17264
rect 17034 17252 17040 17264
rect 15120 17224 17040 17252
rect 5077 17187 5135 17193
rect 5077 17184 5089 17187
rect 4632 17156 5089 17184
rect 5077 17153 5089 17156
rect 5123 17153 5135 17187
rect 5077 17147 5135 17153
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 8398 17187 8456 17193
rect 8398 17184 8410 17187
rect 8076 17156 8410 17184
rect 8076 17144 8082 17156
rect 8398 17153 8410 17156
rect 8444 17153 8456 17187
rect 8662 17184 8668 17196
rect 8623 17156 8668 17184
rect 8398 17147 8456 17153
rect 8662 17144 8668 17156
rect 8720 17184 8726 17196
rect 9122 17184 9128 17196
rect 8720 17156 9128 17184
rect 8720 17144 8726 17156
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 12069 17187 12127 17193
rect 12069 17153 12081 17187
rect 12115 17184 12127 17187
rect 12434 17184 12440 17196
rect 12115 17156 12440 17184
rect 12115 17153 12127 17156
rect 12069 17147 12127 17153
rect 12434 17144 12440 17156
rect 12492 17144 12498 17196
rect 13814 17144 13820 17196
rect 13872 17184 13878 17196
rect 13955 17187 14013 17193
rect 13955 17184 13967 17187
rect 13872 17156 13967 17184
rect 13872 17144 13878 17156
rect 13955 17153 13967 17156
rect 14001 17153 14013 17187
rect 13955 17147 14013 17153
rect 14093 17187 14151 17193
rect 14093 17153 14105 17187
rect 14139 17153 14151 17187
rect 14093 17147 14151 17153
rect 4706 17116 4712 17128
rect 4667 17088 4712 17116
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 5169 17119 5227 17125
rect 5169 17085 5181 17119
rect 5215 17116 5227 17119
rect 5626 17116 5632 17128
rect 5215 17088 5632 17116
rect 5215 17085 5227 17088
rect 5169 17079 5227 17085
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 14108 17116 14136 17147
rect 14274 17144 14280 17196
rect 14332 17193 14338 17196
rect 14332 17187 14371 17193
rect 14359 17153 14371 17187
rect 14458 17184 14464 17196
rect 14419 17156 14464 17184
rect 14332 17147 14371 17153
rect 14332 17144 14338 17147
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 15120 17184 15148 17224
rect 17034 17212 17040 17224
rect 17092 17212 17098 17264
rect 17954 17252 17960 17264
rect 17915 17224 17960 17252
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 24872 17252 24900 17292
rect 25682 17280 25688 17292
rect 25740 17280 25746 17332
rect 25869 17323 25927 17329
rect 25869 17289 25881 17323
rect 25915 17320 25927 17323
rect 26142 17320 26148 17332
rect 25915 17292 26148 17320
rect 25915 17289 25927 17292
rect 25869 17283 25927 17289
rect 26142 17280 26148 17292
rect 26200 17280 26206 17332
rect 26878 17280 26884 17332
rect 26936 17320 26942 17332
rect 26936 17292 31754 17320
rect 26936 17280 26942 17292
rect 18156 17224 24900 17252
rect 14568 17156 15148 17184
rect 15197 17187 15255 17193
rect 14568 17116 14596 17156
rect 15197 17153 15209 17187
rect 15243 17184 15255 17187
rect 15746 17184 15752 17196
rect 15243 17156 15752 17184
rect 15243 17153 15255 17156
rect 15197 17147 15255 17153
rect 15746 17144 15752 17156
rect 15804 17144 15810 17196
rect 16666 17144 16672 17196
rect 16724 17184 16730 17196
rect 18156 17184 18184 17224
rect 25958 17212 25964 17264
rect 26016 17252 26022 17264
rect 26053 17255 26111 17261
rect 26053 17252 26065 17255
rect 26016 17224 26065 17252
rect 26016 17212 26022 17224
rect 26053 17221 26065 17224
rect 26099 17221 26111 17255
rect 31570 17252 31576 17264
rect 26053 17215 26111 17221
rect 26160 17224 31576 17252
rect 18874 17184 18880 17196
rect 16724 17156 18184 17184
rect 18835 17156 18880 17184
rect 16724 17144 16730 17156
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17184 20131 17187
rect 20346 17184 20352 17196
rect 20119 17156 20352 17184
rect 20119 17153 20131 17156
rect 20073 17147 20131 17153
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 22554 17144 22560 17196
rect 22612 17184 22618 17196
rect 23017 17187 23075 17193
rect 23017 17184 23029 17187
rect 22612 17156 23029 17184
rect 22612 17144 22618 17156
rect 23017 17153 23029 17156
rect 23063 17153 23075 17187
rect 23017 17147 23075 17153
rect 23753 17187 23811 17193
rect 23753 17153 23765 17187
rect 23799 17184 23811 17187
rect 24762 17184 24768 17196
rect 23799 17156 24768 17184
rect 23799 17153 23811 17156
rect 23753 17147 23811 17153
rect 24762 17144 24768 17156
rect 24820 17144 24826 17196
rect 24946 17193 24952 17196
rect 24932 17187 24952 17193
rect 24932 17153 24944 17187
rect 24932 17147 24952 17153
rect 24946 17144 24952 17147
rect 25004 17144 25010 17196
rect 25225 17187 25283 17193
rect 25225 17153 25237 17187
rect 25271 17184 25283 17187
rect 26160 17184 26188 17224
rect 31570 17212 31576 17224
rect 31628 17212 31634 17264
rect 31726 17252 31754 17292
rect 32766 17280 32772 17332
rect 32824 17320 32830 17332
rect 33502 17320 33508 17332
rect 32824 17292 33508 17320
rect 32824 17280 32830 17292
rect 33502 17280 33508 17292
rect 33560 17280 33566 17332
rect 34146 17280 34152 17332
rect 34204 17320 34210 17332
rect 34701 17323 34759 17329
rect 34701 17320 34713 17323
rect 34204 17292 34713 17320
rect 34204 17280 34210 17292
rect 34701 17289 34713 17292
rect 34747 17289 34759 17323
rect 34701 17283 34759 17289
rect 35802 17280 35808 17332
rect 35860 17320 35866 17332
rect 37277 17323 37335 17329
rect 37277 17320 37289 17323
rect 35860 17292 37289 17320
rect 35860 17280 35866 17292
rect 37277 17289 37289 17292
rect 37323 17289 37335 17323
rect 37277 17283 37335 17289
rect 33134 17261 33140 17264
rect 33128 17252 33140 17261
rect 31726 17224 32996 17252
rect 33095 17224 33140 17252
rect 25271 17156 26188 17184
rect 26237 17187 26295 17193
rect 25271 17153 25283 17156
rect 25225 17147 25283 17153
rect 26237 17153 26249 17187
rect 26283 17184 26295 17187
rect 26970 17184 26976 17196
rect 26283 17156 26976 17184
rect 26283 17153 26295 17156
rect 26237 17147 26295 17153
rect 26970 17144 26976 17156
rect 27028 17144 27034 17196
rect 27157 17187 27215 17193
rect 27157 17153 27169 17187
rect 27203 17153 27215 17187
rect 27157 17147 27215 17153
rect 14108 17088 14596 17116
rect 14642 17076 14648 17128
rect 14700 17116 14706 17128
rect 14921 17119 14979 17125
rect 14921 17116 14933 17119
rect 14700 17088 14933 17116
rect 14700 17076 14706 17088
rect 14921 17085 14933 17088
rect 14967 17085 14979 17119
rect 14921 17079 14979 17085
rect 15930 17076 15936 17128
rect 15988 17116 15994 17128
rect 19981 17119 20039 17125
rect 15988 17088 19932 17116
rect 15988 17076 15994 17088
rect 16669 17051 16727 17057
rect 16669 17048 16681 17051
rect 14660 17020 16681 17048
rect 5353 16983 5411 16989
rect 5353 16949 5365 16983
rect 5399 16980 5411 16983
rect 6638 16980 6644 16992
rect 5399 16952 6644 16980
rect 5399 16949 5411 16952
rect 5353 16943 5411 16949
rect 6638 16940 6644 16952
rect 6696 16940 6702 16992
rect 7190 16940 7196 16992
rect 7248 16980 7254 16992
rect 7285 16983 7343 16989
rect 7285 16980 7297 16983
rect 7248 16952 7297 16980
rect 7248 16940 7254 16952
rect 7285 16949 7297 16952
rect 7331 16949 7343 16983
rect 7285 16943 7343 16949
rect 11514 16940 11520 16992
rect 11572 16980 11578 16992
rect 14660 16980 14688 17020
rect 16669 17017 16681 17020
rect 16715 17048 16727 17051
rect 16942 17048 16948 17060
rect 16715 17020 16948 17048
rect 16715 17017 16727 17020
rect 16669 17011 16727 17017
rect 16942 17008 16948 17020
rect 17000 17008 17006 17060
rect 17405 17051 17463 17057
rect 17405 17017 17417 17051
rect 17451 17048 17463 17051
rect 17954 17048 17960 17060
rect 17451 17020 17960 17048
rect 17451 17017 17463 17020
rect 17405 17011 17463 17017
rect 17954 17008 17960 17020
rect 18012 17048 18018 17060
rect 18874 17048 18880 17060
rect 18012 17020 18880 17048
rect 18012 17008 18018 17020
rect 18874 17008 18880 17020
rect 18932 17008 18938 17060
rect 19904 16989 19932 17088
rect 19981 17085 19993 17119
rect 20027 17116 20039 17119
rect 22741 17119 22799 17125
rect 20027 17088 22094 17116
rect 20027 17085 20039 17088
rect 19981 17079 20039 17085
rect 22066 17048 22094 17088
rect 22741 17085 22753 17119
rect 22787 17116 22799 17119
rect 23290 17116 23296 17128
rect 22787 17088 23296 17116
rect 22787 17085 22799 17088
rect 22741 17079 22799 17085
rect 23290 17076 23296 17088
rect 23348 17076 23354 17128
rect 23474 17116 23480 17128
rect 23435 17088 23480 17116
rect 23474 17076 23480 17088
rect 23532 17076 23538 17128
rect 25041 17119 25099 17125
rect 25041 17085 25053 17119
rect 25087 17085 25099 17119
rect 25041 17079 25099 17085
rect 24765 17051 24823 17057
rect 24765 17048 24777 17051
rect 22066 17020 24777 17048
rect 24765 17017 24777 17020
rect 24811 17017 24823 17051
rect 25056 17048 25084 17079
rect 25866 17076 25872 17128
rect 25924 17116 25930 17128
rect 27172 17116 27200 17147
rect 30926 17144 30932 17196
rect 30984 17184 30990 17196
rect 32861 17187 32919 17193
rect 32861 17184 32873 17187
rect 30984 17156 32873 17184
rect 30984 17144 30990 17156
rect 32861 17153 32873 17156
rect 32907 17153 32919 17187
rect 32968 17184 32996 17224
rect 33128 17215 33140 17224
rect 33134 17212 33140 17215
rect 33192 17212 33198 17264
rect 35066 17252 35072 17264
rect 34440 17224 35072 17252
rect 34440 17184 34468 17224
rect 35066 17212 35072 17224
rect 35124 17212 35130 17264
rect 39942 17252 39948 17264
rect 36096 17224 39948 17252
rect 32968 17156 34468 17184
rect 32861 17147 32919 17153
rect 34514 17144 34520 17196
rect 34572 17184 34578 17196
rect 36096 17193 36124 17224
rect 39942 17212 39948 17224
rect 40000 17212 40006 17264
rect 35814 17187 35872 17193
rect 35814 17184 35826 17187
rect 34572 17156 35826 17184
rect 34572 17144 34578 17156
rect 35814 17153 35826 17156
rect 35860 17153 35872 17187
rect 35814 17147 35872 17153
rect 36081 17187 36139 17193
rect 36081 17153 36093 17187
rect 36127 17153 36139 17187
rect 37458 17184 37464 17196
rect 37419 17156 37464 17184
rect 36081 17147 36139 17153
rect 37458 17144 37464 17156
rect 37516 17144 37522 17196
rect 37642 17184 37648 17196
rect 37603 17156 37648 17184
rect 37642 17144 37648 17156
rect 37700 17144 37706 17196
rect 39209 17187 39267 17193
rect 39209 17153 39221 17187
rect 39255 17184 39267 17187
rect 39758 17184 39764 17196
rect 39255 17156 39764 17184
rect 39255 17153 39267 17156
rect 39209 17147 39267 17153
rect 39758 17144 39764 17156
rect 39816 17144 39822 17196
rect 29454 17116 29460 17128
rect 25924 17088 27200 17116
rect 27264 17088 29460 17116
rect 25924 17076 25930 17088
rect 24765 17011 24823 17017
rect 24872 17020 25084 17048
rect 11572 16952 14688 16980
rect 19889 16983 19947 16989
rect 11572 16940 11578 16952
rect 19889 16949 19901 16983
rect 19935 16949 19947 16983
rect 19889 16943 19947 16949
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 21358 16980 21364 16992
rect 21315 16952 21364 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21358 16940 21364 16952
rect 21416 16980 21422 16992
rect 21818 16980 21824 16992
rect 21416 16952 21824 16980
rect 21416 16940 21422 16952
rect 21818 16940 21824 16952
rect 21876 16940 21882 16992
rect 23382 16940 23388 16992
rect 23440 16980 23446 16992
rect 24872 16980 24900 17020
rect 25682 17008 25688 17060
rect 25740 17048 25746 17060
rect 27264 17048 27292 17088
rect 29454 17076 29460 17088
rect 29512 17076 29518 17128
rect 30374 17076 30380 17128
rect 30432 17116 30438 17128
rect 30745 17119 30803 17125
rect 30745 17116 30757 17119
rect 30432 17088 30757 17116
rect 30432 17076 30438 17088
rect 30745 17085 30757 17088
rect 30791 17085 30803 17119
rect 30745 17079 30803 17085
rect 31021 17119 31079 17125
rect 31021 17085 31033 17119
rect 31067 17116 31079 17119
rect 32674 17116 32680 17128
rect 31067 17088 32680 17116
rect 31067 17085 31079 17088
rect 31021 17079 31079 17085
rect 32674 17076 32680 17088
rect 32732 17076 32738 17128
rect 39485 17119 39543 17125
rect 39485 17085 39497 17119
rect 39531 17116 39543 17119
rect 39850 17116 39856 17128
rect 39531 17088 39856 17116
rect 39531 17085 39543 17088
rect 39485 17079 39543 17085
rect 39850 17076 39856 17088
rect 39908 17076 39914 17128
rect 25740 17020 27292 17048
rect 27341 17051 27399 17057
rect 25740 17008 25746 17020
rect 27341 17017 27353 17051
rect 27387 17048 27399 17051
rect 28166 17048 28172 17060
rect 27387 17020 28172 17048
rect 27387 17017 27399 17020
rect 27341 17011 27399 17017
rect 28166 17008 28172 17020
rect 28224 17008 28230 17060
rect 33870 17008 33876 17060
rect 33928 17048 33934 17060
rect 34241 17051 34299 17057
rect 34241 17048 34253 17051
rect 33928 17020 34253 17048
rect 33928 17008 33934 17020
rect 34241 17017 34253 17020
rect 34287 17017 34299 17051
rect 58158 17048 58164 17060
rect 58119 17020 58164 17048
rect 34241 17011 34299 17017
rect 58158 17008 58164 17020
rect 58216 17008 58222 17060
rect 25130 16980 25136 16992
rect 23440 16952 24900 16980
rect 25091 16952 25136 16980
rect 23440 16940 23446 16952
rect 25130 16940 25136 16952
rect 25188 16940 25194 16992
rect 27798 16940 27804 16992
rect 27856 16980 27862 16992
rect 27893 16983 27951 16989
rect 27893 16980 27905 16983
rect 27856 16952 27905 16980
rect 27856 16940 27862 16952
rect 27893 16949 27905 16952
rect 27939 16980 27951 16983
rect 28626 16980 28632 16992
rect 27939 16952 28632 16980
rect 27939 16949 27951 16952
rect 27893 16943 27951 16949
rect 28626 16940 28632 16952
rect 28684 16940 28690 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 7282 16736 7288 16788
rect 7340 16776 7346 16788
rect 7742 16776 7748 16788
rect 7340 16748 7748 16776
rect 7340 16736 7346 16748
rect 7742 16736 7748 16748
rect 7800 16736 7806 16788
rect 8018 16776 8024 16788
rect 7979 16748 8024 16776
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 12158 16736 12164 16788
rect 12216 16776 12222 16788
rect 14921 16779 14979 16785
rect 14921 16776 14933 16779
rect 12216 16748 14933 16776
rect 12216 16736 12222 16748
rect 14921 16745 14933 16748
rect 14967 16776 14979 16779
rect 15746 16776 15752 16788
rect 14967 16748 15752 16776
rect 14967 16745 14979 16748
rect 14921 16739 14979 16745
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 20625 16779 20683 16785
rect 20625 16776 20637 16779
rect 16356 16748 20637 16776
rect 16356 16736 16362 16748
rect 20625 16745 20637 16748
rect 20671 16776 20683 16779
rect 25866 16776 25872 16788
rect 20671 16748 21128 16776
rect 25827 16748 25872 16776
rect 20671 16745 20683 16748
rect 20625 16739 20683 16745
rect 5626 16708 5632 16720
rect 5092 16680 5632 16708
rect 5092 16649 5120 16680
rect 5626 16668 5632 16680
rect 5684 16668 5690 16720
rect 7374 16668 7380 16720
rect 7432 16708 7438 16720
rect 7432 16680 7696 16708
rect 7432 16668 7438 16680
rect 7668 16649 7696 16680
rect 16758 16668 16764 16720
rect 16816 16708 16822 16720
rect 21100 16717 21128 16748
rect 25866 16736 25872 16748
rect 25924 16736 25930 16788
rect 28350 16736 28356 16788
rect 28408 16776 28414 16788
rect 32306 16776 32312 16788
rect 28408 16748 32312 16776
rect 28408 16736 28414 16748
rect 32306 16736 32312 16748
rect 32364 16736 32370 16788
rect 38102 16776 38108 16788
rect 36004 16748 38108 16776
rect 21085 16711 21143 16717
rect 16816 16680 18092 16708
rect 16816 16668 16822 16680
rect 5077 16643 5135 16649
rect 5077 16609 5089 16643
rect 5123 16609 5135 16643
rect 5077 16603 5135 16609
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16640 5319 16643
rect 7561 16643 7619 16649
rect 7561 16640 7573 16643
rect 5307 16612 7573 16640
rect 5307 16609 5319 16612
rect 5261 16603 5319 16609
rect 7561 16609 7573 16612
rect 7607 16609 7619 16643
rect 7561 16603 7619 16609
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16609 7711 16643
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 7653 16603 7711 16609
rect 7852 16612 8953 16640
rect 2409 16575 2467 16581
rect 2409 16541 2421 16575
rect 2455 16572 2467 16575
rect 2498 16572 2504 16584
rect 2455 16544 2504 16572
rect 2455 16541 2467 16544
rect 2409 16535 2467 16541
rect 2498 16532 2504 16544
rect 2556 16532 2562 16584
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4985 16575 5043 16581
rect 4985 16572 4997 16575
rect 4396 16544 4997 16572
rect 4396 16532 4402 16544
rect 4985 16541 4997 16544
rect 5031 16541 5043 16575
rect 7282 16572 7288 16584
rect 7243 16544 7288 16572
rect 4985 16535 5043 16541
rect 7282 16532 7288 16544
rect 7340 16532 7346 16584
rect 7466 16572 7472 16584
rect 7427 16544 7472 16572
rect 7466 16532 7472 16544
rect 7524 16532 7530 16584
rect 7852 16581 7880 16612
rect 8941 16609 8953 16612
rect 8987 16609 8999 16643
rect 8941 16603 8999 16609
rect 12529 16643 12587 16649
rect 12529 16609 12541 16643
rect 12575 16640 12587 16643
rect 12618 16640 12624 16652
rect 12575 16612 12624 16640
rect 12575 16609 12587 16612
rect 12529 16603 12587 16609
rect 12618 16600 12624 16612
rect 12676 16640 12682 16652
rect 16298 16640 16304 16652
rect 12676 16612 16304 16640
rect 12676 16600 12682 16612
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 17954 16640 17960 16652
rect 16592 16612 17960 16640
rect 7837 16575 7895 16581
rect 7837 16541 7849 16575
rect 7883 16574 7895 16575
rect 7883 16546 7917 16574
rect 15746 16572 15752 16584
rect 7883 16541 7895 16546
rect 15707 16544 15752 16572
rect 7837 16535 7895 16541
rect 3970 16464 3976 16516
rect 4028 16504 4034 16516
rect 7190 16504 7196 16516
rect 4028 16476 7196 16504
rect 4028 16464 4034 16476
rect 7190 16464 7196 16476
rect 7248 16504 7254 16516
rect 7852 16504 7880 16535
rect 15746 16532 15752 16544
rect 15804 16532 15810 16584
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 14182 16504 14188 16516
rect 7248 16476 7880 16504
rect 10520 16476 14188 16504
rect 7248 16464 7254 16476
rect 2225 16439 2283 16445
rect 2225 16405 2237 16439
rect 2271 16436 2283 16439
rect 2314 16436 2320 16448
rect 2271 16408 2320 16436
rect 2271 16405 2283 16408
rect 2225 16399 2283 16405
rect 2314 16396 2320 16408
rect 2372 16396 2378 16448
rect 4617 16439 4675 16445
rect 4617 16405 4629 16439
rect 4663 16436 4675 16439
rect 4706 16436 4712 16448
rect 4663 16408 4712 16436
rect 4663 16405 4675 16408
rect 4617 16399 4675 16405
rect 4706 16396 4712 16408
rect 4764 16436 4770 16448
rect 5258 16436 5264 16448
rect 4764 16408 5264 16436
rect 4764 16396 4770 16408
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 8478 16396 8484 16448
rect 8536 16436 8542 16448
rect 9953 16439 10011 16445
rect 9953 16436 9965 16439
rect 8536 16408 9965 16436
rect 8536 16396 8542 16408
rect 9953 16405 9965 16408
rect 9999 16436 10011 16439
rect 10318 16436 10324 16448
rect 9999 16408 10324 16436
rect 9999 16405 10011 16408
rect 9953 16399 10011 16405
rect 10318 16396 10324 16408
rect 10376 16436 10382 16448
rect 10520 16445 10548 16476
rect 14182 16464 14188 16476
rect 14240 16464 14246 16516
rect 15856 16504 15884 16535
rect 15930 16532 15936 16584
rect 15988 16572 15994 16584
rect 15988 16544 16033 16572
rect 15988 16532 15994 16544
rect 16114 16532 16120 16584
rect 16172 16572 16178 16584
rect 16592 16581 16620 16612
rect 17954 16600 17960 16612
rect 18012 16600 18018 16652
rect 18064 16640 18092 16680
rect 21085 16677 21097 16711
rect 21131 16708 21143 16711
rect 21174 16708 21180 16720
rect 21131 16680 21180 16708
rect 21131 16677 21143 16680
rect 21085 16671 21143 16677
rect 21174 16668 21180 16680
rect 21232 16668 21238 16720
rect 19981 16643 20039 16649
rect 19981 16640 19993 16643
rect 18064 16612 19993 16640
rect 19981 16609 19993 16612
rect 20027 16640 20039 16643
rect 20990 16640 20996 16652
rect 20027 16612 20996 16640
rect 20027 16609 20039 16612
rect 19981 16603 20039 16609
rect 20990 16600 20996 16612
rect 21048 16600 21054 16652
rect 22370 16600 22376 16652
rect 22428 16640 22434 16652
rect 22646 16640 22652 16652
rect 22428 16612 22652 16640
rect 22428 16600 22434 16612
rect 22646 16600 22652 16612
rect 22704 16640 22710 16652
rect 22833 16643 22891 16649
rect 22833 16640 22845 16643
rect 22704 16612 22845 16640
rect 22704 16600 22710 16612
rect 22833 16609 22845 16612
rect 22879 16609 22891 16643
rect 27246 16640 27252 16652
rect 27207 16612 27252 16640
rect 22833 16603 22891 16609
rect 27246 16600 27252 16612
rect 27304 16600 27310 16652
rect 27338 16600 27344 16652
rect 27396 16640 27402 16652
rect 27798 16640 27804 16652
rect 27396 16612 27804 16640
rect 27396 16600 27402 16612
rect 27798 16600 27804 16612
rect 27856 16640 27862 16652
rect 27856 16612 27936 16640
rect 27856 16600 27862 16612
rect 16577 16575 16635 16581
rect 16577 16572 16589 16575
rect 16172 16544 16589 16572
rect 16172 16532 16178 16544
rect 16577 16541 16589 16544
rect 16623 16541 16635 16575
rect 16758 16572 16764 16584
rect 16719 16544 16764 16572
rect 16577 16535 16635 16541
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16541 16911 16575
rect 16853 16535 16911 16541
rect 16868 16504 16896 16535
rect 16942 16532 16948 16584
rect 17000 16572 17006 16584
rect 17972 16572 18000 16600
rect 18049 16575 18107 16581
rect 18049 16572 18061 16575
rect 17000 16544 17045 16572
rect 17972 16544 18061 16572
rect 17000 16532 17006 16544
rect 18049 16541 18061 16544
rect 18095 16541 18107 16575
rect 18230 16572 18236 16584
rect 18191 16544 18236 16572
rect 18049 16535 18107 16541
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 18325 16575 18383 16581
rect 18325 16541 18337 16575
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16541 18475 16575
rect 22554 16572 22560 16584
rect 22515 16544 22560 16572
rect 18417 16535 18475 16541
rect 17770 16504 17776 16516
rect 15856 16476 17776 16504
rect 17770 16464 17776 16476
rect 17828 16504 17834 16516
rect 18340 16504 18368 16535
rect 17828 16476 18368 16504
rect 17828 16464 17834 16476
rect 10505 16439 10563 16445
rect 10505 16436 10517 16439
rect 10376 16408 10517 16436
rect 10376 16396 10382 16408
rect 10505 16405 10517 16408
rect 10551 16405 10563 16439
rect 11146 16436 11152 16448
rect 11107 16408 11152 16436
rect 10505 16399 10563 16405
rect 11146 16396 11152 16408
rect 11204 16396 11210 16448
rect 12802 16396 12808 16448
rect 12860 16436 12866 16448
rect 12989 16439 13047 16445
rect 12989 16436 13001 16439
rect 12860 16408 13001 16436
rect 12860 16396 12866 16408
rect 12989 16405 13001 16408
rect 13035 16405 13047 16439
rect 12989 16399 13047 16405
rect 15378 16396 15384 16448
rect 15436 16436 15442 16448
rect 15473 16439 15531 16445
rect 15473 16436 15485 16439
rect 15436 16408 15485 16436
rect 15436 16396 15442 16408
rect 15473 16405 15485 16408
rect 15519 16405 15531 16439
rect 17218 16436 17224 16448
rect 17179 16408 17224 16436
rect 15473 16399 15531 16405
rect 17218 16396 17224 16408
rect 17276 16396 17282 16448
rect 18046 16396 18052 16448
rect 18104 16436 18110 16448
rect 18432 16436 18460 16535
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 27908 16572 27936 16612
rect 28092 16612 28580 16640
rect 28092 16581 28120 16612
rect 27965 16575 28023 16581
rect 27965 16572 27977 16575
rect 27908 16544 27977 16572
rect 27965 16541 27977 16544
rect 28011 16541 28023 16575
rect 27965 16535 28023 16541
rect 28074 16575 28132 16581
rect 28074 16541 28086 16575
rect 28120 16541 28132 16575
rect 28074 16535 28132 16541
rect 28166 16532 28172 16584
rect 28224 16572 28230 16584
rect 28224 16544 28269 16572
rect 28224 16532 28230 16544
rect 28350 16532 28356 16584
rect 28408 16572 28414 16584
rect 28408 16544 28453 16572
rect 28408 16532 28414 16544
rect 27004 16507 27062 16513
rect 27004 16473 27016 16507
rect 27050 16504 27062 16507
rect 27709 16507 27767 16513
rect 27709 16504 27721 16507
rect 27050 16476 27721 16504
rect 27050 16473 27062 16476
rect 27004 16467 27062 16473
rect 27709 16473 27721 16476
rect 27755 16473 27767 16507
rect 27709 16467 27767 16473
rect 18690 16436 18696 16448
rect 18104 16408 18460 16436
rect 18651 16408 18696 16436
rect 18104 16396 18110 16408
rect 18690 16396 18696 16408
rect 18748 16396 18754 16448
rect 19426 16436 19432 16448
rect 19387 16408 19432 16436
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 22094 16396 22100 16448
rect 22152 16436 22158 16448
rect 22152 16408 22197 16436
rect 22152 16396 22158 16408
rect 27154 16396 27160 16448
rect 27212 16436 27218 16448
rect 28552 16436 28580 16612
rect 32674 16600 32680 16652
rect 32732 16640 32738 16652
rect 36004 16649 36032 16748
rect 38102 16736 38108 16748
rect 38160 16736 38166 16788
rect 38194 16736 38200 16788
rect 38252 16776 38258 16788
rect 38930 16776 38936 16788
rect 38252 16748 38936 16776
rect 38252 16736 38258 16748
rect 38930 16736 38936 16748
rect 38988 16736 38994 16788
rect 40313 16779 40371 16785
rect 40313 16745 40325 16779
rect 40359 16776 40371 16779
rect 40770 16776 40776 16788
rect 40359 16748 40776 16776
rect 40359 16745 40371 16748
rect 40313 16739 40371 16745
rect 40770 16736 40776 16748
rect 40828 16736 40834 16788
rect 37369 16711 37427 16717
rect 37369 16677 37381 16711
rect 37415 16708 37427 16711
rect 37458 16708 37464 16720
rect 37415 16680 37464 16708
rect 37415 16677 37427 16680
rect 37369 16671 37427 16677
rect 37458 16668 37464 16680
rect 37516 16668 37522 16720
rect 35989 16643 36047 16649
rect 32732 16612 33088 16640
rect 32732 16600 32738 16612
rect 28626 16532 28632 16584
rect 28684 16572 28690 16584
rect 28684 16544 30880 16572
rect 28684 16532 28690 16544
rect 30374 16504 30380 16516
rect 28966 16476 30380 16504
rect 28966 16436 28994 16476
rect 30374 16464 30380 16476
rect 30432 16464 30438 16516
rect 30558 16464 30564 16516
rect 30616 16504 30622 16516
rect 30754 16507 30812 16513
rect 30754 16504 30766 16507
rect 30616 16476 30766 16504
rect 30616 16464 30622 16476
rect 30754 16473 30766 16476
rect 30800 16473 30812 16507
rect 30852 16504 30880 16544
rect 30926 16532 30932 16584
rect 30984 16572 30990 16584
rect 31021 16575 31079 16581
rect 31021 16572 31033 16575
rect 30984 16544 31033 16572
rect 30984 16532 30990 16544
rect 31021 16541 31033 16544
rect 31067 16541 31079 16575
rect 31021 16535 31079 16541
rect 32030 16532 32036 16584
rect 32088 16572 32094 16584
rect 32490 16572 32496 16584
rect 32088 16544 32496 16572
rect 32088 16532 32094 16544
rect 32490 16532 32496 16544
rect 32548 16572 32554 16584
rect 32769 16575 32827 16581
rect 32769 16572 32781 16575
rect 32548 16544 32781 16572
rect 32548 16532 32554 16544
rect 32769 16541 32781 16544
rect 32815 16541 32827 16575
rect 32950 16572 32956 16584
rect 32911 16544 32956 16572
rect 32769 16535 32827 16541
rect 32950 16532 32956 16544
rect 33008 16532 33014 16584
rect 33060 16581 33088 16612
rect 35989 16609 36001 16643
rect 36035 16609 36047 16643
rect 35989 16603 36047 16609
rect 33045 16575 33103 16581
rect 33045 16541 33057 16575
rect 33091 16541 33103 16575
rect 33045 16535 33103 16541
rect 33137 16575 33195 16581
rect 33137 16541 33149 16575
rect 33183 16572 33195 16575
rect 33962 16572 33968 16584
rect 33183 16544 33968 16572
rect 33183 16541 33195 16544
rect 33137 16535 33195 16541
rect 31478 16504 31484 16516
rect 30852 16476 31484 16504
rect 30754 16467 30812 16473
rect 31478 16464 31484 16476
rect 31536 16464 31542 16516
rect 32306 16504 32312 16516
rect 32219 16476 32312 16504
rect 32306 16464 32312 16476
rect 32364 16504 32370 16516
rect 33152 16504 33180 16535
rect 33962 16532 33968 16544
rect 34020 16532 34026 16584
rect 36262 16581 36268 16584
rect 36256 16572 36268 16581
rect 36223 16544 36268 16572
rect 36256 16535 36268 16544
rect 36262 16532 36268 16535
rect 36320 16532 36326 16584
rect 32364 16476 33180 16504
rect 33413 16507 33471 16513
rect 32364 16464 32370 16476
rect 33413 16473 33425 16507
rect 33459 16504 33471 16507
rect 34514 16504 34520 16516
rect 33459 16476 34520 16504
rect 33459 16473 33471 16476
rect 33413 16467 33471 16473
rect 34514 16464 34520 16476
rect 34572 16464 34578 16516
rect 40405 16507 40463 16513
rect 40405 16473 40417 16507
rect 40451 16504 40463 16507
rect 40494 16504 40500 16516
rect 40451 16476 40500 16504
rect 40451 16473 40463 16476
rect 40405 16467 40463 16473
rect 40494 16464 40500 16476
rect 40552 16464 40558 16516
rect 27212 16408 28994 16436
rect 29641 16439 29699 16445
rect 27212 16396 27218 16408
rect 29641 16405 29653 16439
rect 29687 16436 29699 16439
rect 29822 16436 29828 16448
rect 29687 16408 29828 16436
rect 29687 16405 29699 16408
rect 29641 16399 29699 16405
rect 29822 16396 29828 16408
rect 29880 16396 29886 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 3421 16235 3479 16241
rect 3421 16201 3433 16235
rect 3467 16232 3479 16235
rect 4338 16232 4344 16244
rect 3467 16204 4344 16232
rect 3467 16201 3479 16204
rect 3421 16195 3479 16201
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 5169 16235 5227 16241
rect 5169 16201 5181 16235
rect 5215 16232 5227 16235
rect 6178 16232 6184 16244
rect 5215 16204 6184 16232
rect 5215 16201 5227 16204
rect 5169 16195 5227 16201
rect 2866 16164 2872 16176
rect 2056 16136 2872 16164
rect 2056 16105 2084 16136
rect 2866 16124 2872 16136
rect 2924 16124 2930 16176
rect 4249 16167 4307 16173
rect 4249 16133 4261 16167
rect 4295 16164 4307 16167
rect 5184 16164 5212 16195
rect 6178 16192 6184 16204
rect 6236 16192 6242 16244
rect 10870 16232 10876 16244
rect 10831 16204 10876 16232
rect 10870 16192 10876 16204
rect 10928 16192 10934 16244
rect 12713 16235 12771 16241
rect 12713 16201 12725 16235
rect 12759 16232 12771 16235
rect 13722 16232 13728 16244
rect 12759 16204 13728 16232
rect 12759 16201 12771 16204
rect 12713 16195 12771 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 15930 16192 15936 16244
rect 15988 16232 15994 16244
rect 16669 16235 16727 16241
rect 16669 16232 16681 16235
rect 15988 16204 16681 16232
rect 15988 16192 15994 16204
rect 16669 16201 16681 16204
rect 16715 16201 16727 16235
rect 16669 16195 16727 16201
rect 16758 16192 16764 16244
rect 16816 16232 16822 16244
rect 17497 16235 17555 16241
rect 17497 16232 17509 16235
rect 16816 16204 17509 16232
rect 16816 16192 16822 16204
rect 17497 16201 17509 16204
rect 17543 16201 17555 16235
rect 17497 16195 17555 16201
rect 18230 16192 18236 16244
rect 18288 16232 18294 16244
rect 19061 16235 19119 16241
rect 19061 16232 19073 16235
rect 18288 16204 19073 16232
rect 18288 16192 18294 16204
rect 19061 16201 19073 16204
rect 19107 16201 19119 16235
rect 19061 16195 19119 16201
rect 20809 16235 20867 16241
rect 20809 16201 20821 16235
rect 20855 16232 20867 16235
rect 26326 16232 26332 16244
rect 20855 16204 26332 16232
rect 20855 16201 20867 16204
rect 20809 16195 20867 16201
rect 26326 16192 26332 16204
rect 26384 16192 26390 16244
rect 26970 16192 26976 16244
rect 27028 16232 27034 16244
rect 27157 16235 27215 16241
rect 27157 16232 27169 16235
rect 27028 16204 27169 16232
rect 27028 16192 27034 16204
rect 27157 16201 27169 16204
rect 27203 16232 27215 16235
rect 31386 16232 31392 16244
rect 27203 16204 31392 16232
rect 27203 16201 27215 16204
rect 27157 16195 27215 16201
rect 31386 16192 31392 16204
rect 31444 16192 31450 16244
rect 31478 16192 31484 16244
rect 31536 16232 31542 16244
rect 37277 16235 37335 16241
rect 31536 16204 35112 16232
rect 31536 16192 31542 16204
rect 4295 16136 5212 16164
rect 11885 16167 11943 16173
rect 4295 16133 4307 16136
rect 4249 16127 4307 16133
rect 11885 16133 11897 16167
rect 11931 16164 11943 16167
rect 15010 16164 15016 16176
rect 11931 16136 15016 16164
rect 11931 16133 11943 16136
rect 11885 16127 11943 16133
rect 15010 16124 15016 16136
rect 15068 16124 15074 16176
rect 16114 16164 16120 16176
rect 16075 16136 16120 16164
rect 16114 16124 16120 16136
rect 16172 16124 16178 16176
rect 17037 16167 17095 16173
rect 17037 16133 17049 16167
rect 17083 16164 17095 16167
rect 17865 16167 17923 16173
rect 17865 16164 17877 16167
rect 17083 16136 17877 16164
rect 17083 16133 17095 16136
rect 17037 16127 17095 16133
rect 17865 16133 17877 16136
rect 17911 16164 17923 16167
rect 19334 16164 19340 16176
rect 17911 16136 19340 16164
rect 17911 16133 17923 16136
rect 17865 16127 17923 16133
rect 19334 16124 19340 16136
rect 19392 16164 19398 16176
rect 19429 16167 19487 16173
rect 19429 16164 19441 16167
rect 19392 16136 19441 16164
rect 19392 16124 19398 16136
rect 19429 16133 19441 16136
rect 19475 16133 19487 16167
rect 19429 16127 19487 16133
rect 19886 16124 19892 16176
rect 19944 16164 19950 16176
rect 19944 16136 26188 16164
rect 19944 16124 19950 16136
rect 2314 16105 2320 16108
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16065 2099 16099
rect 2308 16096 2320 16105
rect 2275 16068 2320 16096
rect 2041 16059 2099 16065
rect 2308 16059 2320 16068
rect 2314 16056 2320 16059
rect 2372 16056 2378 16108
rect 10137 16099 10195 16105
rect 10137 16065 10149 16099
rect 10183 16065 10195 16099
rect 10318 16096 10324 16108
rect 10279 16068 10324 16096
rect 10137 16059 10195 16065
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 16028 4583 16031
rect 4706 16028 4712 16040
rect 4571 16000 4712 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 10152 16028 10180 16059
rect 10318 16056 10324 16068
rect 10376 16096 10382 16108
rect 10781 16099 10839 16105
rect 10781 16096 10793 16099
rect 10376 16068 10793 16096
rect 10376 16056 10382 16068
rect 10781 16065 10793 16068
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16065 11023 16099
rect 10965 16059 11023 16065
rect 10980 16028 11008 16059
rect 11422 16056 11428 16108
rect 11480 16096 11486 16108
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 11480 16068 11529 16096
rect 11480 16056 11486 16068
rect 11517 16065 11529 16068
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 11664 16068 11709 16096
rect 11664 16056 11670 16068
rect 11790 16056 11796 16108
rect 11848 16096 11854 16108
rect 11974 16096 11980 16108
rect 11848 16068 11893 16096
rect 11933 16068 11980 16096
rect 11848 16056 11854 16068
rect 11974 16056 11980 16068
rect 12032 16105 12038 16108
rect 12032 16099 12081 16105
rect 12032 16065 12035 16099
rect 12069 16096 12081 16099
rect 12618 16096 12624 16108
rect 12069 16068 12434 16096
rect 12579 16068 12624 16096
rect 12069 16065 12081 16068
rect 12032 16059 12081 16065
rect 12032 16056 12038 16059
rect 11146 16028 11152 16040
rect 9723 16000 10916 16028
rect 10980 16000 11152 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 10321 15963 10379 15969
rect 10321 15929 10333 15963
rect 10367 15960 10379 15963
rect 10778 15960 10784 15972
rect 10367 15932 10784 15960
rect 10367 15929 10379 15932
rect 10321 15923 10379 15929
rect 10778 15920 10784 15932
rect 10836 15920 10842 15972
rect 10888 15960 10916 16000
rect 11146 15988 11152 16000
rect 11204 16028 11210 16040
rect 11698 16028 11704 16040
rect 11204 16000 11704 16028
rect 11204 15988 11210 16000
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 12406 16028 12434 16068
rect 12618 16056 12624 16068
rect 12676 16056 12682 16108
rect 12802 16096 12808 16108
rect 12763 16068 12808 16096
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 13814 16056 13820 16108
rect 13872 16056 13878 16108
rect 14274 16096 14280 16108
rect 14187 16068 14280 16096
rect 14274 16056 14280 16068
rect 14332 16096 14338 16108
rect 14642 16096 14648 16108
rect 14332 16068 14648 16096
rect 14332 16056 14338 16068
rect 14642 16056 14648 16068
rect 14700 16056 14706 16108
rect 16853 16099 16911 16105
rect 16853 16065 16865 16099
rect 16899 16096 16911 16099
rect 16942 16096 16948 16108
rect 16899 16068 16948 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 17681 16099 17739 16105
rect 17681 16065 17693 16099
rect 17727 16096 17739 16099
rect 18230 16096 18236 16108
rect 17727 16068 18236 16096
rect 17727 16065 17739 16068
rect 17681 16059 17739 16065
rect 18230 16056 18236 16068
rect 18288 16056 18294 16108
rect 19245 16099 19303 16105
rect 19245 16065 19257 16099
rect 19291 16096 19303 16099
rect 19291 16068 20024 16096
rect 19291 16065 19303 16068
rect 19245 16059 19303 16065
rect 13832 16028 13860 16056
rect 14550 16028 14556 16040
rect 12406 16000 13860 16028
rect 14511 16000 14556 16028
rect 14550 15988 14556 16000
rect 14608 15988 14614 16040
rect 19426 15988 19432 16040
rect 19484 16028 19490 16040
rect 19886 16028 19892 16040
rect 19484 16000 19892 16028
rect 19484 15988 19490 16000
rect 19886 15988 19892 16000
rect 19944 15988 19950 16040
rect 19996 16028 20024 16068
rect 20070 16056 20076 16108
rect 20128 16096 20134 16108
rect 20717 16099 20775 16105
rect 20128 16068 20173 16096
rect 20128 16056 20134 16068
rect 20717 16065 20729 16099
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16096 20959 16099
rect 20990 16096 20996 16108
rect 20947 16068 20996 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 20622 16028 20628 16040
rect 19996 16000 20628 16028
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 20732 16028 20760 16059
rect 20990 16056 20996 16068
rect 21048 16056 21054 16108
rect 23017 16099 23075 16105
rect 23017 16065 23029 16099
rect 23063 16096 23075 16099
rect 23474 16096 23480 16108
rect 23063 16068 23480 16096
rect 23063 16065 23075 16068
rect 23017 16059 23075 16065
rect 23474 16056 23480 16068
rect 23532 16056 23538 16108
rect 26160 16096 26188 16136
rect 26234 16124 26240 16176
rect 26292 16164 26298 16176
rect 26292 16136 32628 16164
rect 26292 16124 26298 16136
rect 26160 16068 26464 16096
rect 21174 16028 21180 16040
rect 20732 16000 21180 16028
rect 21174 15988 21180 16000
rect 21232 15988 21238 16040
rect 26436 16037 26464 16068
rect 27154 16056 27160 16108
rect 27212 16096 27218 16108
rect 27341 16099 27399 16105
rect 27341 16096 27353 16099
rect 27212 16068 27353 16096
rect 27212 16056 27218 16068
rect 27341 16065 27353 16068
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 29089 16099 29147 16105
rect 29089 16065 29101 16099
rect 29135 16065 29147 16099
rect 29089 16059 29147 16065
rect 29273 16099 29331 16105
rect 29273 16065 29285 16099
rect 29319 16096 29331 16099
rect 29822 16096 29828 16108
rect 29319 16068 29828 16096
rect 29319 16065 29331 16068
rect 29273 16059 29331 16065
rect 23293 16031 23351 16037
rect 23293 15997 23305 16031
rect 23339 15997 23351 16031
rect 23293 15991 23351 15997
rect 26421 16031 26479 16037
rect 26421 15997 26433 16031
rect 26467 16028 26479 16031
rect 27522 16028 27528 16040
rect 26467 16000 27528 16028
rect 26467 15997 26479 16000
rect 26421 15991 26479 15997
rect 13817 15963 13875 15969
rect 10888 15932 12296 15960
rect 3878 15892 3884 15904
rect 3839 15864 3884 15892
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 7098 15892 7104 15904
rect 7059 15864 7104 15892
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 12161 15895 12219 15901
rect 12161 15892 12173 15895
rect 9732 15864 12173 15892
rect 9732 15852 9738 15864
rect 12161 15861 12173 15864
rect 12207 15861 12219 15895
rect 12268 15892 12296 15932
rect 13817 15929 13829 15963
rect 13863 15960 13875 15963
rect 14182 15960 14188 15972
rect 13863 15932 14188 15960
rect 13863 15929 13875 15932
rect 13817 15923 13875 15929
rect 14182 15920 14188 15932
rect 14240 15960 14246 15972
rect 22094 15960 22100 15972
rect 14240 15932 22100 15960
rect 14240 15920 14246 15932
rect 22094 15920 22100 15932
rect 22152 15920 22158 15972
rect 23198 15920 23204 15972
rect 23256 15960 23262 15972
rect 23308 15960 23336 15991
rect 27522 15988 27528 16000
rect 27580 15988 27586 16040
rect 27154 15960 27160 15972
rect 23256 15932 27160 15960
rect 23256 15920 23262 15932
rect 27154 15920 27160 15932
rect 27212 15920 27218 15972
rect 29104 15960 29132 16059
rect 29822 16056 29828 16068
rect 29880 16056 29886 16108
rect 30374 16056 30380 16108
rect 30432 16096 30438 16108
rect 30745 16099 30803 16105
rect 30745 16096 30757 16099
rect 30432 16068 30757 16096
rect 30432 16056 30438 16068
rect 30745 16065 30757 16068
rect 30791 16065 30803 16099
rect 31386 16096 31392 16108
rect 31347 16068 31392 16096
rect 30745 16059 30803 16065
rect 31386 16056 31392 16068
rect 31444 16056 31450 16108
rect 29914 15988 29920 16040
rect 29972 16028 29978 16040
rect 30469 16031 30527 16037
rect 30469 16028 30481 16031
rect 29972 16000 30481 16028
rect 29972 15988 29978 16000
rect 30469 15997 30481 16000
rect 30515 16028 30527 16031
rect 30650 16028 30656 16040
rect 30515 16000 30656 16028
rect 30515 15997 30527 16000
rect 30469 15991 30527 15997
rect 30650 15988 30656 16000
rect 30708 15988 30714 16040
rect 30926 15988 30932 16040
rect 30984 16028 30990 16040
rect 32493 16031 32551 16037
rect 32493 16028 32505 16031
rect 30984 16000 32505 16028
rect 30984 15988 30990 16000
rect 32493 15997 32505 16000
rect 32539 15997 32551 16031
rect 32493 15991 32551 15997
rect 29822 15960 29828 15972
rect 29104 15932 29828 15960
rect 29822 15920 29828 15932
rect 29880 15960 29886 15972
rect 31205 15963 31263 15969
rect 31205 15960 31217 15963
rect 29880 15932 31217 15960
rect 29880 15920 29886 15932
rect 31205 15929 31217 15932
rect 31251 15929 31263 15963
rect 31205 15923 31263 15929
rect 32600 15904 32628 16136
rect 34241 16099 34299 16105
rect 34241 16065 34253 16099
rect 34287 16065 34299 16099
rect 34241 16059 34299 16065
rect 12802 15892 12808 15904
rect 12268 15864 12808 15892
rect 12161 15855 12219 15861
rect 12802 15852 12808 15864
rect 12860 15852 12866 15904
rect 20257 15895 20315 15901
rect 20257 15861 20269 15895
rect 20303 15892 20315 15895
rect 21450 15892 21456 15904
rect 20303 15864 21456 15892
rect 20303 15861 20315 15864
rect 20257 15855 20315 15861
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 22186 15852 22192 15904
rect 22244 15892 22250 15904
rect 22281 15895 22339 15901
rect 22281 15892 22293 15895
rect 22244 15864 22293 15892
rect 22244 15852 22250 15864
rect 22281 15861 22293 15864
rect 22327 15861 22339 15895
rect 22281 15855 22339 15861
rect 29457 15895 29515 15901
rect 29457 15861 29469 15895
rect 29503 15892 29515 15895
rect 30374 15892 30380 15904
rect 29503 15864 30380 15892
rect 29503 15861 29515 15864
rect 29457 15855 29515 15861
rect 30374 15852 30380 15864
rect 30432 15852 30438 15904
rect 32582 15852 32588 15904
rect 32640 15892 32646 15904
rect 34256 15892 34284 16059
rect 35084 15960 35112 16204
rect 37277 16201 37289 16235
rect 37323 16232 37335 16235
rect 37366 16232 37372 16244
rect 37323 16204 37372 16232
rect 37323 16201 37335 16204
rect 37277 16195 37335 16201
rect 37366 16192 37372 16204
rect 37424 16192 37430 16244
rect 39942 16192 39948 16244
rect 40000 16232 40006 16244
rect 40000 16204 40264 16232
rect 40000 16192 40006 16204
rect 37090 16164 37096 16176
rect 37003 16136 37096 16164
rect 35161 16031 35219 16037
rect 35161 15997 35173 16031
rect 35207 16028 35219 16031
rect 35342 16028 35348 16040
rect 35207 16000 35348 16028
rect 35207 15997 35219 16000
rect 35161 15991 35219 15997
rect 35342 15988 35348 16000
rect 35400 15988 35406 16040
rect 35437 16031 35495 16037
rect 35437 15997 35449 16031
rect 35483 16028 35495 16031
rect 37016 16028 37044 16136
rect 37090 16124 37096 16136
rect 37148 16164 37154 16176
rect 37645 16167 37703 16173
rect 37645 16164 37657 16167
rect 37148 16136 37657 16164
rect 37148 16124 37154 16136
rect 37645 16133 37657 16136
rect 37691 16133 37703 16167
rect 37645 16127 37703 16133
rect 37182 16056 37188 16108
rect 37240 16096 37246 16108
rect 37461 16099 37519 16105
rect 37461 16096 37473 16099
rect 37240 16068 37473 16096
rect 37240 16056 37246 16068
rect 37461 16065 37473 16068
rect 37507 16065 37519 16099
rect 37461 16059 37519 16065
rect 37553 16099 37611 16105
rect 37553 16065 37565 16099
rect 37599 16065 37611 16099
rect 37553 16059 37611 16065
rect 37829 16099 37887 16105
rect 37829 16065 37841 16099
rect 37875 16096 37887 16099
rect 38654 16096 38660 16108
rect 37875 16068 38660 16096
rect 37875 16065 37887 16068
rect 37829 16059 37887 16065
rect 35483 16000 37044 16028
rect 37568 16028 37596 16059
rect 38654 16056 38660 16068
rect 38712 16056 38718 16108
rect 39965 16099 40023 16105
rect 39965 16065 39977 16099
rect 40011 16096 40023 16099
rect 40126 16096 40132 16108
rect 40011 16068 40132 16096
rect 40011 16065 40023 16068
rect 39965 16059 40023 16065
rect 40126 16056 40132 16068
rect 40184 16056 40190 16108
rect 40236 16105 40264 16204
rect 40221 16099 40279 16105
rect 40221 16065 40233 16099
rect 40267 16065 40279 16099
rect 40221 16059 40279 16065
rect 37568 16000 38884 16028
rect 35483 15997 35495 16000
rect 35437 15991 35495 15997
rect 38289 15963 38347 15969
rect 38289 15960 38301 15963
rect 35084 15932 38301 15960
rect 38289 15929 38301 15932
rect 38335 15960 38347 15963
rect 38746 15960 38752 15972
rect 38335 15932 38752 15960
rect 38335 15929 38347 15932
rect 38289 15923 38347 15929
rect 38746 15920 38752 15932
rect 38804 15920 38810 15972
rect 36906 15892 36912 15904
rect 32640 15864 36912 15892
rect 32640 15852 32646 15864
rect 36906 15852 36912 15864
rect 36964 15852 36970 15904
rect 38856 15901 38884 16000
rect 38841 15895 38899 15901
rect 38841 15861 38853 15895
rect 38887 15892 38899 15895
rect 38930 15892 38936 15904
rect 38887 15864 38936 15892
rect 38887 15861 38899 15864
rect 38841 15855 38899 15861
rect 38930 15852 38936 15864
rect 38988 15852 38994 15904
rect 58158 15892 58164 15904
rect 58119 15864 58164 15892
rect 58158 15852 58164 15864
rect 58216 15852 58222 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2498 15688 2504 15700
rect 2459 15660 2504 15688
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 6822 15688 6828 15700
rect 6783 15660 6828 15688
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 7745 15691 7803 15697
rect 7745 15657 7757 15691
rect 7791 15688 7803 15691
rect 7834 15688 7840 15700
rect 7791 15660 7840 15688
rect 7791 15657 7803 15660
rect 7745 15651 7803 15657
rect 7834 15648 7840 15660
rect 7892 15648 7898 15700
rect 9306 15688 9312 15700
rect 9267 15660 9312 15688
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 11974 15688 11980 15700
rect 10152 15660 11980 15688
rect 6454 15580 6460 15632
rect 6512 15620 6518 15632
rect 7377 15623 7435 15629
rect 7377 15620 7389 15623
rect 6512 15592 7389 15620
rect 6512 15580 6518 15592
rect 7377 15589 7389 15592
rect 7423 15589 7435 15623
rect 7377 15583 7435 15589
rect 9953 15623 10011 15629
rect 9953 15589 9965 15623
rect 9999 15589 10011 15623
rect 9953 15583 10011 15589
rect 6825 15555 6883 15561
rect 6825 15521 6837 15555
rect 6871 15552 6883 15555
rect 7098 15552 7104 15564
rect 6871 15524 7104 15552
rect 6871 15521 6883 15524
rect 6825 15515 6883 15521
rect 7098 15512 7104 15524
rect 7156 15552 7162 15564
rect 7558 15552 7564 15564
rect 7156 15524 7564 15552
rect 7156 15512 7162 15524
rect 7558 15512 7564 15524
rect 7616 15512 7622 15564
rect 9968 15552 9996 15583
rect 7760 15524 9996 15552
rect 2222 15484 2228 15496
rect 2183 15456 2228 15484
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15484 2375 15487
rect 3878 15484 3884 15496
rect 2363 15456 3884 15484
rect 2363 15453 2375 15456
rect 2317 15447 2375 15453
rect 3878 15444 3884 15456
rect 3936 15444 3942 15496
rect 6917 15487 6975 15493
rect 6917 15453 6929 15487
rect 6963 15453 6975 15487
rect 7650 15484 7656 15496
rect 7611 15456 7656 15484
rect 6917 15447 6975 15453
rect 5074 15376 5080 15428
rect 5132 15416 5138 15428
rect 6730 15416 6736 15428
rect 5132 15388 6736 15416
rect 5132 15376 5138 15388
rect 6730 15376 6736 15388
rect 6788 15376 6794 15428
rect 6932 15416 6960 15447
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 7760 15493 7788 15524
rect 7745 15487 7803 15493
rect 7745 15453 7757 15487
rect 7791 15453 7803 15487
rect 9398 15484 9404 15496
rect 9359 15456 9404 15484
rect 7745 15447 7803 15453
rect 9398 15444 9404 15456
rect 9456 15444 9462 15496
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15484 9551 15487
rect 9674 15484 9680 15496
rect 9539 15456 9680 15484
rect 9539 15453 9551 15456
rect 9493 15447 9551 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 10152 15493 10180 15660
rect 11974 15648 11980 15660
rect 12032 15648 12038 15700
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 14274 15688 14280 15700
rect 12492 15660 12537 15688
rect 14235 15660 14280 15688
rect 12492 15648 12498 15660
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 21269 15691 21327 15697
rect 21269 15657 21281 15691
rect 21315 15688 21327 15691
rect 21542 15688 21548 15700
rect 21315 15660 21548 15688
rect 21315 15657 21327 15660
rect 21269 15651 21327 15657
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 22465 15691 22523 15697
rect 22465 15657 22477 15691
rect 22511 15688 22523 15691
rect 22554 15688 22560 15700
rect 22511 15660 22560 15688
rect 22511 15657 22523 15660
rect 22465 15651 22523 15657
rect 22554 15648 22560 15660
rect 22612 15648 22618 15700
rect 23293 15691 23351 15697
rect 23293 15657 23305 15691
rect 23339 15688 23351 15691
rect 23474 15688 23480 15700
rect 23339 15660 23480 15688
rect 23339 15657 23351 15660
rect 23293 15651 23351 15657
rect 23474 15648 23480 15660
rect 23532 15648 23538 15700
rect 27062 15688 27068 15700
rect 27023 15660 27068 15688
rect 27062 15648 27068 15660
rect 27120 15648 27126 15700
rect 29546 15688 29552 15700
rect 29507 15660 29552 15688
rect 29546 15648 29552 15660
rect 29604 15648 29610 15700
rect 30650 15648 30656 15700
rect 30708 15688 30714 15700
rect 32582 15688 32588 15700
rect 30708 15660 31754 15688
rect 32543 15660 32588 15688
rect 30708 15648 30714 15660
rect 10870 15552 10876 15564
rect 10244 15524 10876 15552
rect 10244 15493 10272 15524
rect 10870 15512 10876 15524
rect 10928 15512 10934 15564
rect 11054 15552 11060 15564
rect 11015 15524 11060 15552
rect 11054 15512 11060 15524
rect 11112 15512 11118 15564
rect 12452 15552 12480 15648
rect 30926 15580 30932 15632
rect 30984 15580 30990 15632
rect 14550 15552 14556 15564
rect 12452 15524 13032 15552
rect 10132 15487 10190 15493
rect 10132 15453 10144 15487
rect 10178 15453 10190 15487
rect 10132 15447 10190 15453
rect 10229 15487 10287 15493
rect 10229 15453 10241 15487
rect 10275 15453 10287 15487
rect 10502 15484 10508 15496
rect 10463 15456 10508 15484
rect 10229 15447 10287 15453
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 10594 15444 10600 15496
rect 10652 15484 10658 15496
rect 11324 15487 11382 15493
rect 10652 15456 10697 15484
rect 10652 15444 10658 15456
rect 11324 15453 11336 15487
rect 11370 15484 11382 15487
rect 11882 15484 11888 15496
rect 11370 15456 11888 15484
rect 11370 15453 11382 15456
rect 11324 15447 11382 15453
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 12894 15484 12900 15496
rect 12855 15456 12900 15484
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 13004 15493 13032 15524
rect 13188 15524 14556 15552
rect 13188 15493 13216 15524
rect 14550 15512 14556 15524
rect 14608 15512 14614 15564
rect 19242 15552 19248 15564
rect 19203 15524 19248 15552
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 20990 15512 20996 15564
rect 21048 15552 21054 15564
rect 23753 15555 23811 15561
rect 23753 15552 23765 15555
rect 21048 15524 23765 15552
rect 21048 15512 21054 15524
rect 12990 15487 13048 15493
rect 12990 15453 13002 15487
rect 13036 15453 13048 15487
rect 12990 15447 13048 15453
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15453 13231 15487
rect 13173 15447 13231 15453
rect 13403 15487 13461 15493
rect 13403 15453 13415 15487
rect 13449 15484 13461 15487
rect 13814 15484 13820 15496
rect 13449 15456 13820 15484
rect 13449 15453 13461 15456
rect 13403 15447 13461 15453
rect 10321 15419 10379 15425
rect 6932 15388 9260 15416
rect 6546 15348 6552 15360
rect 6507 15320 6552 15348
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 8386 15308 8392 15360
rect 8444 15348 8450 15360
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 8444 15320 9137 15348
rect 8444 15308 8450 15320
rect 9125 15317 9137 15320
rect 9171 15317 9183 15351
rect 9232 15348 9260 15388
rect 10321 15385 10333 15419
rect 10367 15416 10379 15419
rect 11790 15416 11796 15428
rect 10367 15388 11796 15416
rect 10367 15385 10379 15388
rect 10321 15379 10379 15385
rect 11790 15376 11796 15388
rect 11848 15416 11854 15428
rect 13188 15416 13216 15447
rect 13814 15444 13820 15456
rect 13872 15444 13878 15496
rect 14093 15487 14151 15493
rect 14093 15453 14105 15487
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 11848 15388 13216 15416
rect 11848 15376 11854 15388
rect 13262 15376 13268 15428
rect 13320 15416 13326 15428
rect 14108 15416 14136 15447
rect 14182 15444 14188 15496
rect 14240 15484 14246 15496
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 14240 15456 14289 15484
rect 14240 15444 14246 15456
rect 14277 15453 14289 15456
rect 14323 15453 14335 15487
rect 15102 15484 15108 15496
rect 15063 15456 15108 15484
rect 14277 15447 14335 15453
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15378 15493 15384 15496
rect 15372 15484 15384 15493
rect 15339 15456 15384 15484
rect 15372 15447 15384 15456
rect 15378 15444 15384 15447
rect 15436 15444 15442 15496
rect 18690 15444 18696 15496
rect 18748 15484 18754 15496
rect 19501 15487 19559 15493
rect 19501 15484 19513 15487
rect 18748 15456 19513 15484
rect 18748 15444 18754 15456
rect 19501 15453 19513 15456
rect 19547 15453 19559 15487
rect 19501 15447 19559 15453
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15453 21143 15487
rect 21266 15484 21272 15496
rect 21227 15456 21272 15484
rect 21085 15447 21143 15453
rect 14366 15416 14372 15428
rect 13320 15388 13365 15416
rect 14108 15388 14372 15416
rect 13320 15376 13326 15388
rect 14366 15376 14372 15388
rect 14424 15376 14430 15428
rect 21100 15416 21128 15447
rect 21266 15444 21272 15456
rect 21324 15444 21330 15496
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 23124 15493 23152 15524
rect 23753 15521 23765 15524
rect 23799 15521 23811 15555
rect 23753 15515 23811 15521
rect 22465 15487 22523 15493
rect 22465 15484 22477 15487
rect 22152 15456 22477 15484
rect 22152 15444 22158 15456
rect 22465 15453 22477 15456
rect 22511 15453 22523 15487
rect 22465 15447 22523 15453
rect 22649 15487 22707 15493
rect 22649 15453 22661 15487
rect 22695 15453 22707 15487
rect 22649 15447 22707 15453
rect 23109 15487 23167 15493
rect 23109 15453 23121 15487
rect 23155 15453 23167 15487
rect 23290 15484 23296 15496
rect 23109 15447 23167 15453
rect 23216 15456 23296 15484
rect 21174 15416 21180 15428
rect 21100 15388 21180 15416
rect 21174 15376 21180 15388
rect 21232 15376 21238 15428
rect 22186 15376 22192 15428
rect 22244 15416 22250 15428
rect 22664 15416 22692 15447
rect 23216 15416 23244 15456
rect 23290 15444 23296 15456
rect 23348 15484 23354 15496
rect 24397 15487 24455 15493
rect 24397 15484 24409 15487
rect 23348 15456 24409 15484
rect 23348 15444 23354 15456
rect 24397 15453 24409 15456
rect 24443 15453 24455 15487
rect 26970 15484 26976 15496
rect 26931 15456 26976 15484
rect 24397 15447 24455 15453
rect 26970 15444 26976 15456
rect 27028 15444 27034 15496
rect 27154 15484 27160 15496
rect 27115 15456 27160 15484
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 30944 15493 30972 15580
rect 31726 15552 31754 15660
rect 32582 15648 32588 15660
rect 32640 15648 32646 15700
rect 36906 15688 36912 15700
rect 36867 15660 36912 15688
rect 36906 15648 36912 15660
rect 36964 15648 36970 15700
rect 40126 15648 40132 15700
rect 40184 15688 40190 15700
rect 41785 15691 41843 15697
rect 41785 15688 41797 15691
rect 40184 15660 41797 15688
rect 40184 15648 40190 15660
rect 41785 15657 41797 15660
rect 41831 15657 41843 15691
rect 41785 15651 41843 15657
rect 39574 15580 39580 15632
rect 39632 15620 39638 15632
rect 40494 15620 40500 15632
rect 39632 15592 40500 15620
rect 39632 15580 39638 15592
rect 40494 15580 40500 15592
rect 40552 15620 40558 15632
rect 40552 15592 41460 15620
rect 40552 15580 40558 15592
rect 35713 15555 35771 15561
rect 31726 15524 31800 15552
rect 30929 15487 30987 15493
rect 30929 15453 30941 15487
rect 30975 15453 30987 15487
rect 30929 15447 30987 15453
rect 31018 15444 31024 15496
rect 31076 15484 31082 15496
rect 31772 15493 31800 15524
rect 35713 15521 35725 15555
rect 35759 15552 35771 15555
rect 37182 15552 37188 15564
rect 35759 15524 37188 15552
rect 35759 15521 35771 15524
rect 35713 15515 35771 15521
rect 37182 15512 37188 15524
rect 37240 15512 37246 15564
rect 37826 15512 37832 15564
rect 37884 15552 37890 15564
rect 40405 15555 40463 15561
rect 37884 15524 38516 15552
rect 37884 15512 37890 15524
rect 31665 15487 31723 15493
rect 31665 15484 31677 15487
rect 31076 15456 31677 15484
rect 31076 15444 31082 15456
rect 31665 15453 31677 15456
rect 31711 15453 31723 15487
rect 31665 15447 31723 15453
rect 31757 15487 31815 15493
rect 31757 15453 31769 15487
rect 31803 15453 31815 15487
rect 31757 15447 31815 15453
rect 31849 15487 31907 15493
rect 31849 15453 31861 15487
rect 31895 15453 31907 15487
rect 32030 15484 32036 15496
rect 31991 15456 32036 15484
rect 31849 15447 31907 15453
rect 22244 15388 22692 15416
rect 22756 15388 23244 15416
rect 26988 15416 27016 15444
rect 27617 15419 27675 15425
rect 27617 15416 27629 15419
rect 26988 15388 27629 15416
rect 22244 15376 22250 15388
rect 22756 15360 22784 15388
rect 27617 15385 27629 15388
rect 27663 15385 27675 15419
rect 27617 15379 27675 15385
rect 30684 15419 30742 15425
rect 30684 15385 30696 15419
rect 30730 15416 30742 15419
rect 31389 15419 31447 15425
rect 31389 15416 31401 15419
rect 30730 15388 31401 15416
rect 30730 15385 30742 15388
rect 30684 15379 30742 15385
rect 31389 15385 31401 15388
rect 31435 15385 31447 15419
rect 31389 15379 31447 15385
rect 31478 15376 31484 15428
rect 31536 15416 31542 15428
rect 31864 15416 31892 15447
rect 32030 15444 32036 15456
rect 32088 15444 32094 15496
rect 33226 15444 33232 15496
rect 33284 15484 33290 15496
rect 33321 15487 33379 15493
rect 33321 15484 33333 15487
rect 33284 15456 33333 15484
rect 33284 15444 33290 15456
rect 33321 15453 33333 15456
rect 33367 15453 33379 15487
rect 33594 15484 33600 15496
rect 33555 15456 33600 15484
rect 33321 15447 33379 15453
rect 33594 15444 33600 15456
rect 33652 15444 33658 15496
rect 34698 15444 34704 15496
rect 34756 15484 34762 15496
rect 35437 15487 35495 15493
rect 35437 15484 35449 15487
rect 34756 15456 35449 15484
rect 34756 15444 34762 15456
rect 35437 15453 35449 15456
rect 35483 15453 35495 15487
rect 35437 15447 35495 15453
rect 37369 15487 37427 15493
rect 37369 15453 37381 15487
rect 37415 15484 37427 15487
rect 37642 15484 37648 15496
rect 37415 15456 37648 15484
rect 37415 15453 37427 15456
rect 37369 15447 37427 15453
rect 37642 15444 37648 15456
rect 37700 15444 37706 15496
rect 38194 15484 38200 15496
rect 38155 15456 38200 15484
rect 38194 15444 38200 15456
rect 38252 15444 38258 15496
rect 38488 15493 38516 15524
rect 40405 15521 40417 15555
rect 40451 15552 40463 15555
rect 40451 15524 41184 15552
rect 40451 15521 40463 15524
rect 40405 15515 40463 15521
rect 41156 15496 41184 15524
rect 38360 15484 38418 15490
rect 38360 15481 38372 15484
rect 38304 15453 38372 15481
rect 31536 15388 31892 15416
rect 37553 15419 37611 15425
rect 31536 15376 31542 15388
rect 37553 15385 37565 15419
rect 37599 15385 37611 15419
rect 37553 15379 37611 15385
rect 37737 15419 37795 15425
rect 37737 15385 37749 15419
rect 37783 15416 37795 15419
rect 38304 15416 38332 15453
rect 38360 15450 38372 15453
rect 38406 15450 38418 15484
rect 38360 15444 38418 15450
rect 38473 15487 38531 15493
rect 38473 15453 38485 15487
rect 38519 15453 38531 15487
rect 38473 15447 38531 15453
rect 38611 15487 38669 15493
rect 38611 15453 38623 15487
rect 38657 15484 38669 15487
rect 38746 15484 38752 15496
rect 38657 15456 38752 15484
rect 38657 15453 38669 15456
rect 38611 15447 38669 15453
rect 38746 15444 38752 15456
rect 38804 15444 38810 15496
rect 40678 15484 40684 15496
rect 40639 15456 40684 15484
rect 40678 15444 40684 15456
rect 40736 15444 40742 15496
rect 41138 15484 41144 15496
rect 41099 15456 41144 15484
rect 41138 15444 41144 15456
rect 41196 15444 41202 15496
rect 41322 15484 41328 15496
rect 41283 15456 41328 15484
rect 41322 15444 41328 15456
rect 41380 15444 41386 15496
rect 41432 15493 41460 15592
rect 41417 15487 41475 15493
rect 41417 15453 41429 15487
rect 41463 15453 41475 15487
rect 41417 15447 41475 15453
rect 41506 15444 41512 15496
rect 41564 15484 41570 15496
rect 41564 15456 41609 15484
rect 41564 15444 41570 15456
rect 37783 15388 38332 15416
rect 37783 15385 37795 15388
rect 37737 15379 37795 15385
rect 13541 15351 13599 15357
rect 13541 15348 13553 15351
rect 9232 15320 13553 15348
rect 9125 15311 9183 15317
rect 13541 15317 13553 15320
rect 13587 15317 13599 15351
rect 13541 15311 13599 15317
rect 16485 15351 16543 15357
rect 16485 15317 16497 15351
rect 16531 15348 16543 15351
rect 16942 15348 16948 15360
rect 16531 15320 16948 15348
rect 16531 15317 16543 15320
rect 16485 15311 16543 15317
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 18417 15351 18475 15357
rect 18417 15317 18429 15351
rect 18463 15348 18475 15351
rect 18782 15348 18788 15360
rect 18463 15320 18788 15348
rect 18463 15317 18475 15320
rect 18417 15311 18475 15317
rect 18782 15308 18788 15320
rect 18840 15308 18846 15360
rect 20622 15348 20628 15360
rect 20583 15320 20628 15348
rect 20622 15308 20628 15320
rect 20680 15308 20686 15360
rect 21910 15348 21916 15360
rect 21871 15320 21916 15348
rect 21910 15308 21916 15320
rect 21968 15348 21974 15360
rect 22738 15348 22744 15360
rect 21968 15320 22744 15348
rect 21968 15308 21974 15320
rect 22738 15308 22744 15320
rect 22796 15308 22802 15360
rect 37568 15348 37596 15379
rect 38654 15348 38660 15360
rect 37568 15320 38660 15348
rect 38654 15308 38660 15320
rect 38712 15308 38718 15360
rect 38838 15348 38844 15360
rect 38799 15320 38844 15348
rect 38838 15308 38844 15320
rect 38896 15308 38902 15360
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 7742 15144 7748 15156
rect 7655 15116 7748 15144
rect 7742 15104 7748 15116
rect 7800 15144 7806 15156
rect 7800 15116 9812 15144
rect 7800 15104 7806 15116
rect 6730 15036 6736 15088
rect 6788 15076 6794 15088
rect 8880 15079 8938 15085
rect 6788 15048 6960 15076
rect 6788 15036 6794 15048
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 2866 14968 2872 15020
rect 2924 15008 2930 15020
rect 3033 15011 3091 15017
rect 3033 15008 3045 15011
rect 2924 14980 3045 15008
rect 2924 14968 2930 14980
rect 3033 14977 3045 14980
rect 3079 14977 3091 15011
rect 5626 15008 5632 15020
rect 5587 14980 5632 15008
rect 3033 14971 3091 14977
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 6362 15008 6368 15020
rect 6323 14980 6368 15008
rect 6362 14968 6368 14980
rect 6420 14968 6426 15020
rect 6546 15008 6552 15020
rect 6507 14980 6552 15008
rect 6546 14968 6552 14980
rect 6604 14968 6610 15020
rect 6638 14968 6644 15020
rect 6696 15008 6702 15020
rect 6932 15017 6960 15048
rect 8880 15045 8892 15079
rect 8926 15076 8938 15079
rect 9585 15079 9643 15085
rect 9585 15076 9597 15079
rect 8926 15048 9597 15076
rect 8926 15045 8938 15048
rect 8880 15039 8938 15045
rect 9585 15045 9597 15048
rect 9631 15045 9643 15079
rect 9585 15039 9643 15045
rect 6917 15011 6975 15017
rect 6696 14980 6741 15008
rect 6696 14968 6702 14980
rect 6917 14977 6929 15011
rect 6963 14977 6975 15011
rect 9122 15008 9128 15020
rect 9083 14980 9128 15008
rect 6917 14971 6975 14977
rect 9122 14968 9128 14980
rect 9180 14968 9186 15020
rect 9784 15017 9812 15116
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 13078 15144 13084 15156
rect 12860 15116 13084 15144
rect 12860 15104 12866 15116
rect 13078 15104 13084 15116
rect 13136 15144 13142 15156
rect 13136 15116 17356 15144
rect 13136 15104 13142 15116
rect 14277 15079 14335 15085
rect 14277 15045 14289 15079
rect 14323 15076 14335 15079
rect 16666 15076 16672 15088
rect 14323 15048 16672 15076
rect 14323 15045 14335 15048
rect 14277 15039 14335 15045
rect 16666 15036 16672 15048
rect 16724 15036 16730 15088
rect 17120 15079 17178 15085
rect 17120 15045 17132 15079
rect 17166 15076 17178 15079
rect 17218 15076 17224 15088
rect 17166 15048 17224 15076
rect 17166 15045 17178 15048
rect 17120 15039 17178 15045
rect 17218 15036 17224 15048
rect 17276 15036 17282 15088
rect 17328 15076 17356 15116
rect 18506 15104 18512 15156
rect 18564 15144 18570 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 18564 15116 18797 15144
rect 18564 15104 18570 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 24210 15144 24216 15156
rect 24171 15116 24216 15144
rect 18785 15107 18843 15113
rect 24210 15104 24216 15116
rect 24268 15104 24274 15156
rect 25038 15144 25044 15156
rect 24999 15116 25044 15144
rect 25038 15104 25044 15116
rect 25096 15104 25102 15156
rect 25590 15104 25596 15156
rect 25648 15144 25654 15156
rect 27614 15144 27620 15156
rect 25648 15116 27620 15144
rect 25648 15104 25654 15116
rect 27614 15104 27620 15116
rect 27672 15104 27678 15156
rect 28258 15144 28264 15156
rect 28219 15116 28264 15144
rect 28258 15104 28264 15116
rect 28316 15104 28322 15156
rect 29917 15147 29975 15153
rect 29917 15113 29929 15147
rect 29963 15144 29975 15147
rect 30558 15144 30564 15156
rect 29963 15116 30564 15144
rect 29963 15113 29975 15116
rect 29917 15107 29975 15113
rect 30558 15104 30564 15116
rect 30616 15104 30622 15156
rect 37461 15147 37519 15153
rect 37461 15113 37473 15147
rect 37507 15144 37519 15147
rect 37826 15144 37832 15156
rect 37507 15116 37832 15144
rect 37507 15113 37519 15116
rect 37461 15107 37519 15113
rect 37826 15104 37832 15116
rect 37884 15144 37890 15156
rect 38562 15144 38568 15156
rect 37884 15116 38568 15144
rect 37884 15104 37890 15116
rect 38562 15104 38568 15116
rect 38620 15104 38626 15156
rect 38654 15104 38660 15156
rect 38712 15144 38718 15156
rect 40221 15147 40279 15153
rect 40221 15144 40233 15147
rect 38712 15116 40233 15144
rect 38712 15104 38718 15116
rect 40221 15113 40233 15116
rect 40267 15113 40279 15147
rect 40221 15107 40279 15113
rect 19429 15079 19487 15085
rect 19429 15076 19441 15079
rect 17328 15048 19441 15076
rect 9769 15011 9827 15017
rect 9769 14977 9781 15011
rect 9815 14977 9827 15011
rect 10134 15008 10140 15020
rect 10095 14980 10140 15008
rect 9769 14971 9827 14977
rect 10134 14968 10140 14980
rect 10192 14968 10198 15020
rect 10321 15011 10379 15017
rect 10321 14977 10333 15011
rect 10367 15008 10379 15011
rect 11054 15008 11060 15020
rect 10367 14980 11060 15008
rect 10367 14977 10379 14980
rect 10321 14971 10379 14977
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 18708 15017 18736 15048
rect 19429 15045 19441 15048
rect 19475 15076 19487 15079
rect 22094 15076 22100 15088
rect 19475 15048 22100 15076
rect 19475 15045 19487 15048
rect 19429 15039 19487 15045
rect 22094 15036 22100 15048
rect 22152 15076 22158 15088
rect 22649 15079 22707 15085
rect 22152 15048 22600 15076
rect 22152 15036 22158 15048
rect 14093 15011 14151 15017
rect 14093 15008 14105 15011
rect 12032 14980 14105 15008
rect 12032 14968 12038 14980
rect 14093 14977 14105 14980
rect 14139 14977 14151 15011
rect 14093 14971 14151 14977
rect 18693 15011 18751 15017
rect 18693 14977 18705 15011
rect 18739 14977 18751 15011
rect 18693 14971 18751 14977
rect 18782 14968 18788 15020
rect 18840 15008 18846 15020
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 18840 14980 18889 15008
rect 18840 14968 18846 14980
rect 18877 14977 18889 14980
rect 18923 14977 18935 15011
rect 18877 14971 18935 14977
rect 20070 14968 20076 15020
rect 20128 15008 20134 15020
rect 22572 15017 22600 15048
rect 22649 15045 22661 15079
rect 22695 15076 22707 15079
rect 22695 15048 32720 15076
rect 22695 15045 22707 15048
rect 22649 15039 22707 15045
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 20128 14980 20453 15008
rect 20128 14968 20134 14980
rect 20441 14977 20453 14980
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 22557 15011 22615 15017
rect 22557 14977 22569 15011
rect 22603 14977 22615 15011
rect 22738 15008 22744 15020
rect 22699 14980 22744 15008
rect 22557 14971 22615 14977
rect 22738 14968 22744 14980
rect 22796 14968 22802 15020
rect 23201 15011 23259 15017
rect 23201 14977 23213 15011
rect 23247 14977 23259 15011
rect 23201 14971 23259 14977
rect 1949 14943 2007 14949
rect 1949 14909 1961 14943
rect 1995 14940 2007 14943
rect 2222 14940 2228 14952
rect 1995 14912 2228 14940
rect 1995 14909 2007 14912
rect 1949 14903 2007 14909
rect 2222 14900 2228 14912
rect 2280 14940 2286 14952
rect 2682 14940 2688 14952
rect 2280 14912 2688 14940
rect 2280 14900 2286 14912
rect 2682 14900 2688 14912
rect 2740 14900 2746 14952
rect 2777 14943 2835 14949
rect 2777 14909 2789 14943
rect 2823 14909 2835 14943
rect 2777 14903 2835 14909
rect 5169 14943 5227 14949
rect 5169 14909 5181 14943
rect 5215 14940 5227 14943
rect 5258 14940 5264 14952
rect 5215 14912 5264 14940
rect 5215 14909 5227 14912
rect 5169 14903 5227 14909
rect 2317 14807 2375 14813
rect 2317 14773 2329 14807
rect 2363 14804 2375 14807
rect 2590 14804 2596 14816
rect 2363 14776 2596 14804
rect 2363 14773 2375 14776
rect 2317 14767 2375 14773
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 2792 14804 2820 14903
rect 5258 14900 5264 14912
rect 5316 14900 5322 14952
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14909 5595 14943
rect 5537 14903 5595 14909
rect 6733 14943 6791 14949
rect 6733 14909 6745 14943
rect 6779 14940 6791 14943
rect 7374 14940 7380 14952
rect 6779 14912 7380 14940
rect 6779 14909 6791 14912
rect 6733 14903 6791 14909
rect 3786 14804 3792 14816
rect 2792 14776 3792 14804
rect 3786 14764 3792 14776
rect 3844 14764 3850 14816
rect 4157 14807 4215 14813
rect 4157 14773 4169 14807
rect 4203 14804 4215 14807
rect 4982 14804 4988 14816
rect 4203 14776 4988 14804
rect 4203 14773 4215 14776
rect 4157 14767 4215 14773
rect 4982 14764 4988 14776
rect 5040 14804 5046 14816
rect 5552 14804 5580 14903
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14909 10011 14943
rect 9953 14903 10011 14909
rect 9766 14832 9772 14884
rect 9824 14872 9830 14884
rect 9968 14872 9996 14903
rect 10042 14900 10048 14952
rect 10100 14940 10106 14952
rect 10100 14912 10145 14940
rect 10100 14900 10106 14912
rect 15102 14900 15108 14952
rect 15160 14940 15166 14952
rect 16850 14940 16856 14952
rect 15160 14912 16856 14940
rect 15160 14900 15166 14912
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 20162 14940 20168 14952
rect 20123 14912 20168 14940
rect 20162 14900 20168 14912
rect 20220 14900 20226 14952
rect 22186 14900 22192 14952
rect 22244 14940 22250 14952
rect 23216 14940 23244 14971
rect 23290 14968 23296 15020
rect 23348 15008 23354 15020
rect 23385 15011 23443 15017
rect 23385 15008 23397 15011
rect 23348 14980 23397 15008
rect 23348 14968 23354 14980
rect 23385 14977 23397 14980
rect 23431 14977 23443 15011
rect 23385 14971 23443 14977
rect 24118 14968 24124 15020
rect 24176 15008 24182 15020
rect 27525 15011 27583 15017
rect 27525 15008 27537 15011
rect 24176 14980 27537 15008
rect 24176 14968 24182 14980
rect 27525 14977 27537 14980
rect 27571 15008 27583 15011
rect 27614 15008 27620 15020
rect 27571 14980 27620 15008
rect 27571 14977 27583 14980
rect 27525 14971 27583 14977
rect 27614 14968 27620 14980
rect 27672 14968 27678 15020
rect 27709 15011 27767 15017
rect 27709 14977 27721 15011
rect 27755 14977 27767 15011
rect 27709 14971 27767 14977
rect 22244 14912 23244 14940
rect 27724 14940 27752 14971
rect 29638 14968 29644 15020
rect 29696 15008 29702 15020
rect 30193 15011 30251 15017
rect 30193 15008 30205 15011
rect 29696 14980 30205 15008
rect 29696 14968 29702 14980
rect 30193 14977 30205 14980
rect 30239 14977 30251 15011
rect 30193 14971 30251 14977
rect 30285 15011 30343 15017
rect 30285 14977 30297 15011
rect 30331 14977 30343 15011
rect 30285 14971 30343 14977
rect 29822 14940 29828 14952
rect 27724 14912 29828 14940
rect 22244 14900 22250 14912
rect 29822 14900 29828 14912
rect 29880 14900 29886 14952
rect 29914 14900 29920 14952
rect 29972 14940 29978 14952
rect 30300 14940 30328 14971
rect 30374 14968 30380 15020
rect 30432 15008 30438 15020
rect 30432 14980 30477 15008
rect 30432 14968 30438 14980
rect 30558 14968 30564 15020
rect 30616 15008 30622 15020
rect 32030 15008 32036 15020
rect 30616 14980 32036 15008
rect 30616 14968 30622 14980
rect 32030 14968 32036 14980
rect 32088 14968 32094 15020
rect 32692 15008 32720 15048
rect 38838 15036 38844 15088
rect 38896 15076 38902 15088
rect 39086 15079 39144 15085
rect 39086 15076 39098 15079
rect 38896 15048 39098 15076
rect 38896 15036 38902 15048
rect 39086 15045 39098 15048
rect 39132 15045 39144 15079
rect 39086 15039 39144 15045
rect 35342 15008 35348 15020
rect 32692 14980 35348 15008
rect 35268 14978 35348 14980
rect 35342 14968 35348 14978
rect 35400 14968 35406 15020
rect 35710 14968 35716 15020
rect 35768 15008 35774 15020
rect 35989 15011 36047 15017
rect 35989 15008 36001 15011
rect 35768 14980 36001 15008
rect 35768 14968 35774 14980
rect 35989 14977 36001 14980
rect 36035 14977 36047 15011
rect 35989 14971 36047 14977
rect 37277 15011 37335 15017
rect 37277 14977 37289 15011
rect 37323 14977 37335 15011
rect 37277 14971 37335 14977
rect 29972 14912 30328 14940
rect 35069 14943 35127 14949
rect 29972 14900 29978 14912
rect 35069 14909 35081 14943
rect 35115 14940 35127 14943
rect 35618 14940 35624 14952
rect 35115 14912 35624 14940
rect 35115 14909 35127 14912
rect 35069 14903 35127 14909
rect 35618 14900 35624 14912
rect 35676 14900 35682 14952
rect 35802 14940 35808 14952
rect 35763 14912 35808 14940
rect 35802 14900 35808 14912
rect 35860 14940 35866 14952
rect 36633 14943 36691 14949
rect 36633 14940 36645 14943
rect 35860 14912 36645 14940
rect 35860 14900 35866 14912
rect 36633 14909 36645 14912
rect 36679 14909 36691 14943
rect 36633 14903 36691 14909
rect 9824 14844 9996 14872
rect 9824 14832 9830 14844
rect 13814 14832 13820 14884
rect 13872 14872 13878 14884
rect 18230 14872 18236 14884
rect 13872 14844 14872 14872
rect 18143 14844 18236 14872
rect 13872 14832 13878 14844
rect 5810 14804 5816 14816
rect 5040 14776 5580 14804
rect 5771 14776 5816 14804
rect 5040 14764 5046 14776
rect 5810 14764 5816 14776
rect 5868 14764 5874 14816
rect 7098 14804 7104 14816
rect 7059 14776 7104 14804
rect 7098 14764 7104 14776
rect 7156 14764 7162 14816
rect 14366 14764 14372 14816
rect 14424 14804 14430 14816
rect 14737 14807 14795 14813
rect 14737 14804 14749 14807
rect 14424 14776 14749 14804
rect 14424 14764 14430 14776
rect 14737 14773 14749 14776
rect 14783 14773 14795 14807
rect 14844 14804 14872 14844
rect 18230 14832 18236 14844
rect 18288 14872 18294 14884
rect 22830 14872 22836 14884
rect 18288 14844 22836 14872
rect 18288 14832 18294 14844
rect 22830 14832 22836 14844
rect 22888 14832 22894 14884
rect 23385 14875 23443 14881
rect 23385 14841 23397 14875
rect 23431 14872 23443 14875
rect 34698 14872 34704 14884
rect 23431 14844 34704 14872
rect 23431 14841 23443 14844
rect 23385 14835 23443 14841
rect 34698 14832 34704 14844
rect 34756 14832 34762 14884
rect 35636 14872 35664 14900
rect 37292 14872 37320 14971
rect 37458 14968 37464 15020
rect 37516 15008 37522 15020
rect 37921 15011 37979 15017
rect 37921 15008 37933 15011
rect 37516 14980 37933 15008
rect 37516 14968 37522 14980
rect 37921 14977 37933 14980
rect 37967 14977 37979 15011
rect 37921 14971 37979 14977
rect 38746 14968 38752 15020
rect 38804 15008 38810 15020
rect 40957 15011 41015 15017
rect 40957 15008 40969 15011
rect 38804 14980 40969 15008
rect 38804 14968 38810 14980
rect 40957 14977 40969 14980
rect 41003 15008 41015 15011
rect 41506 15008 41512 15020
rect 41003 14980 41512 15008
rect 41003 14977 41015 14980
rect 40957 14971 41015 14977
rect 41506 14968 41512 14980
rect 41564 14968 41570 15020
rect 38102 14900 38108 14952
rect 38160 14940 38166 14952
rect 38841 14943 38899 14949
rect 38841 14940 38853 14943
rect 38160 14912 38853 14940
rect 38160 14900 38166 14912
rect 38841 14909 38853 14912
rect 38887 14909 38899 14943
rect 38841 14903 38899 14909
rect 35636 14844 37320 14872
rect 20346 14804 20352 14816
rect 14844 14776 20352 14804
rect 14737 14767 14795 14773
rect 20346 14764 20352 14776
rect 20404 14764 20410 14816
rect 20806 14764 20812 14816
rect 20864 14804 20870 14816
rect 20990 14804 20996 14816
rect 20864 14776 20996 14804
rect 20864 14764 20870 14776
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 22097 14807 22155 14813
rect 22097 14773 22109 14807
rect 22143 14804 22155 14807
rect 22186 14804 22192 14816
rect 22143 14776 22192 14804
rect 22143 14773 22155 14776
rect 22097 14767 22155 14773
rect 22186 14764 22192 14776
rect 22244 14764 22250 14816
rect 23474 14764 23480 14816
rect 23532 14804 23538 14816
rect 26970 14804 26976 14816
rect 23532 14776 26976 14804
rect 23532 14764 23538 14776
rect 26970 14764 26976 14776
rect 27028 14764 27034 14816
rect 27341 14807 27399 14813
rect 27341 14773 27353 14807
rect 27387 14804 27399 14807
rect 27706 14804 27712 14816
rect 27387 14776 27712 14804
rect 27387 14773 27399 14776
rect 27341 14767 27399 14773
rect 27706 14764 27712 14776
rect 27764 14764 27770 14816
rect 29457 14807 29515 14813
rect 29457 14773 29469 14807
rect 29503 14804 29515 14807
rect 29638 14804 29644 14816
rect 29503 14776 29644 14804
rect 29503 14773 29515 14776
rect 29457 14767 29515 14773
rect 29638 14764 29644 14776
rect 29696 14764 29702 14816
rect 31018 14764 31024 14816
rect 31076 14804 31082 14816
rect 31205 14807 31263 14813
rect 31205 14804 31217 14807
rect 31076 14776 31217 14804
rect 31076 14764 31082 14776
rect 31205 14773 31217 14776
rect 31251 14773 31263 14807
rect 33226 14804 33232 14816
rect 33187 14776 33232 14804
rect 31205 14767 31263 14773
rect 33226 14764 33232 14776
rect 33284 14764 33290 14816
rect 36173 14807 36231 14813
rect 36173 14773 36185 14807
rect 36219 14804 36231 14807
rect 36722 14804 36728 14816
rect 36219 14776 36728 14804
rect 36219 14773 36231 14776
rect 36173 14767 36231 14773
rect 36722 14764 36728 14776
rect 36780 14764 36786 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14600 2835 14603
rect 2866 14600 2872 14612
rect 2823 14572 2872 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 2866 14560 2872 14572
rect 2924 14560 2930 14612
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 10042 14600 10048 14612
rect 5868 14572 10048 14600
rect 5868 14560 5874 14572
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 10226 14560 10232 14612
rect 10284 14600 10290 14612
rect 10413 14603 10471 14609
rect 10413 14600 10425 14603
rect 10284 14572 10425 14600
rect 10284 14560 10290 14572
rect 10413 14569 10425 14572
rect 10459 14569 10471 14603
rect 10413 14563 10471 14569
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 16669 14603 16727 14609
rect 16669 14600 16681 14603
rect 16632 14572 16681 14600
rect 16632 14560 16638 14572
rect 16669 14569 16681 14572
rect 16715 14569 16727 14603
rect 18601 14603 18659 14609
rect 18601 14600 18613 14603
rect 16669 14563 16727 14569
rect 16776 14572 18613 14600
rect 2130 14492 2136 14544
rect 2188 14532 2194 14544
rect 4525 14535 4583 14541
rect 4525 14532 4537 14535
rect 2188 14504 4537 14532
rect 2188 14492 2194 14504
rect 4525 14501 4537 14504
rect 4571 14501 4583 14535
rect 4525 14495 4583 14501
rect 4890 14492 4896 14544
rect 4948 14532 4954 14544
rect 6365 14535 6423 14541
rect 6365 14532 6377 14535
rect 4948 14504 6377 14532
rect 4948 14492 4954 14504
rect 6365 14501 6377 14504
rect 6411 14532 6423 14535
rect 6730 14532 6736 14544
rect 6411 14504 6736 14532
rect 6411 14501 6423 14504
rect 6365 14495 6423 14501
rect 6730 14492 6736 14504
rect 6788 14492 6794 14544
rect 16776 14532 16804 14572
rect 18601 14569 18613 14572
rect 18647 14600 18659 14603
rect 18782 14600 18788 14612
rect 18647 14572 18788 14600
rect 18647 14569 18659 14572
rect 18601 14563 18659 14569
rect 18782 14560 18788 14572
rect 18840 14600 18846 14612
rect 19610 14600 19616 14612
rect 18840 14572 19616 14600
rect 18840 14560 18846 14572
rect 19610 14560 19616 14572
rect 19668 14600 19674 14612
rect 20806 14600 20812 14612
rect 19668 14572 20812 14600
rect 19668 14560 19674 14572
rect 20806 14560 20812 14572
rect 20864 14560 20870 14612
rect 20901 14603 20959 14609
rect 20901 14569 20913 14603
rect 20947 14600 20959 14603
rect 20990 14600 20996 14612
rect 20947 14572 20996 14600
rect 20947 14569 20959 14572
rect 20901 14563 20959 14569
rect 20990 14560 20996 14572
rect 21048 14560 21054 14612
rect 23385 14603 23443 14609
rect 23385 14569 23397 14603
rect 23431 14600 23443 14603
rect 24581 14603 24639 14609
rect 24581 14600 24593 14603
rect 23431 14572 24593 14600
rect 23431 14569 23443 14572
rect 23385 14563 23443 14569
rect 24581 14569 24593 14572
rect 24627 14569 24639 14603
rect 24581 14563 24639 14569
rect 30193 14603 30251 14609
rect 30193 14569 30205 14603
rect 30239 14600 30251 14603
rect 31478 14600 31484 14612
rect 30239 14572 31484 14600
rect 30239 14569 30251 14572
rect 30193 14563 30251 14569
rect 31478 14560 31484 14572
rect 31536 14560 31542 14612
rect 40221 14603 40279 14609
rect 40221 14569 40233 14603
rect 40267 14600 40279 14603
rect 41322 14600 41328 14612
rect 40267 14572 41328 14600
rect 40267 14569 40279 14572
rect 40221 14563 40279 14569
rect 41322 14560 41328 14572
rect 41380 14560 41386 14612
rect 10428 14504 16804 14532
rect 4982 14464 4988 14476
rect 4943 14436 4988 14464
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 5169 14467 5227 14473
rect 5169 14433 5181 14467
rect 5215 14464 5227 14467
rect 5994 14464 6000 14476
rect 5215 14436 6000 14464
rect 5215 14433 5227 14436
rect 5169 14427 5227 14433
rect 5994 14424 6000 14436
rect 6052 14424 6058 14476
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 10428 14464 10456 14504
rect 16942 14492 16948 14544
rect 17000 14532 17006 14544
rect 22373 14535 22431 14541
rect 17000 14504 21864 14532
rect 17000 14492 17006 14504
rect 17129 14467 17187 14473
rect 17129 14464 17141 14467
rect 9732 14436 10456 14464
rect 9732 14424 9738 14436
rect 2590 14396 2596 14408
rect 2551 14368 2596 14396
rect 2590 14356 2596 14368
rect 2648 14356 2654 14408
rect 7098 14356 7104 14408
rect 7156 14396 7162 14408
rect 7478 14399 7536 14405
rect 7478 14396 7490 14399
rect 7156 14368 7490 14396
rect 7156 14356 7162 14368
rect 7478 14365 7490 14368
rect 7524 14365 7536 14399
rect 7742 14396 7748 14408
rect 7703 14368 7748 14396
rect 7478 14359 7536 14365
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 10428 14405 10456 14436
rect 16500 14436 17141 14464
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14365 10287 14399
rect 10229 14359 10287 14365
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14365 10471 14399
rect 11974 14396 11980 14408
rect 11935 14368 11980 14396
rect 10413 14359 10471 14365
rect 10244 14328 10272 14359
rect 11974 14356 11980 14368
rect 12032 14356 12038 14408
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 16500 14405 16528 14436
rect 17129 14433 17141 14436
rect 17175 14464 17187 14467
rect 19521 14467 19579 14473
rect 17175 14436 19472 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 16485 14399 16543 14405
rect 16485 14396 16497 14399
rect 14424 14368 16497 14396
rect 14424 14356 14430 14368
rect 16485 14365 16497 14368
rect 16531 14365 16543 14399
rect 16485 14359 16543 14365
rect 16669 14399 16727 14405
rect 16669 14365 16681 14399
rect 16715 14365 16727 14399
rect 16669 14359 16727 14365
rect 16684 14328 16712 14359
rect 19334 14356 19340 14408
rect 19392 14396 19398 14408
rect 19444 14405 19472 14436
rect 19521 14433 19533 14467
rect 19567 14464 19579 14467
rect 19567 14436 20208 14464
rect 19567 14433 19579 14436
rect 19521 14427 19579 14433
rect 20180 14408 20208 14436
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 19392 14368 19441 14396
rect 19392 14356 19398 14368
rect 19429 14365 19441 14368
rect 19475 14365 19487 14399
rect 19610 14396 19616 14408
rect 19571 14368 19616 14396
rect 19429 14359 19487 14365
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 20162 14396 20168 14408
rect 20123 14368 20168 14396
rect 20162 14356 20168 14368
rect 20220 14356 20226 14408
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20809 14399 20867 14405
rect 20809 14396 20821 14399
rect 20404 14368 20821 14396
rect 20404 14356 20410 14368
rect 20809 14365 20821 14368
rect 20855 14365 20867 14399
rect 20809 14359 20867 14365
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14396 21051 14399
rect 21358 14396 21364 14408
rect 21039 14368 21364 14396
rect 21039 14365 21051 14368
rect 20993 14359 21051 14365
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 21836 14405 21864 14504
rect 22373 14501 22385 14535
rect 22419 14532 22431 14535
rect 24946 14532 24952 14544
rect 22419 14504 24952 14532
rect 22419 14501 22431 14504
rect 22373 14495 22431 14501
rect 24946 14492 24952 14504
rect 25004 14492 25010 14544
rect 26970 14492 26976 14544
rect 27028 14532 27034 14544
rect 27028 14504 31754 14532
rect 27028 14492 27034 14504
rect 22554 14464 22560 14476
rect 22020 14436 22560 14464
rect 22020 14405 22048 14436
rect 22554 14424 22560 14436
rect 22612 14464 22618 14476
rect 24118 14464 24124 14476
rect 22612 14436 23060 14464
rect 22612 14424 22618 14436
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14365 21879 14399
rect 21821 14359 21879 14365
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 22189 14399 22247 14405
rect 22189 14365 22201 14399
rect 22235 14396 22247 14399
rect 22646 14396 22652 14408
rect 22235 14368 22652 14396
rect 22235 14365 22247 14368
rect 22189 14359 22247 14365
rect 22646 14356 22652 14368
rect 22704 14356 22710 14408
rect 22830 14396 22836 14408
rect 22791 14368 22836 14396
rect 22830 14356 22836 14368
rect 22888 14356 22894 14408
rect 23032 14405 23060 14436
rect 23124 14436 24124 14464
rect 23124 14405 23152 14436
rect 24118 14424 24124 14436
rect 24176 14424 24182 14476
rect 24394 14424 24400 14476
rect 24452 14464 24458 14476
rect 24673 14467 24731 14473
rect 24673 14464 24685 14467
rect 24452 14436 24685 14464
rect 24452 14424 24458 14436
rect 24673 14433 24685 14436
rect 24719 14433 24731 14467
rect 28353 14467 28411 14473
rect 28353 14464 28365 14467
rect 24673 14427 24731 14433
rect 27724 14436 28365 14464
rect 23017 14399 23075 14405
rect 23017 14365 23029 14399
rect 23063 14365 23075 14399
rect 23017 14359 23075 14365
rect 23109 14399 23167 14405
rect 23109 14365 23121 14399
rect 23155 14365 23167 14399
rect 23109 14359 23167 14365
rect 23198 14356 23204 14408
rect 23256 14396 23262 14408
rect 24581 14399 24639 14405
rect 23256 14368 23301 14396
rect 23256 14356 23262 14368
rect 24581 14365 24593 14399
rect 24627 14396 24639 14399
rect 24762 14396 24768 14408
rect 24627 14368 24768 14396
rect 24627 14365 24639 14368
rect 24581 14359 24639 14365
rect 24762 14356 24768 14368
rect 24820 14356 24826 14408
rect 24857 14399 24915 14405
rect 24857 14365 24869 14399
rect 24903 14396 24915 14399
rect 25038 14396 25044 14408
rect 24903 14368 25044 14396
rect 24903 14365 24915 14368
rect 24857 14359 24915 14365
rect 25038 14356 25044 14368
rect 25096 14356 25102 14408
rect 26789 14399 26847 14405
rect 26789 14365 26801 14399
rect 26835 14396 26847 14399
rect 26970 14396 26976 14408
rect 26835 14368 26976 14396
rect 26835 14365 26847 14368
rect 26789 14359 26847 14365
rect 26970 14356 26976 14368
rect 27028 14356 27034 14408
rect 27522 14396 27528 14408
rect 27483 14368 27528 14396
rect 27522 14356 27528 14368
rect 27580 14356 27586 14408
rect 27724 14405 27752 14436
rect 28353 14433 28365 14436
rect 28399 14433 28411 14467
rect 28353 14427 28411 14433
rect 27617 14399 27675 14405
rect 27617 14365 27629 14399
rect 27663 14365 27675 14399
rect 27617 14359 27675 14365
rect 27709 14399 27767 14405
rect 27709 14365 27721 14399
rect 27755 14365 27767 14399
rect 27709 14359 27767 14365
rect 27893 14399 27951 14405
rect 27893 14365 27905 14399
rect 27939 14396 27951 14399
rect 28258 14396 28264 14408
rect 27939 14368 28264 14396
rect 27939 14365 27951 14368
rect 27893 14359 27951 14365
rect 21726 14328 21732 14340
rect 10244 14300 10824 14328
rect 10796 14272 10824 14300
rect 16684 14300 21732 14328
rect 4893 14263 4951 14269
rect 4893 14229 4905 14263
rect 4939 14260 4951 14263
rect 5810 14260 5816 14272
rect 4939 14232 5816 14260
rect 4939 14229 4951 14232
rect 4893 14223 4951 14229
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 9674 14260 9680 14272
rect 9635 14232 9680 14260
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 10873 14263 10931 14269
rect 10873 14260 10885 14263
rect 10836 14232 10885 14260
rect 10836 14220 10842 14232
rect 10873 14229 10885 14232
rect 10919 14229 10931 14263
rect 12066 14260 12072 14272
rect 12027 14232 12072 14260
rect 10873 14223 10931 14229
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 15933 14263 15991 14269
rect 15933 14260 15945 14263
rect 13688 14232 15945 14260
rect 13688 14220 13694 14232
rect 15933 14229 15945 14232
rect 15979 14260 15991 14263
rect 16684 14260 16712 14300
rect 21726 14288 21732 14300
rect 21784 14328 21790 14340
rect 21910 14328 21916 14340
rect 21784 14300 21916 14328
rect 21784 14288 21790 14300
rect 21910 14288 21916 14300
rect 21968 14288 21974 14340
rect 22097 14331 22155 14337
rect 22097 14297 22109 14331
rect 22143 14297 22155 14331
rect 22097 14291 22155 14297
rect 15979 14232 16712 14260
rect 22112 14260 22140 14291
rect 23290 14288 23296 14340
rect 23348 14328 23354 14340
rect 26544 14331 26602 14337
rect 23348 14300 25452 14328
rect 23348 14288 23354 14300
rect 23934 14260 23940 14272
rect 22112 14232 23940 14260
rect 15979 14229 15991 14232
rect 15933 14223 15991 14229
rect 23934 14220 23940 14232
rect 23992 14220 23998 14272
rect 24302 14220 24308 14272
rect 24360 14260 24366 14272
rect 25424 14269 25452 14300
rect 26544 14297 26556 14331
rect 26590 14328 26602 14331
rect 27249 14331 27307 14337
rect 27249 14328 27261 14331
rect 26590 14300 27261 14328
rect 26590 14297 26602 14300
rect 26544 14291 26602 14297
rect 27249 14297 27261 14300
rect 27295 14297 27307 14331
rect 27632 14328 27660 14359
rect 28258 14356 28264 14368
rect 28316 14356 28322 14408
rect 28721 14399 28779 14405
rect 28721 14365 28733 14399
rect 28767 14396 28779 14399
rect 29362 14396 29368 14408
rect 28767 14368 29368 14396
rect 28767 14365 28779 14368
rect 28721 14359 28779 14365
rect 29362 14356 29368 14368
rect 29420 14396 29426 14408
rect 29822 14396 29828 14408
rect 29420 14368 29828 14396
rect 29420 14356 29426 14368
rect 29822 14356 29828 14368
rect 29880 14356 29886 14408
rect 31726 14396 31754 14504
rect 40862 14492 40868 14544
rect 40920 14532 40926 14544
rect 40957 14535 41015 14541
rect 40957 14532 40969 14535
rect 40920 14504 40969 14532
rect 40920 14492 40926 14504
rect 40957 14501 40969 14504
rect 41003 14501 41015 14535
rect 40957 14495 41015 14501
rect 32030 14424 32036 14476
rect 32088 14464 32094 14476
rect 33505 14467 33563 14473
rect 33505 14464 33517 14467
rect 32088 14436 33517 14464
rect 32088 14424 32094 14436
rect 33505 14433 33517 14436
rect 33551 14433 33563 14467
rect 33505 14427 33563 14433
rect 33594 14424 33600 14476
rect 33652 14464 33658 14476
rect 33781 14467 33839 14473
rect 33781 14464 33793 14467
rect 33652 14436 33793 14464
rect 33652 14424 33658 14436
rect 33781 14433 33793 14436
rect 33827 14433 33839 14467
rect 34698 14464 34704 14476
rect 34659 14436 34704 14464
rect 33781 14427 33839 14433
rect 34698 14424 34704 14436
rect 34756 14424 34762 14476
rect 35802 14424 35808 14476
rect 35860 14464 35866 14476
rect 35989 14467 36047 14473
rect 35989 14464 36001 14467
rect 35860 14436 36001 14464
rect 35860 14424 35866 14436
rect 35989 14433 36001 14436
rect 36035 14433 36047 14467
rect 35989 14427 36047 14433
rect 33410 14396 33416 14408
rect 31726 14368 33416 14396
rect 33410 14356 33416 14368
rect 33468 14356 33474 14408
rect 34790 14356 34796 14408
rect 34848 14396 34854 14408
rect 34977 14399 35035 14405
rect 34977 14396 34989 14399
rect 34848 14368 34989 14396
rect 34848 14356 34854 14368
rect 34977 14365 34989 14368
rect 35023 14396 35035 14399
rect 35710 14396 35716 14408
rect 35023 14368 35716 14396
rect 35023 14365 35035 14368
rect 34977 14359 35035 14365
rect 35710 14356 35716 14368
rect 35768 14356 35774 14408
rect 36173 14399 36231 14405
rect 36173 14365 36185 14399
rect 36219 14365 36231 14399
rect 36173 14359 36231 14365
rect 27798 14328 27804 14340
rect 27632 14300 27804 14328
rect 27249 14291 27307 14297
rect 27798 14288 27804 14300
rect 27856 14288 27862 14340
rect 28537 14331 28595 14337
rect 28537 14297 28549 14331
rect 28583 14297 28595 14331
rect 28537 14291 28595 14297
rect 24397 14263 24455 14269
rect 24397 14260 24409 14263
rect 24360 14232 24409 14260
rect 24360 14220 24366 14232
rect 24397 14229 24409 14232
rect 24443 14229 24455 14263
rect 24397 14223 24455 14229
rect 25409 14263 25467 14269
rect 25409 14229 25421 14263
rect 25455 14260 25467 14263
rect 28552 14260 28580 14291
rect 29546 14288 29552 14340
rect 29604 14328 29610 14340
rect 30009 14331 30067 14337
rect 30009 14328 30021 14331
rect 29604 14300 30021 14328
rect 29604 14288 29610 14300
rect 30009 14297 30021 14300
rect 30055 14297 30067 14331
rect 36188 14328 36216 14359
rect 36906 14356 36912 14408
rect 36964 14396 36970 14408
rect 37182 14396 37188 14408
rect 36964 14368 37188 14396
rect 36964 14356 36970 14368
rect 37182 14356 37188 14368
rect 37240 14356 37246 14408
rect 38930 14356 38936 14408
rect 38988 14396 38994 14408
rect 40037 14399 40095 14405
rect 40037 14396 40049 14399
rect 38988 14368 40049 14396
rect 38988 14356 38994 14368
rect 40037 14365 40049 14368
rect 40083 14365 40095 14399
rect 40037 14359 40095 14365
rect 40678 14356 40684 14408
rect 40736 14396 40742 14408
rect 40773 14399 40831 14405
rect 40773 14396 40785 14399
rect 40736 14368 40785 14396
rect 40736 14356 40742 14368
rect 40773 14365 40785 14368
rect 40819 14365 40831 14399
rect 58158 14396 58164 14408
rect 58119 14368 58164 14396
rect 40773 14359 40831 14365
rect 58158 14356 58164 14368
rect 58216 14356 58222 14408
rect 30009 14291 30067 14297
rect 35728 14300 36216 14328
rect 35728 14272 35756 14300
rect 39482 14288 39488 14340
rect 39540 14328 39546 14340
rect 39850 14328 39856 14340
rect 39540 14300 39856 14328
rect 39540 14288 39546 14300
rect 39850 14288 39856 14300
rect 39908 14288 39914 14340
rect 25455 14232 28580 14260
rect 25455 14229 25467 14232
rect 25409 14223 25467 14229
rect 35710 14220 35716 14272
rect 35768 14220 35774 14272
rect 36357 14263 36415 14269
rect 36357 14229 36369 14263
rect 36403 14260 36415 14263
rect 37642 14260 37648 14272
rect 36403 14232 37648 14260
rect 36403 14229 36415 14232
rect 36357 14223 36415 14229
rect 37642 14220 37648 14232
rect 37700 14220 37706 14272
rect 38102 14220 38108 14272
rect 38160 14260 38166 14272
rect 38473 14263 38531 14269
rect 38473 14260 38485 14263
rect 38160 14232 38485 14260
rect 38160 14220 38166 14232
rect 38473 14229 38485 14232
rect 38519 14229 38531 14263
rect 38473 14223 38531 14229
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 2682 14016 2688 14068
rect 2740 14056 2746 14068
rect 2961 14059 3019 14065
rect 2961 14056 2973 14059
rect 2740 14028 2973 14056
rect 2740 14016 2746 14028
rect 2961 14025 2973 14028
rect 3007 14025 3019 14059
rect 19334 14056 19340 14068
rect 19295 14028 19340 14056
rect 2961 14019 3019 14025
rect 19334 14016 19340 14028
rect 19392 14056 19398 14068
rect 20717 14059 20775 14065
rect 20717 14056 20729 14059
rect 19392 14028 20729 14056
rect 19392 14016 19398 14028
rect 20717 14025 20729 14028
rect 20763 14056 20775 14059
rect 21266 14056 21272 14068
rect 20763 14028 21272 14056
rect 20763 14025 20775 14028
rect 20717 14019 20775 14025
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 22094 14016 22100 14068
rect 22152 14056 22158 14068
rect 22152 14028 22197 14056
rect 22152 14016 22158 14028
rect 22554 14016 22560 14068
rect 22612 14056 22618 14068
rect 23658 14056 23664 14068
rect 22612 14028 22784 14056
rect 23619 14028 23664 14056
rect 22612 14016 22618 14028
rect 10778 13948 10784 14000
rect 10836 13988 10842 14000
rect 22186 13988 22192 14000
rect 10836 13960 22192 13988
rect 10836 13948 10842 13960
rect 22186 13948 22192 13960
rect 22244 13948 22250 14000
rect 22756 13997 22784 14028
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 23934 14016 23940 14068
rect 23992 14056 23998 14068
rect 24578 14056 24584 14068
rect 23992 14028 24440 14056
rect 24539 14028 24584 14056
rect 23992 14016 23998 14028
rect 22741 13991 22799 13997
rect 22741 13957 22753 13991
rect 22787 13957 22799 13991
rect 22741 13951 22799 13957
rect 22833 13991 22891 13997
rect 22833 13957 22845 13991
rect 22879 13988 22891 13991
rect 23290 13988 23296 14000
rect 22879 13960 23296 13988
rect 22879 13957 22891 13960
rect 22833 13951 22891 13957
rect 23290 13948 23296 13960
rect 23348 13948 23354 14000
rect 24121 13991 24179 13997
rect 24121 13957 24133 13991
rect 24167 13988 24179 13991
rect 24210 13988 24216 14000
rect 24167 13960 24216 13988
rect 24167 13957 24179 13960
rect 24121 13951 24179 13957
rect 24210 13948 24216 13960
rect 24268 13948 24274 14000
rect 24412 13988 24440 14028
rect 24578 14016 24584 14028
rect 24636 14016 24642 14068
rect 25590 14056 25596 14068
rect 25551 14028 25596 14056
rect 25590 14016 25596 14028
rect 25648 14016 25654 14068
rect 26421 14059 26479 14065
rect 26421 14025 26433 14059
rect 26467 14056 26479 14059
rect 26602 14056 26608 14068
rect 26467 14028 26608 14056
rect 26467 14025 26479 14028
rect 26421 14019 26479 14025
rect 26602 14016 26608 14028
rect 26660 14056 26666 14068
rect 27522 14056 27528 14068
rect 26660 14028 27528 14056
rect 26660 14016 26666 14028
rect 27522 14016 27528 14028
rect 27580 14016 27586 14068
rect 27614 14016 27620 14068
rect 27672 14056 27678 14068
rect 28353 14059 28411 14065
rect 28353 14056 28365 14059
rect 27672 14028 28365 14056
rect 27672 14016 27678 14028
rect 28353 14025 28365 14028
rect 28399 14025 28411 14059
rect 37458 14056 37464 14068
rect 28353 14019 28411 14025
rect 34532 14028 37464 14056
rect 24412 13960 27614 13988
rect 3145 13923 3203 13929
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 4614 13920 4620 13932
rect 3191 13892 4620 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 6362 13880 6368 13932
rect 6420 13920 6426 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 6420 13892 7297 13920
rect 6420 13880 6426 13892
rect 7285 13889 7297 13892
rect 7331 13920 7343 13923
rect 12066 13920 12072 13932
rect 7331 13892 12072 13920
rect 7331 13889 7343 13892
rect 7285 13883 7343 13889
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 14274 13920 14280 13932
rect 14332 13929 14338 13932
rect 14244 13892 14280 13920
rect 14274 13880 14280 13892
rect 14332 13883 14344 13929
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13920 14611 13923
rect 15102 13920 15108 13932
rect 14599 13892 15108 13920
rect 14599 13889 14611 13892
rect 14553 13883 14611 13889
rect 14332 13880 14338 13883
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 20622 13880 20628 13932
rect 20680 13920 20686 13932
rect 22557 13923 22615 13929
rect 22557 13920 22569 13923
rect 20680 13892 22569 13920
rect 20680 13880 20686 13892
rect 22557 13889 22569 13892
rect 22603 13889 22615 13923
rect 22557 13883 22615 13889
rect 22646 13880 22652 13932
rect 22704 13920 22710 13932
rect 22925 13923 22983 13929
rect 22925 13920 22937 13923
rect 22704 13892 22937 13920
rect 22704 13880 22710 13892
rect 22925 13889 22937 13892
rect 22971 13920 22983 13923
rect 23198 13920 23204 13932
rect 22971 13892 23204 13920
rect 22971 13889 22983 13892
rect 22925 13883 22983 13889
rect 23198 13880 23204 13892
rect 23256 13880 23262 13932
rect 23845 13923 23903 13929
rect 23845 13889 23857 13923
rect 23891 13920 23903 13923
rect 24486 13920 24492 13932
rect 23891 13892 24492 13920
rect 23891 13889 23903 13892
rect 23845 13883 23903 13889
rect 24486 13880 24492 13892
rect 24544 13880 24550 13932
rect 24765 13923 24823 13929
rect 24765 13920 24777 13923
rect 24688 13892 24777 13920
rect 3786 13812 3792 13864
rect 3844 13852 3850 13864
rect 7742 13852 7748 13864
rect 3844 13824 7748 13852
rect 3844 13812 3850 13824
rect 7742 13812 7748 13824
rect 7800 13812 7806 13864
rect 21358 13812 21364 13864
rect 21416 13852 21422 13864
rect 23474 13852 23480 13864
rect 21416 13824 23480 13852
rect 21416 13812 21422 13824
rect 23474 13812 23480 13824
rect 23532 13812 23538 13864
rect 23566 13812 23572 13864
rect 23624 13852 23630 13864
rect 23937 13855 23995 13861
rect 23937 13852 23949 13855
rect 23624 13824 23949 13852
rect 23624 13812 23630 13824
rect 23937 13821 23949 13824
rect 23983 13821 23995 13855
rect 23937 13815 23995 13821
rect 23109 13787 23167 13793
rect 23109 13753 23121 13787
rect 23155 13784 23167 13787
rect 24688 13784 24716 13892
rect 24765 13889 24777 13892
rect 24811 13889 24823 13923
rect 24765 13883 24823 13889
rect 25041 13923 25099 13929
rect 25041 13889 25053 13923
rect 25087 13920 25099 13923
rect 25590 13920 25596 13932
rect 25087 13892 25596 13920
rect 25087 13889 25099 13892
rect 25041 13883 25099 13889
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 26142 13880 26148 13932
rect 26200 13920 26206 13932
rect 26970 13920 26976 13932
rect 26200 13892 26976 13920
rect 26200 13880 26206 13892
rect 26970 13880 26976 13892
rect 27028 13880 27034 13932
rect 27246 13929 27252 13932
rect 27240 13883 27252 13929
rect 27304 13920 27310 13932
rect 27586 13920 27614 13960
rect 27304 13892 27340 13920
rect 27586 13892 29592 13920
rect 27246 13880 27252 13883
rect 27304 13880 27310 13892
rect 24854 13852 24860 13864
rect 24815 13824 24860 13852
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 29564 13796 29592 13892
rect 30374 13880 30380 13932
rect 30432 13920 30438 13932
rect 30662 13923 30720 13929
rect 30662 13920 30674 13923
rect 30432 13892 30674 13920
rect 30432 13880 30438 13892
rect 30662 13889 30674 13892
rect 30708 13889 30720 13923
rect 30926 13920 30932 13932
rect 30887 13892 30932 13920
rect 30662 13883 30720 13889
rect 30926 13880 30932 13892
rect 30984 13880 30990 13932
rect 33410 13880 33416 13932
rect 33468 13920 33474 13932
rect 33965 13923 34023 13929
rect 33965 13920 33977 13923
rect 33468 13892 33977 13920
rect 33468 13880 33474 13892
rect 33965 13889 33977 13892
rect 34011 13920 34023 13923
rect 34425 13923 34483 13929
rect 34425 13920 34437 13923
rect 34011 13892 34437 13920
rect 34011 13889 34023 13892
rect 33965 13883 34023 13889
rect 34425 13889 34437 13892
rect 34471 13920 34483 13923
rect 34532 13920 34560 14028
rect 37458 14016 37464 14028
rect 37516 14016 37522 14068
rect 36538 13988 36544 14000
rect 36499 13960 36544 13988
rect 36538 13948 36544 13960
rect 36596 13948 36602 14000
rect 39209 13991 39267 13997
rect 39209 13988 39221 13991
rect 36648 13960 39221 13988
rect 34471 13892 34560 13920
rect 34609 13923 34667 13929
rect 34471 13889 34483 13892
rect 34425 13883 34483 13889
rect 34609 13889 34621 13923
rect 34655 13920 34667 13923
rect 34790 13920 34796 13932
rect 34655 13892 34796 13920
rect 34655 13889 34667 13892
rect 34609 13883 34667 13889
rect 34790 13880 34796 13892
rect 34848 13880 34854 13932
rect 35897 13923 35955 13929
rect 35897 13920 35909 13923
rect 35452 13892 35909 13920
rect 33594 13812 33600 13864
rect 33652 13852 33658 13864
rect 35452 13852 35480 13892
rect 35897 13889 35909 13892
rect 35943 13920 35955 13923
rect 36648 13920 36676 13960
rect 39209 13957 39221 13960
rect 39255 13988 39267 13991
rect 40678 13988 40684 14000
rect 39255 13960 40684 13988
rect 39255 13957 39267 13960
rect 39209 13951 39267 13957
rect 40678 13948 40684 13960
rect 40736 13948 40742 14000
rect 35943 13892 36676 13920
rect 35943 13889 35955 13892
rect 35897 13883 35955 13889
rect 36722 13880 36728 13932
rect 36780 13920 36786 13932
rect 38562 13920 38568 13932
rect 36780 13892 38240 13920
rect 38523 13892 38568 13920
rect 36780 13880 36786 13892
rect 35618 13852 35624 13864
rect 33652 13824 35480 13852
rect 35579 13824 35624 13852
rect 33652 13812 33658 13824
rect 35618 13812 35624 13824
rect 35676 13812 35682 13864
rect 25866 13784 25872 13796
rect 23155 13756 23888 13784
rect 24688 13756 25872 13784
rect 23155 13753 23167 13756
rect 23109 13747 23167 13753
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 7745 13719 7803 13725
rect 7745 13716 7757 13719
rect 7708 13688 7757 13716
rect 7708 13676 7714 13688
rect 7745 13685 7757 13688
rect 7791 13685 7803 13719
rect 13170 13716 13176 13728
rect 13131 13688 13176 13716
rect 7745 13679 7803 13685
rect 13170 13676 13176 13688
rect 13228 13676 13234 13728
rect 18690 13716 18696 13728
rect 18651 13688 18696 13716
rect 18690 13676 18696 13688
rect 18748 13676 18754 13728
rect 19889 13719 19947 13725
rect 19889 13685 19901 13719
rect 19935 13716 19947 13719
rect 20070 13716 20076 13728
rect 19935 13688 20076 13716
rect 19935 13685 19947 13688
rect 19889 13679 19947 13685
rect 20070 13676 20076 13688
rect 20128 13676 20134 13728
rect 23860 13725 23888 13756
rect 25866 13744 25872 13756
rect 25924 13744 25930 13796
rect 29546 13784 29552 13796
rect 29459 13756 29552 13784
rect 29546 13744 29552 13756
rect 29604 13744 29610 13796
rect 34517 13787 34575 13793
rect 34517 13753 34529 13787
rect 34563 13784 34575 13787
rect 35986 13784 35992 13796
rect 34563 13756 35992 13784
rect 34563 13753 34575 13756
rect 34517 13747 34575 13753
rect 35986 13744 35992 13756
rect 36044 13744 36050 13796
rect 38212 13784 38240 13892
rect 38562 13880 38568 13892
rect 38620 13880 38626 13932
rect 38289 13855 38347 13861
rect 38289 13821 38301 13855
rect 38335 13852 38347 13855
rect 38378 13852 38384 13864
rect 38335 13824 38384 13852
rect 38335 13821 38347 13824
rect 38289 13815 38347 13821
rect 38378 13812 38384 13824
rect 38436 13812 38442 13864
rect 39482 13852 39488 13864
rect 38580 13824 39488 13852
rect 38580 13784 38608 13824
rect 39482 13812 39488 13824
rect 39540 13812 39546 13864
rect 40402 13852 40408 13864
rect 39960 13824 40408 13852
rect 39960 13784 39988 13824
rect 40402 13812 40408 13824
rect 40460 13812 40466 13864
rect 38212 13756 38608 13784
rect 39316 13756 39988 13784
rect 39316 13728 39344 13756
rect 23845 13719 23903 13725
rect 23845 13685 23857 13719
rect 23891 13685 23903 13719
rect 24946 13716 24952 13728
rect 24907 13688 24952 13716
rect 23845 13679 23903 13685
rect 24946 13676 24952 13688
rect 25004 13676 25010 13728
rect 35894 13676 35900 13728
rect 35952 13716 35958 13728
rect 36357 13719 36415 13725
rect 36357 13716 36369 13719
rect 35952 13688 36369 13716
rect 35952 13676 35958 13688
rect 36357 13685 36369 13688
rect 36403 13685 36415 13719
rect 39298 13716 39304 13728
rect 39259 13688 39304 13716
rect 36357 13679 36415 13685
rect 39298 13676 39304 13688
rect 39356 13676 39362 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 14274 13512 14280 13524
rect 14235 13484 14280 13512
rect 14274 13472 14280 13484
rect 14332 13472 14338 13524
rect 18782 13472 18788 13524
rect 18840 13512 18846 13524
rect 22002 13512 22008 13524
rect 18840 13484 22008 13512
rect 18840 13472 18846 13484
rect 22002 13472 22008 13484
rect 22060 13512 22066 13524
rect 23658 13512 23664 13524
rect 22060 13484 23664 13512
rect 22060 13472 22066 13484
rect 23658 13472 23664 13484
rect 23716 13472 23722 13524
rect 27246 13512 27252 13524
rect 27207 13484 27252 13512
rect 27246 13472 27252 13484
rect 27304 13472 27310 13524
rect 28997 13515 29055 13521
rect 28997 13481 29009 13515
rect 29043 13512 29055 13515
rect 29086 13512 29092 13524
rect 29043 13484 29092 13512
rect 29043 13481 29055 13484
rect 28997 13475 29055 13481
rect 29086 13472 29092 13484
rect 29144 13512 29150 13524
rect 30006 13512 30012 13524
rect 29144 13484 30012 13512
rect 29144 13472 29150 13484
rect 30006 13472 30012 13484
rect 30064 13472 30070 13524
rect 30285 13515 30343 13521
rect 30285 13481 30297 13515
rect 30331 13512 30343 13515
rect 30374 13512 30380 13524
rect 30331 13484 30380 13512
rect 30331 13481 30343 13484
rect 30285 13475 30343 13481
rect 30374 13472 30380 13484
rect 30432 13472 30438 13524
rect 34977 13515 35035 13521
rect 34977 13481 34989 13515
rect 35023 13512 35035 13515
rect 35802 13512 35808 13524
rect 35023 13484 35808 13512
rect 35023 13481 35035 13484
rect 34977 13475 35035 13481
rect 35802 13472 35808 13484
rect 35860 13472 35866 13524
rect 36538 13472 36544 13524
rect 36596 13512 36602 13524
rect 36817 13515 36875 13521
rect 36817 13512 36829 13515
rect 36596 13484 36829 13512
rect 36596 13472 36602 13484
rect 36817 13481 36829 13484
rect 36863 13481 36875 13515
rect 36817 13475 36875 13481
rect 17678 13404 17684 13456
rect 17736 13444 17742 13456
rect 19337 13447 19395 13453
rect 19337 13444 19349 13447
rect 17736 13416 19349 13444
rect 17736 13404 17742 13416
rect 19337 13413 19349 13416
rect 19383 13413 19395 13447
rect 19337 13407 19395 13413
rect 12526 13336 12532 13388
rect 12584 13376 12590 13388
rect 19058 13376 19064 13388
rect 12584 13348 19064 13376
rect 12584 13336 12590 13348
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13308 5963 13311
rect 7653 13311 7711 13317
rect 5951 13280 6914 13308
rect 5951 13277 5963 13280
rect 5905 13271 5963 13277
rect 6886 13172 6914 13280
rect 7653 13277 7665 13311
rect 7699 13308 7711 13311
rect 7742 13308 7748 13320
rect 7699 13280 7748 13308
rect 7699 13277 7711 13280
rect 7653 13271 7711 13277
rect 7742 13268 7748 13280
rect 7800 13308 7806 13320
rect 8754 13308 8760 13320
rect 7800 13280 8760 13308
rect 7800 13268 7806 13280
rect 8754 13268 8760 13280
rect 8812 13308 8818 13320
rect 9677 13311 9735 13317
rect 9677 13308 9689 13311
rect 8812 13280 9689 13308
rect 8812 13268 8818 13280
rect 9677 13277 9689 13280
rect 9723 13277 9735 13311
rect 9677 13271 9735 13277
rect 13541 13311 13599 13317
rect 13541 13277 13553 13311
rect 13587 13308 13599 13311
rect 14274 13308 14280 13320
rect 13587 13280 14280 13308
rect 13587 13277 13599 13280
rect 13541 13271 13599 13277
rect 14274 13268 14280 13280
rect 14332 13308 14338 13320
rect 14553 13311 14611 13317
rect 14553 13308 14565 13311
rect 14332 13280 14565 13308
rect 14332 13268 14338 13280
rect 14553 13277 14565 13280
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 14645 13311 14703 13317
rect 14645 13277 14657 13311
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 14737 13311 14795 13317
rect 14737 13277 14749 13311
rect 14783 13308 14795 13311
rect 14826 13308 14832 13320
rect 14783 13280 14832 13308
rect 14783 13277 14795 13280
rect 14737 13271 14795 13277
rect 9766 13200 9772 13252
rect 9824 13240 9830 13252
rect 9922 13243 9980 13249
rect 9922 13240 9934 13243
rect 9824 13212 9934 13240
rect 9824 13200 9830 13212
rect 9922 13209 9934 13212
rect 9968 13209 9980 13243
rect 9922 13203 9980 13209
rect 8205 13175 8263 13181
rect 8205 13172 8217 13175
rect 6886 13144 8217 13172
rect 8205 13141 8217 13144
rect 8251 13172 8263 13175
rect 8294 13172 8300 13184
rect 8251 13144 8300 13172
rect 8251 13141 8263 13144
rect 8205 13135 8263 13141
rect 8294 13132 8300 13144
rect 8352 13172 8358 13184
rect 9030 13172 9036 13184
rect 8352 13144 9036 13172
rect 8352 13132 8358 13144
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 10502 13132 10508 13184
rect 10560 13172 10566 13184
rect 11057 13175 11115 13181
rect 11057 13172 11069 13175
rect 10560 13144 11069 13172
rect 10560 13132 10566 13144
rect 11057 13141 11069 13144
rect 11103 13141 11115 13175
rect 11057 13135 11115 13141
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 14660 13172 14688 13271
rect 14826 13268 14832 13280
rect 14884 13268 14890 13320
rect 14921 13311 14979 13317
rect 14921 13277 14933 13311
rect 14967 13308 14979 13311
rect 15010 13308 15016 13320
rect 14967 13280 15016 13308
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 16390 13268 16396 13320
rect 16448 13308 16454 13320
rect 17773 13311 17831 13317
rect 17773 13308 17785 13311
rect 16448 13280 17785 13308
rect 16448 13268 16454 13280
rect 17773 13277 17785 13280
rect 17819 13277 17831 13311
rect 19352 13308 19380 13407
rect 21726 13404 21732 13456
rect 21784 13444 21790 13456
rect 22189 13447 22247 13453
rect 22189 13444 22201 13447
rect 21784 13416 22201 13444
rect 21784 13404 21790 13416
rect 22189 13413 22201 13416
rect 22235 13413 22247 13447
rect 22189 13407 22247 13413
rect 24762 13404 24768 13456
rect 24820 13444 24826 13456
rect 24820 13416 31754 13444
rect 24820 13404 24826 13416
rect 23569 13379 23627 13385
rect 23569 13345 23581 13379
rect 23615 13376 23627 13379
rect 24578 13376 24584 13388
rect 23615 13348 24584 13376
rect 23615 13345 23627 13348
rect 23569 13339 23627 13345
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 27798 13376 27804 13388
rect 27632 13348 27804 13376
rect 19981 13311 20039 13317
rect 19981 13308 19993 13311
rect 19352 13280 19993 13308
rect 17773 13271 17831 13277
rect 19981 13277 19993 13280
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 23750 13268 23756 13320
rect 23808 13308 23814 13320
rect 27632 13317 27660 13348
rect 27798 13336 27804 13348
rect 27856 13336 27862 13388
rect 28258 13376 28264 13388
rect 27908 13348 28264 13376
rect 23845 13311 23903 13317
rect 23845 13308 23857 13311
rect 23808 13280 23857 13308
rect 23808 13268 23814 13280
rect 23845 13277 23857 13280
rect 23891 13308 23903 13311
rect 24765 13311 24823 13317
rect 24765 13308 24777 13311
rect 23891 13280 24777 13308
rect 23891 13277 23903 13280
rect 23845 13271 23903 13277
rect 24765 13277 24777 13280
rect 24811 13277 24823 13311
rect 27525 13311 27583 13317
rect 27525 13308 27537 13311
rect 24765 13271 24823 13277
rect 26804 13280 27537 13308
rect 16666 13200 16672 13252
rect 16724 13240 16730 13252
rect 17589 13243 17647 13249
rect 17589 13240 17601 13243
rect 16724 13212 17601 13240
rect 16724 13200 16730 13212
rect 17589 13209 17601 13212
rect 17635 13209 17647 13243
rect 17589 13203 17647 13209
rect 20165 13243 20223 13249
rect 20165 13209 20177 13243
rect 20211 13240 20223 13243
rect 22186 13240 22192 13252
rect 20211 13212 22192 13240
rect 20211 13209 20223 13212
rect 20165 13203 20223 13209
rect 22186 13200 22192 13212
rect 22244 13200 22250 13252
rect 22370 13200 22376 13252
rect 22428 13240 22434 13252
rect 24949 13243 25007 13249
rect 24949 13240 24961 13243
rect 22428 13212 24961 13240
rect 22428 13200 22434 13212
rect 24949 13209 24961 13212
rect 24995 13240 25007 13243
rect 25498 13240 25504 13252
rect 24995 13212 25504 13240
rect 24995 13209 25007 13212
rect 24949 13203 25007 13209
rect 25498 13200 25504 13212
rect 25556 13200 25562 13252
rect 26804 13184 26832 13280
rect 27525 13277 27537 13280
rect 27571 13277 27583 13311
rect 27525 13271 27583 13277
rect 27617 13311 27675 13317
rect 27617 13277 27629 13311
rect 27663 13277 27675 13311
rect 27617 13271 27675 13277
rect 14608 13144 14688 13172
rect 14608 13132 14614 13144
rect 14734 13132 14740 13184
rect 14792 13172 14798 13184
rect 15102 13172 15108 13184
rect 14792 13144 15108 13172
rect 14792 13132 14798 13144
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 17957 13175 18015 13181
rect 17957 13141 17969 13175
rect 18003 13172 18015 13175
rect 18506 13172 18512 13184
rect 18003 13144 18512 13172
rect 18003 13141 18015 13144
rect 17957 13135 18015 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 18693 13175 18751 13181
rect 18693 13141 18705 13175
rect 18739 13172 18751 13175
rect 18966 13172 18972 13184
rect 18739 13144 18972 13172
rect 18739 13141 18751 13144
rect 18693 13135 18751 13141
rect 18966 13132 18972 13144
rect 19024 13132 19030 13184
rect 21177 13175 21235 13181
rect 21177 13141 21189 13175
rect 21223 13172 21235 13175
rect 21358 13172 21364 13184
rect 21223 13144 21364 13172
rect 21223 13141 21235 13144
rect 21177 13135 21235 13141
rect 21358 13132 21364 13144
rect 21416 13132 21422 13184
rect 26786 13172 26792 13184
rect 26747 13144 26792 13172
rect 26786 13132 26792 13144
rect 26844 13132 26850 13184
rect 27632 13172 27660 13271
rect 27706 13268 27712 13320
rect 27764 13308 27770 13320
rect 27908 13317 27936 13348
rect 28258 13336 28264 13348
rect 28316 13376 28322 13388
rect 28353 13379 28411 13385
rect 28353 13376 28365 13379
rect 28316 13348 28365 13376
rect 28316 13336 28322 13348
rect 28353 13345 28365 13348
rect 28399 13345 28411 13379
rect 30558 13376 30564 13388
rect 28353 13339 28411 13345
rect 29656 13348 30564 13376
rect 29656 13317 29684 13348
rect 30558 13336 30564 13348
rect 30616 13336 30622 13388
rect 27893 13311 27951 13317
rect 27764 13280 27809 13308
rect 27764 13268 27770 13280
rect 27893 13277 27905 13311
rect 27939 13277 27951 13311
rect 27893 13271 27951 13277
rect 29641 13311 29699 13317
rect 29641 13277 29653 13311
rect 29687 13277 29699 13311
rect 29641 13271 29699 13277
rect 29730 13268 29736 13320
rect 29788 13308 29794 13320
rect 29825 13311 29883 13317
rect 29825 13308 29837 13311
rect 29788 13280 29837 13308
rect 29788 13268 29794 13280
rect 29825 13277 29837 13280
rect 29871 13277 29883 13311
rect 29825 13271 29883 13277
rect 29917 13311 29975 13317
rect 29917 13277 29929 13311
rect 29963 13277 29975 13311
rect 29917 13271 29975 13277
rect 29932 13184 29960 13271
rect 30006 13268 30012 13320
rect 30064 13308 30070 13320
rect 30064 13280 30109 13308
rect 30064 13268 30070 13280
rect 30650 13268 30656 13320
rect 30708 13308 30714 13320
rect 30837 13311 30895 13317
rect 30837 13308 30849 13311
rect 30708 13280 30849 13308
rect 30708 13268 30714 13280
rect 30837 13277 30849 13280
rect 30883 13308 30895 13311
rect 31202 13308 31208 13320
rect 30883 13280 31208 13308
rect 30883 13277 30895 13280
rect 30837 13271 30895 13277
rect 31202 13268 31208 13280
rect 31260 13268 31266 13320
rect 31726 13308 31754 13416
rect 38378 13404 38384 13456
rect 38436 13444 38442 13456
rect 38436 13416 38608 13444
rect 38436 13404 38442 13416
rect 34149 13379 34207 13385
rect 34149 13345 34161 13379
rect 34195 13376 34207 13379
rect 35437 13379 35495 13385
rect 35437 13376 35449 13379
rect 34195 13348 35449 13376
rect 34195 13345 34207 13348
rect 34149 13339 34207 13345
rect 35437 13345 35449 13348
rect 35483 13345 35495 13379
rect 35437 13339 35495 13345
rect 37737 13379 37795 13385
rect 37737 13345 37749 13379
rect 37783 13376 37795 13379
rect 38580 13376 38608 13416
rect 37783 13348 38424 13376
rect 37783 13345 37795 13348
rect 37737 13339 37795 13345
rect 34422 13308 34428 13320
rect 31726 13280 34428 13308
rect 34422 13268 34428 13280
rect 34480 13268 34486 13320
rect 35452 13308 35480 13339
rect 38102 13308 38108 13320
rect 35452 13280 38108 13308
rect 38102 13268 38108 13280
rect 38160 13268 38166 13320
rect 38396 13317 38424 13348
rect 38488 13348 38608 13376
rect 38488 13317 38516 13348
rect 38197 13311 38255 13317
rect 38197 13277 38209 13311
rect 38243 13277 38255 13311
rect 38197 13271 38255 13277
rect 38381 13311 38439 13317
rect 38381 13277 38393 13311
rect 38427 13277 38439 13311
rect 38381 13271 38439 13277
rect 38473 13311 38531 13317
rect 38473 13277 38485 13311
rect 38519 13277 38531 13311
rect 38473 13271 38531 13277
rect 31021 13243 31079 13249
rect 31021 13209 31033 13243
rect 31067 13240 31079 13243
rect 32306 13240 32312 13252
rect 31067 13212 32312 13240
rect 31067 13209 31079 13212
rect 31021 13203 31079 13209
rect 32306 13200 32312 13212
rect 32364 13200 32370 13252
rect 33318 13200 33324 13252
rect 33376 13240 33382 13252
rect 33882 13243 33940 13249
rect 33882 13240 33894 13243
rect 33376 13212 33894 13240
rect 33376 13200 33382 13212
rect 33882 13209 33894 13212
rect 33928 13209 33940 13243
rect 33882 13203 33940 13209
rect 35434 13200 35440 13252
rect 35492 13240 35498 13252
rect 35682 13243 35740 13249
rect 35682 13240 35694 13243
rect 35492 13212 35694 13240
rect 35492 13200 35498 13212
rect 35682 13209 35694 13212
rect 35728 13209 35740 13243
rect 35682 13203 35740 13209
rect 37090 13200 37096 13252
rect 37148 13240 37154 13252
rect 37369 13243 37427 13249
rect 37369 13240 37381 13243
rect 37148 13212 37381 13240
rect 37148 13200 37154 13212
rect 37369 13209 37381 13212
rect 37415 13209 37427 13243
rect 37369 13203 37427 13209
rect 37553 13243 37611 13249
rect 37553 13209 37565 13243
rect 37599 13209 37611 13243
rect 38212 13240 38240 13271
rect 38562 13268 38568 13320
rect 38620 13308 38626 13320
rect 39853 13311 39911 13317
rect 39853 13308 39865 13311
rect 38620 13280 39865 13308
rect 38620 13268 38626 13280
rect 39853 13277 39865 13280
rect 39899 13277 39911 13311
rect 58158 13308 58164 13320
rect 58119 13280 58164 13308
rect 39853 13271 39911 13277
rect 58158 13268 58164 13280
rect 58216 13268 58222 13320
rect 39298 13240 39304 13252
rect 38212 13212 39304 13240
rect 37553 13203 37611 13209
rect 29914 13172 29920 13184
rect 27632 13144 29920 13172
rect 29914 13132 29920 13144
rect 29972 13132 29978 13184
rect 32582 13132 32588 13184
rect 32640 13172 32646 13184
rect 32769 13175 32827 13181
rect 32769 13172 32781 13175
rect 32640 13144 32781 13172
rect 32640 13132 32646 13144
rect 32769 13141 32781 13144
rect 32815 13141 32827 13175
rect 32769 13135 32827 13141
rect 37274 13132 37280 13184
rect 37332 13172 37338 13184
rect 37568 13172 37596 13203
rect 39298 13200 39304 13212
rect 39356 13200 39362 13252
rect 38838 13172 38844 13184
rect 37332 13144 37596 13172
rect 38799 13144 38844 13172
rect 37332 13132 37338 13144
rect 38838 13132 38844 13144
rect 38896 13132 38902 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 4985 12971 5043 12977
rect 4985 12937 4997 12971
rect 5031 12937 5043 12971
rect 4985 12931 5043 12937
rect 6733 12971 6791 12977
rect 6733 12937 6745 12971
rect 6779 12968 6791 12971
rect 7650 12968 7656 12980
rect 6779 12940 7656 12968
rect 6779 12937 6791 12940
rect 6733 12931 6791 12937
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 5000 12832 5028 12931
rect 7650 12928 7656 12940
rect 7708 12928 7714 12980
rect 10137 12971 10195 12977
rect 10137 12937 10149 12971
rect 10183 12968 10195 12971
rect 14093 12971 14151 12977
rect 10183 12940 12434 12968
rect 10183 12937 10195 12940
rect 10137 12931 10195 12937
rect 9585 12903 9643 12909
rect 9585 12869 9597 12903
rect 9631 12900 9643 12903
rect 10152 12900 10180 12931
rect 11054 12900 11060 12912
rect 9631 12872 10180 12900
rect 10967 12872 11060 12900
rect 9631 12869 9643 12872
rect 9585 12863 9643 12869
rect 11054 12860 11060 12872
rect 11112 12900 11118 12912
rect 12406 12900 12434 12940
rect 14093 12937 14105 12971
rect 14139 12968 14151 12971
rect 14826 12968 14832 12980
rect 14139 12940 14832 12968
rect 14139 12937 14151 12940
rect 14093 12931 14151 12937
rect 14826 12928 14832 12940
rect 14884 12928 14890 12980
rect 15746 12928 15752 12980
rect 15804 12968 15810 12980
rect 15841 12971 15899 12977
rect 15841 12968 15853 12971
rect 15804 12940 15853 12968
rect 15804 12928 15810 12940
rect 15841 12937 15853 12940
rect 15887 12968 15899 12971
rect 16022 12968 16028 12980
rect 15887 12940 16028 12968
rect 15887 12937 15899 12940
rect 15841 12931 15899 12937
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 18782 12968 18788 12980
rect 16776 12940 18788 12968
rect 16776 12900 16804 12940
rect 18782 12928 18788 12940
rect 18840 12928 18846 12980
rect 20073 12971 20131 12977
rect 20073 12937 20085 12971
rect 20119 12968 20131 12971
rect 21082 12968 21088 12980
rect 20119 12940 21088 12968
rect 20119 12937 20131 12940
rect 20073 12931 20131 12937
rect 21082 12928 21088 12940
rect 21140 12968 21146 12980
rect 23474 12968 23480 12980
rect 21140 12940 23480 12968
rect 21140 12928 21146 12940
rect 23474 12928 23480 12940
rect 23532 12928 23538 12980
rect 23750 12928 23756 12980
rect 23808 12968 23814 12980
rect 23937 12971 23995 12977
rect 23937 12968 23949 12971
rect 23808 12940 23949 12968
rect 23808 12928 23814 12940
rect 23937 12937 23949 12940
rect 23983 12937 23995 12971
rect 29730 12968 29736 12980
rect 29691 12940 29736 12968
rect 23937 12931 23995 12937
rect 29730 12928 29736 12940
rect 29788 12928 29794 12980
rect 30650 12968 30656 12980
rect 30611 12940 30656 12968
rect 30650 12928 30656 12940
rect 30708 12968 30714 12980
rect 30834 12968 30840 12980
rect 30708 12940 30840 12968
rect 30708 12928 30714 12940
rect 30834 12928 30840 12940
rect 30892 12928 30898 12980
rect 32217 12971 32275 12977
rect 32217 12937 32229 12971
rect 32263 12968 32275 12971
rect 32306 12968 32312 12980
rect 32263 12940 32312 12968
rect 32263 12937 32275 12940
rect 32217 12931 32275 12937
rect 32306 12928 32312 12940
rect 32364 12928 32370 12980
rect 33318 12968 33324 12980
rect 33279 12940 33324 12968
rect 33318 12928 33324 12940
rect 33376 12928 33382 12980
rect 35434 12968 35440 12980
rect 35395 12940 35440 12968
rect 35434 12928 35440 12940
rect 35492 12928 35498 12980
rect 35526 12928 35532 12980
rect 35584 12928 35590 12980
rect 37274 12928 37280 12980
rect 37332 12968 37338 12980
rect 39853 12971 39911 12977
rect 39853 12968 39865 12971
rect 37332 12940 39865 12968
rect 37332 12928 37338 12940
rect 39853 12937 39865 12940
rect 39899 12937 39911 12971
rect 39853 12931 39911 12937
rect 11112 12872 12296 12900
rect 12406 12872 16804 12900
rect 11112 12860 11118 12872
rect 5350 12832 5356 12844
rect 2547 12804 5028 12832
rect 5311 12804 5356 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 7834 12792 7840 12844
rect 7892 12832 7898 12844
rect 11072 12832 11100 12860
rect 11698 12832 11704 12844
rect 7892 12804 11100 12832
rect 11659 12804 11704 12832
rect 7892 12792 7898 12804
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12268 12841 12296 12872
rect 16850 12860 16856 12912
rect 16908 12900 16914 12912
rect 16908 12872 18368 12900
rect 16908 12860 16914 12872
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12832 12127 12835
rect 12253 12835 12311 12841
rect 12115 12804 12204 12832
rect 12115 12801 12127 12804
rect 12069 12795 12127 12801
rect 2682 12764 2688 12776
rect 2643 12736 2688 12764
rect 2682 12724 2688 12736
rect 2740 12724 2746 12776
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 3973 12767 4031 12773
rect 3973 12764 3985 12767
rect 2924 12736 3985 12764
rect 2924 12724 2930 12736
rect 3973 12733 3985 12736
rect 4019 12733 4031 12767
rect 3973 12727 4031 12733
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12764 4307 12767
rect 4614 12764 4620 12776
rect 4295 12736 4620 12764
rect 4295 12733 4307 12736
rect 4249 12727 4307 12733
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 5442 12764 5448 12776
rect 5403 12736 5448 12764
rect 5442 12724 5448 12736
rect 5500 12724 5506 12776
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 6822 12764 6828 12776
rect 6783 12736 6828 12764
rect 5537 12727 5595 12733
rect 4706 12656 4712 12708
rect 4764 12696 4770 12708
rect 5552 12696 5580 12727
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 4764 12668 5580 12696
rect 4764 12656 4770 12668
rect 5994 12656 6000 12708
rect 6052 12696 6058 12708
rect 6932 12696 6960 12727
rect 9674 12724 9680 12776
rect 9732 12764 9738 12776
rect 11885 12767 11943 12773
rect 11885 12764 11897 12767
rect 9732 12736 11897 12764
rect 9732 12724 9738 12736
rect 11885 12733 11897 12736
rect 11931 12733 11943 12767
rect 11885 12727 11943 12733
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12176 12764 12204 12804
rect 12253 12801 12265 12835
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 13170 12792 13176 12844
rect 13228 12832 13234 12844
rect 14277 12835 14335 12841
rect 14277 12832 14289 12835
rect 13228 12804 14289 12832
rect 13228 12792 13234 12804
rect 14277 12801 14289 12804
rect 14323 12801 14335 12835
rect 14277 12795 14335 12801
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12832 14519 12835
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14507 12804 14933 12832
rect 14507 12801 14519 12804
rect 14461 12795 14519 12801
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 15102 12832 15108 12844
rect 15063 12804 15108 12832
rect 14921 12795 14979 12801
rect 14936 12764 14964 12795
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 18046 12832 18052 12844
rect 18104 12841 18110 12844
rect 18340 12841 18368 12872
rect 18966 12860 18972 12912
rect 19024 12900 19030 12912
rect 19024 12872 19472 12900
rect 19024 12860 19030 12872
rect 18016 12804 18052 12832
rect 18046 12792 18052 12804
rect 18104 12795 18116 12841
rect 18325 12835 18383 12841
rect 18325 12801 18337 12835
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 18104 12792 18110 12795
rect 18690 12792 18696 12844
rect 18748 12832 18754 12844
rect 19061 12835 19119 12841
rect 19061 12832 19073 12835
rect 18748 12804 19073 12832
rect 18748 12792 18754 12804
rect 19061 12801 19073 12804
rect 19107 12801 19119 12835
rect 19061 12795 19119 12801
rect 19153 12835 19211 12841
rect 19153 12801 19165 12835
rect 19199 12801 19211 12835
rect 19153 12795 19211 12801
rect 16666 12764 16672 12776
rect 12032 12736 12077 12764
rect 12176 12736 12434 12764
rect 14936 12736 16672 12764
rect 12032 12724 12038 12736
rect 6052 12668 6960 12696
rect 12406 12696 12434 12736
rect 16666 12724 16672 12736
rect 16724 12724 16730 12776
rect 18782 12724 18788 12776
rect 18840 12764 18846 12776
rect 19168 12764 19196 12795
rect 19242 12792 19248 12844
rect 19300 12832 19306 12844
rect 19444 12841 19472 12872
rect 20622 12860 20628 12912
rect 20680 12900 20686 12912
rect 20806 12900 20812 12912
rect 20680 12872 20812 12900
rect 20680 12860 20686 12872
rect 20806 12860 20812 12872
rect 20864 12900 20870 12912
rect 20901 12903 20959 12909
rect 20901 12900 20913 12903
rect 20864 12872 20913 12900
rect 20864 12860 20870 12872
rect 20901 12869 20913 12872
rect 20947 12869 20959 12903
rect 26142 12900 26148 12912
rect 26103 12872 26148 12900
rect 20901 12863 20959 12869
rect 26142 12860 26148 12872
rect 26200 12860 26206 12912
rect 29362 12900 29368 12912
rect 29323 12872 29368 12900
rect 29362 12860 29368 12872
rect 29420 12860 29426 12912
rect 29546 12900 29552 12912
rect 29507 12872 29552 12900
rect 29546 12860 29552 12872
rect 29604 12860 29610 12912
rect 32324 12900 32352 12928
rect 32324 12872 33171 12900
rect 19429 12835 19487 12841
rect 19300 12804 19345 12832
rect 19300 12792 19306 12804
rect 19429 12801 19441 12835
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12832 19947 12835
rect 20070 12832 20076 12844
rect 19935 12804 20076 12832
rect 19935 12801 19947 12804
rect 19889 12795 19947 12801
rect 20070 12792 20076 12804
rect 20128 12792 20134 12844
rect 20717 12835 20775 12841
rect 20717 12801 20729 12835
rect 20763 12832 20775 12835
rect 21174 12832 21180 12844
rect 20763 12804 21180 12832
rect 20763 12801 20775 12804
rect 20717 12795 20775 12801
rect 21174 12792 21180 12804
rect 21232 12832 21238 12844
rect 21450 12832 21456 12844
rect 21232 12804 21456 12832
rect 21232 12792 21238 12804
rect 21450 12792 21456 12804
rect 21508 12792 21514 12844
rect 24489 12835 24547 12841
rect 24489 12801 24501 12835
rect 24535 12832 24547 12835
rect 26234 12832 26240 12844
rect 24535 12804 26240 12832
rect 24535 12801 24547 12804
rect 24489 12795 24547 12801
rect 26234 12792 26240 12804
rect 26292 12832 26298 12844
rect 26973 12835 27031 12841
rect 26973 12832 26985 12835
rect 26292 12804 26985 12832
rect 26292 12792 26298 12804
rect 26973 12801 26985 12804
rect 27019 12832 27031 12835
rect 27062 12832 27068 12844
rect 27019 12804 27068 12832
rect 27019 12801 27031 12804
rect 26973 12795 27031 12801
rect 27062 12792 27068 12804
rect 27120 12792 27126 12844
rect 32674 12832 32680 12844
rect 32635 12804 32680 12832
rect 32674 12792 32680 12804
rect 32732 12792 32738 12844
rect 32858 12832 32864 12844
rect 32819 12804 32864 12832
rect 32858 12792 32864 12804
rect 32916 12792 32922 12844
rect 32950 12792 32956 12844
rect 33008 12832 33014 12844
rect 33143 12841 33171 12872
rect 33091 12835 33171 12841
rect 33008 12804 33053 12832
rect 33008 12792 33014 12804
rect 33091 12801 33103 12835
rect 33137 12804 33171 12835
rect 35544 12832 35572 12928
rect 35618 12860 35624 12912
rect 35676 12900 35682 12912
rect 38740 12903 38798 12909
rect 35676 12872 36124 12900
rect 35676 12860 35682 12872
rect 35713 12835 35771 12841
rect 35713 12832 35725 12835
rect 35544 12804 35725 12832
rect 33137 12801 33149 12804
rect 33091 12795 33149 12801
rect 35636 12776 35664 12804
rect 35713 12801 35725 12804
rect 35759 12801 35771 12835
rect 35713 12795 35771 12801
rect 35805 12835 35863 12841
rect 35805 12801 35817 12835
rect 35851 12801 35863 12835
rect 35805 12795 35863 12801
rect 21634 12764 21640 12776
rect 18840 12736 19196 12764
rect 19260 12736 21640 12764
rect 18840 12724 18846 12736
rect 12805 12699 12863 12705
rect 12805 12696 12817 12699
rect 12406 12668 12817 12696
rect 6052 12656 6058 12668
rect 12805 12665 12817 12668
rect 12851 12696 12863 12699
rect 12851 12668 15608 12696
rect 12851 12665 12863 12668
rect 12805 12659 12863 12665
rect 2130 12588 2136 12640
rect 2188 12628 2194 12640
rect 2317 12631 2375 12637
rect 2317 12628 2329 12631
rect 2188 12600 2329 12628
rect 2188 12588 2194 12600
rect 2317 12597 2329 12600
rect 2363 12597 2375 12631
rect 6362 12628 6368 12640
rect 6323 12600 6368 12628
rect 2317 12591 2375 12597
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 8294 12628 8300 12640
rect 8255 12600 8300 12628
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 11514 12628 11520 12640
rect 11475 12600 11520 12628
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 15102 12588 15108 12640
rect 15160 12628 15166 12640
rect 15289 12631 15347 12637
rect 15289 12628 15301 12631
rect 15160 12600 15301 12628
rect 15160 12588 15166 12600
rect 15289 12597 15301 12600
rect 15335 12597 15347 12631
rect 15580 12628 15608 12668
rect 16390 12656 16396 12708
rect 16448 12696 16454 12708
rect 16945 12699 17003 12705
rect 16945 12696 16957 12699
rect 16448 12668 16957 12696
rect 16448 12656 16454 12668
rect 16945 12665 16957 12668
rect 16991 12665 17003 12699
rect 19260 12696 19288 12736
rect 21634 12724 21640 12736
rect 21692 12724 21698 12776
rect 21913 12767 21971 12773
rect 21913 12733 21925 12767
rect 21959 12764 21971 12767
rect 22186 12764 22192 12776
rect 21959 12736 22192 12764
rect 21959 12733 21971 12736
rect 21913 12727 21971 12733
rect 22186 12724 22192 12736
rect 22244 12764 22250 12776
rect 22465 12767 22523 12773
rect 22465 12764 22477 12767
rect 22244 12736 22477 12764
rect 22244 12724 22250 12736
rect 22465 12733 22477 12736
rect 22511 12764 22523 12767
rect 27338 12764 27344 12776
rect 22511 12736 27344 12764
rect 22511 12733 22523 12736
rect 22465 12727 22523 12733
rect 27338 12724 27344 12736
rect 27396 12724 27402 12776
rect 34057 12767 34115 12773
rect 34057 12733 34069 12767
rect 34103 12733 34115 12767
rect 34330 12764 34336 12776
rect 34291 12736 34336 12764
rect 34057 12727 34115 12733
rect 16945 12659 17003 12665
rect 18340 12668 19288 12696
rect 18340 12628 18368 12668
rect 15580 12600 18368 12628
rect 15289 12591 15347 12597
rect 18414 12588 18420 12640
rect 18472 12628 18478 12640
rect 18785 12631 18843 12637
rect 18785 12628 18797 12631
rect 18472 12600 18797 12628
rect 18472 12588 18478 12600
rect 18785 12597 18797 12600
rect 18831 12597 18843 12631
rect 18785 12591 18843 12597
rect 21085 12631 21143 12637
rect 21085 12597 21097 12631
rect 21131 12628 21143 12631
rect 21910 12628 21916 12640
rect 21131 12600 21916 12628
rect 21131 12597 21143 12600
rect 21085 12591 21143 12597
rect 21910 12588 21916 12600
rect 21968 12588 21974 12640
rect 25498 12588 25504 12640
rect 25556 12628 25562 12640
rect 33226 12628 33232 12640
rect 25556 12600 33232 12628
rect 25556 12588 25562 12600
rect 33226 12588 33232 12600
rect 33284 12628 33290 12640
rect 33870 12628 33876 12640
rect 33284 12600 33876 12628
rect 33284 12588 33290 12600
rect 33870 12588 33876 12600
rect 33928 12628 33934 12640
rect 34072 12628 34100 12727
rect 34330 12724 34336 12736
rect 34388 12724 34394 12776
rect 35618 12724 35624 12776
rect 35676 12724 35682 12776
rect 35820 12764 35848 12795
rect 35894 12792 35900 12844
rect 35952 12832 35958 12844
rect 36096 12841 36124 12872
rect 38740 12869 38752 12903
rect 38786 12900 38798 12903
rect 38838 12900 38844 12912
rect 38786 12872 38844 12900
rect 38786 12869 38798 12872
rect 38740 12863 38798 12869
rect 38838 12860 38844 12872
rect 38896 12860 38902 12912
rect 36081 12835 36139 12841
rect 35952 12804 35997 12832
rect 35952 12792 35958 12804
rect 36081 12801 36093 12835
rect 36127 12801 36139 12835
rect 37642 12832 37648 12844
rect 37603 12804 37648 12832
rect 36081 12795 36139 12801
rect 37642 12792 37648 12804
rect 37700 12792 37706 12844
rect 38102 12792 38108 12844
rect 38160 12832 38166 12844
rect 38473 12835 38531 12841
rect 38473 12832 38485 12835
rect 38160 12804 38485 12832
rect 38160 12792 38166 12804
rect 38473 12801 38485 12804
rect 38519 12801 38531 12835
rect 39574 12832 39580 12844
rect 38473 12795 38531 12801
rect 38580 12804 39580 12832
rect 35986 12764 35992 12776
rect 35820 12736 35992 12764
rect 35986 12724 35992 12736
rect 36044 12764 36050 12776
rect 38580 12764 38608 12804
rect 39574 12792 39580 12804
rect 39632 12792 39638 12844
rect 36044 12736 38608 12764
rect 36044 12724 36050 12736
rect 33928 12600 34100 12628
rect 33928 12588 33934 12600
rect 36446 12588 36452 12640
rect 36504 12628 36510 12640
rect 37090 12628 37096 12640
rect 36504 12600 37096 12628
rect 36504 12588 36510 12600
rect 37090 12588 37096 12600
rect 37148 12628 37154 12640
rect 37461 12631 37519 12637
rect 37461 12628 37473 12631
rect 37148 12600 37473 12628
rect 37148 12588 37154 12600
rect 37461 12597 37473 12600
rect 37507 12597 37519 12631
rect 37461 12591 37519 12597
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 6362 12424 6368 12436
rect 2700 12396 6368 12424
rect 2700 12229 2728 12396
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 9766 12424 9772 12436
rect 9723 12396 9772 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 10229 12427 10287 12433
rect 10229 12393 10241 12427
rect 10275 12424 10287 12427
rect 12526 12424 12532 12436
rect 10275 12396 12532 12424
rect 10275 12393 10287 12396
rect 10229 12387 10287 12393
rect 6270 12316 6276 12368
rect 6328 12356 6334 12368
rect 10244 12356 10272 12387
rect 12526 12384 12532 12396
rect 12584 12384 12590 12436
rect 13173 12427 13231 12433
rect 13173 12393 13185 12427
rect 13219 12424 13231 12427
rect 14090 12424 14096 12436
rect 13219 12396 14096 12424
rect 13219 12393 13231 12396
rect 13173 12387 13231 12393
rect 14090 12384 14096 12396
rect 14148 12424 14154 12436
rect 22370 12424 22376 12436
rect 14148 12396 22376 12424
rect 14148 12384 14154 12396
rect 22370 12384 22376 12396
rect 22428 12384 22434 12436
rect 22649 12427 22707 12433
rect 22649 12393 22661 12427
rect 22695 12424 22707 12427
rect 27890 12424 27896 12436
rect 22695 12396 27896 12424
rect 22695 12393 22707 12396
rect 22649 12387 22707 12393
rect 6328 12328 6684 12356
rect 6328 12316 6334 12328
rect 3786 12288 3792 12300
rect 3747 12260 3792 12288
rect 3786 12248 3792 12260
rect 3844 12248 3850 12300
rect 5350 12248 5356 12300
rect 5408 12288 5414 12300
rect 6656 12297 6684 12328
rect 9140 12328 10272 12356
rect 5813 12291 5871 12297
rect 5813 12288 5825 12291
rect 5408 12260 5825 12288
rect 5408 12248 5414 12260
rect 5813 12257 5825 12260
rect 5859 12257 5871 12291
rect 5813 12251 5871 12257
rect 6641 12291 6699 12297
rect 6641 12257 6653 12291
rect 6687 12257 6699 12291
rect 6641 12251 6699 12257
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12288 6791 12291
rect 7374 12288 7380 12300
rect 6779 12260 7380 12288
rect 6779 12257 6791 12260
rect 6733 12251 6791 12257
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7834 12288 7840 12300
rect 7795 12260 7840 12288
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 1857 12223 1915 12229
rect 1857 12189 1869 12223
rect 1903 12220 1915 12223
rect 2501 12223 2559 12229
rect 2501 12220 2513 12223
rect 1903 12192 2513 12220
rect 1903 12189 1915 12192
rect 1857 12183 1915 12189
rect 2501 12189 2513 12192
rect 2547 12189 2559 12223
rect 2501 12183 2559 12189
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12189 2743 12223
rect 2866 12220 2872 12232
rect 2827 12192 2872 12220
rect 2685 12183 2743 12189
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 6178 12180 6184 12232
rect 6236 12220 6242 12232
rect 6365 12223 6423 12229
rect 6365 12220 6377 12223
rect 6236 12192 6377 12220
rect 6236 12180 6242 12192
rect 6365 12189 6377 12192
rect 6411 12189 6423 12223
rect 6365 12183 6423 12189
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 6553 12223 6611 12229
rect 6553 12220 6565 12223
rect 6512 12192 6565 12220
rect 6512 12180 6518 12192
rect 6553 12189 6565 12192
rect 6599 12189 6611 12223
rect 6553 12183 6611 12189
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12220 6975 12223
rect 7006 12220 7012 12232
rect 6963 12192 7012 12220
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 7561 12223 7619 12229
rect 7561 12189 7573 12223
rect 7607 12189 7619 12223
rect 7852 12220 7880 12248
rect 9140 12229 9168 12328
rect 13814 12316 13820 12368
rect 13872 12356 13878 12368
rect 15010 12356 15016 12368
rect 13872 12328 15016 12356
rect 13872 12316 13878 12328
rect 15010 12316 15016 12328
rect 15068 12356 15074 12368
rect 15068 12328 15332 12356
rect 15068 12316 15074 12328
rect 15194 12288 15200 12300
rect 14936 12260 15200 12288
rect 8929 12223 8987 12229
rect 8929 12220 8941 12223
rect 7852 12192 8941 12220
rect 7561 12183 7619 12189
rect 8929 12189 8941 12192
rect 8975 12189 8987 12223
rect 8929 12183 8987 12189
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12189 9183 12223
rect 9125 12183 9183 12189
rect 9217 12223 9275 12229
rect 9217 12189 9229 12223
rect 9263 12189 9275 12223
rect 9217 12183 9275 12189
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9493 12223 9551 12229
rect 9493 12189 9505 12223
rect 9539 12220 9551 12223
rect 10686 12220 10692 12232
rect 9539 12192 10692 12220
rect 9539 12189 9551 12192
rect 9493 12183 9551 12189
rect 4034 12155 4092 12161
rect 4034 12152 4046 12155
rect 2056 12124 4046 12152
rect 2056 12093 2084 12124
rect 4034 12121 4046 12124
rect 4080 12121 4092 12155
rect 4034 12115 4092 12121
rect 4614 12112 4620 12164
rect 4672 12152 4678 12164
rect 7576 12152 7604 12183
rect 4672 12124 6684 12152
rect 4672 12112 4678 12124
rect 2041 12087 2099 12093
rect 2041 12053 2053 12087
rect 2087 12053 2099 12087
rect 2041 12047 2099 12053
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 5534 12084 5540 12096
rect 5215 12056 5540 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5534 12044 5540 12056
rect 5592 12084 5598 12096
rect 6546 12084 6552 12096
rect 5592 12056 6552 12084
rect 5592 12044 5598 12056
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 6656 12084 6684 12124
rect 6932 12124 7604 12152
rect 6932 12084 6960 12124
rect 7098 12084 7104 12096
rect 6656 12056 6960 12084
rect 7059 12056 7104 12084
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 7576 12084 7604 12124
rect 7650 12112 7656 12164
rect 7708 12152 7714 12164
rect 9232 12152 9260 12183
rect 7708 12124 9260 12152
rect 9324 12152 9352 12183
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 11514 12180 11520 12232
rect 11572 12220 11578 12232
rect 12262 12223 12320 12229
rect 12262 12220 12274 12223
rect 11572 12192 12274 12220
rect 11572 12180 11578 12192
rect 12262 12189 12274 12192
rect 12308 12189 12320 12223
rect 12526 12220 12532 12232
rect 12487 12192 12532 12220
rect 12262 12183 12320 12189
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 14936 12229 14964 12260
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 15304 12288 15332 12328
rect 16666 12316 16672 12368
rect 16724 12356 16730 12368
rect 20162 12356 20168 12368
rect 16724 12328 20168 12356
rect 16724 12316 16730 12328
rect 20162 12316 20168 12328
rect 20220 12316 20226 12368
rect 21008 12328 21864 12356
rect 21008 12300 21036 12328
rect 16114 12288 16120 12300
rect 15304 12260 16120 12288
rect 12989 12223 13047 12229
rect 12989 12189 13001 12223
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 15013 12223 15071 12229
rect 15013 12189 15025 12223
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 9766 12152 9772 12164
rect 9324 12124 9772 12152
rect 7708 12112 7714 12124
rect 9766 12112 9772 12124
rect 9824 12112 9830 12164
rect 12066 12152 12072 12164
rect 10520 12124 12072 12152
rect 10520 12084 10548 12124
rect 12066 12112 12072 12124
rect 12124 12112 12130 12164
rect 12342 12112 12348 12164
rect 12400 12152 12406 12164
rect 13004 12152 13032 12183
rect 12400 12124 13032 12152
rect 12400 12112 12406 12124
rect 14550 12112 14556 12164
rect 14608 12152 14614 12164
rect 15028 12152 15056 12183
rect 15102 12180 15108 12232
rect 15160 12220 15166 12232
rect 15304 12229 15332 12260
rect 16114 12248 16120 12260
rect 16172 12248 16178 12300
rect 17126 12248 17132 12300
rect 17184 12288 17190 12300
rect 20990 12288 20996 12300
rect 17184 12260 19472 12288
rect 20951 12260 20996 12288
rect 17184 12248 17190 12260
rect 15289 12223 15347 12229
rect 15160 12192 15205 12220
rect 15160 12180 15166 12192
rect 15289 12189 15301 12223
rect 15335 12189 15347 12223
rect 16022 12220 16028 12232
rect 15289 12183 15347 12189
rect 15396 12192 16028 12220
rect 14608 12124 15056 12152
rect 14608 12112 14614 12124
rect 7576 12056 10548 12084
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 11149 12087 11207 12093
rect 11149 12084 11161 12087
rect 10652 12056 11161 12084
rect 10652 12044 10658 12056
rect 11149 12053 11161 12056
rect 11195 12084 11207 12087
rect 11698 12084 11704 12096
rect 11195 12056 11704 12084
rect 11195 12053 11207 12056
rect 11149 12047 11207 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 13262 12044 13268 12096
rect 13320 12084 13326 12096
rect 14182 12084 14188 12096
rect 13320 12056 14188 12084
rect 13320 12044 13326 12056
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 14642 12084 14648 12096
rect 14603 12056 14648 12084
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 15028 12084 15056 12124
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 15396 12152 15424 12192
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 18138 12180 18144 12232
rect 18196 12214 18202 12232
rect 18305 12223 18363 12229
rect 18305 12220 18317 12223
rect 18248 12214 18317 12220
rect 18196 12192 18317 12214
rect 18196 12186 18276 12192
rect 18305 12189 18317 12192
rect 18351 12189 18363 12223
rect 18196 12180 18202 12186
rect 18305 12183 18363 12189
rect 18417 12217 18475 12223
rect 18417 12183 18429 12217
rect 18463 12183 18475 12217
rect 18417 12177 18475 12183
rect 18506 12180 18512 12232
rect 18564 12220 18570 12232
rect 18693 12223 18751 12229
rect 18564 12192 18609 12220
rect 18564 12180 18570 12192
rect 18693 12189 18705 12223
rect 18739 12220 18751 12223
rect 19058 12220 19064 12232
rect 18739 12192 19064 12220
rect 18739 12189 18751 12192
rect 18693 12183 18751 12189
rect 19058 12180 19064 12192
rect 19116 12180 19122 12232
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 19334 12220 19340 12232
rect 19291 12192 19340 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 19334 12180 19340 12192
rect 19392 12180 19398 12232
rect 19444 12229 19472 12260
rect 20990 12248 20996 12260
rect 21048 12248 21054 12300
rect 21450 12288 21456 12300
rect 21411 12260 21456 12288
rect 21450 12248 21456 12260
rect 21508 12248 21514 12300
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12189 19487 12223
rect 20717 12223 20775 12229
rect 20717 12220 20729 12223
rect 19429 12183 19487 12189
rect 19516 12192 20729 12220
rect 15252 12124 15424 12152
rect 15252 12112 15258 12124
rect 15746 12112 15752 12164
rect 15804 12152 15810 12164
rect 15841 12155 15899 12161
rect 15841 12152 15853 12155
rect 15804 12124 15853 12152
rect 15804 12112 15810 12124
rect 15841 12121 15853 12124
rect 15887 12152 15899 12155
rect 16574 12152 16580 12164
rect 15887 12124 16580 12152
rect 15887 12121 15899 12124
rect 15841 12115 15899 12121
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 18046 12152 18052 12164
rect 16684 12124 17264 12152
rect 18007 12124 18052 12152
rect 16684 12084 16712 12124
rect 15028 12056 16712 12084
rect 16850 12044 16856 12096
rect 16908 12084 16914 12096
rect 17129 12087 17187 12093
rect 17129 12084 17141 12087
rect 16908 12056 17141 12084
rect 16908 12044 16914 12056
rect 17129 12053 17141 12056
rect 17175 12053 17187 12087
rect 17236 12084 17264 12124
rect 18046 12112 18052 12124
rect 18104 12112 18110 12164
rect 18432 12084 18460 12177
rect 18782 12112 18788 12164
rect 18840 12152 18846 12164
rect 19516 12152 19544 12192
rect 20717 12189 20729 12192
rect 20763 12189 20775 12223
rect 21709 12223 21767 12229
rect 21836 12226 21864 12328
rect 22002 12316 22008 12368
rect 22060 12356 22066 12368
rect 22554 12356 22560 12368
rect 22060 12328 22560 12356
rect 22060 12316 22066 12328
rect 22554 12316 22560 12328
rect 22612 12316 22618 12368
rect 21709 12220 21721 12223
rect 21698 12214 21721 12220
rect 20717 12183 20775 12189
rect 21652 12189 21721 12214
rect 21755 12189 21767 12223
rect 21652 12186 21767 12189
rect 18840 12124 19544 12152
rect 19613 12155 19671 12161
rect 18840 12112 18846 12124
rect 19613 12121 19625 12155
rect 19659 12152 19671 12155
rect 20162 12152 20168 12164
rect 19659 12124 20168 12152
rect 19659 12121 19671 12124
rect 19613 12115 19671 12121
rect 20162 12112 20168 12124
rect 20220 12112 20226 12164
rect 21652 12152 21680 12186
rect 21709 12183 21767 12186
rect 21818 12220 21876 12226
rect 21818 12186 21830 12220
rect 21864 12186 21876 12220
rect 21818 12180 21876 12186
rect 21910 12180 21916 12232
rect 21968 12229 21974 12232
rect 21968 12220 21976 12229
rect 21968 12192 22013 12220
rect 21968 12183 21976 12192
rect 21968 12180 21974 12183
rect 22094 12180 22100 12232
rect 22152 12220 22158 12232
rect 22664 12220 22692 12387
rect 27890 12384 27896 12396
rect 27948 12384 27954 12436
rect 32858 12424 32864 12436
rect 32819 12396 32864 12424
rect 32858 12384 32864 12396
rect 32916 12384 32922 12436
rect 33870 12424 33876 12436
rect 33831 12396 33876 12424
rect 33870 12384 33876 12396
rect 33928 12384 33934 12436
rect 35618 12384 35624 12436
rect 35676 12424 35682 12436
rect 35989 12427 36047 12433
rect 35989 12424 36001 12427
rect 35676 12396 36001 12424
rect 35676 12384 35682 12396
rect 35989 12393 36001 12396
rect 36035 12393 36047 12427
rect 35989 12387 36047 12393
rect 35529 12359 35587 12365
rect 35529 12325 35541 12359
rect 35575 12356 35587 12359
rect 36998 12356 37004 12368
rect 35575 12328 37004 12356
rect 35575 12325 35587 12328
rect 35529 12319 35587 12325
rect 36998 12316 37004 12328
rect 37056 12316 37062 12368
rect 38562 12316 38568 12368
rect 38620 12316 38626 12368
rect 30098 12288 30104 12300
rect 30011 12260 30104 12288
rect 30098 12248 30104 12260
rect 30156 12288 30162 12300
rect 30156 12260 30972 12288
rect 30156 12248 30162 12260
rect 25038 12220 25044 12232
rect 22152 12192 22692 12220
rect 24999 12192 25044 12220
rect 22152 12180 22158 12192
rect 25038 12180 25044 12192
rect 25096 12220 25102 12232
rect 26142 12220 26148 12232
rect 25096 12192 26148 12220
rect 25096 12180 25102 12192
rect 26142 12180 26148 12192
rect 26200 12180 26206 12232
rect 28074 12220 28080 12232
rect 26252 12192 28080 12220
rect 22186 12152 22192 12164
rect 21652 12124 22192 12152
rect 22186 12112 22192 12124
rect 22244 12112 22250 12164
rect 25130 12112 25136 12164
rect 25188 12152 25194 12164
rect 25286 12155 25344 12161
rect 25286 12152 25298 12155
rect 25188 12124 25298 12152
rect 25188 12112 25194 12124
rect 25286 12121 25298 12124
rect 25332 12121 25344 12155
rect 26252 12152 26280 12192
rect 28074 12180 28080 12192
rect 28132 12220 28138 12232
rect 28353 12223 28411 12229
rect 28353 12220 28365 12223
rect 28132 12192 28365 12220
rect 28132 12180 28138 12192
rect 28353 12189 28365 12192
rect 28399 12189 28411 12223
rect 30558 12220 30564 12232
rect 30519 12192 30564 12220
rect 28353 12183 28411 12189
rect 30558 12180 30564 12192
rect 30616 12180 30622 12232
rect 30742 12220 30748 12232
rect 30703 12192 30748 12220
rect 30742 12180 30748 12192
rect 30800 12180 30806 12232
rect 30944 12229 30972 12260
rect 31018 12248 31024 12300
rect 31076 12288 31082 12300
rect 38580 12288 38608 12316
rect 31076 12260 38608 12288
rect 31076 12248 31082 12260
rect 39022 12248 39028 12300
rect 39080 12288 39086 12300
rect 40129 12291 40187 12297
rect 40129 12288 40141 12291
rect 39080 12260 40141 12288
rect 39080 12248 39086 12260
rect 40129 12257 40141 12260
rect 40175 12257 40187 12291
rect 40129 12251 40187 12257
rect 30837 12223 30895 12229
rect 30837 12189 30849 12223
rect 30883 12189 30895 12223
rect 30837 12183 30895 12189
rect 30929 12223 30987 12229
rect 30929 12189 30941 12223
rect 30975 12189 30987 12223
rect 31202 12220 31208 12232
rect 30929 12183 30987 12189
rect 31036 12192 31208 12220
rect 25286 12115 25344 12121
rect 25976 12124 26280 12152
rect 27525 12155 27583 12161
rect 18800 12084 18828 12112
rect 17236 12056 18828 12084
rect 17129 12047 17187 12053
rect 19058 12044 19064 12096
rect 19116 12084 19122 12096
rect 25976 12084 26004 12124
rect 27525 12121 27537 12155
rect 27571 12152 27583 12155
rect 28166 12152 28172 12164
rect 27571 12124 28172 12152
rect 27571 12121 27583 12124
rect 27525 12115 27583 12121
rect 28166 12112 28172 12124
rect 28224 12112 28230 12164
rect 30852 12152 30880 12183
rect 31036 12152 31064 12192
rect 31202 12180 31208 12192
rect 31260 12220 31266 12232
rect 32950 12220 32956 12232
rect 31260 12192 32956 12220
rect 31260 12180 31266 12192
rect 32950 12180 32956 12192
rect 33008 12180 33014 12232
rect 34330 12180 34336 12232
rect 34388 12220 34394 12232
rect 35345 12223 35403 12229
rect 35345 12220 35357 12223
rect 34388 12192 35357 12220
rect 34388 12180 34394 12192
rect 35345 12189 35357 12192
rect 35391 12189 35403 12223
rect 38286 12220 38292 12232
rect 38247 12192 38292 12220
rect 35345 12183 35403 12189
rect 38286 12180 38292 12192
rect 38344 12180 38350 12232
rect 38565 12223 38623 12229
rect 38565 12189 38577 12223
rect 38611 12220 38623 12223
rect 39482 12220 39488 12232
rect 38611 12192 39488 12220
rect 38611 12189 38623 12192
rect 38565 12183 38623 12189
rect 39482 12180 39488 12192
rect 39540 12180 39546 12232
rect 39758 12180 39764 12232
rect 39816 12220 39822 12232
rect 39853 12223 39911 12229
rect 39853 12220 39865 12223
rect 39816 12192 39865 12220
rect 39816 12180 39822 12192
rect 39853 12189 39865 12192
rect 39899 12189 39911 12223
rect 39853 12183 39911 12189
rect 32493 12155 32551 12161
rect 32493 12152 32505 12155
rect 30852 12124 31064 12152
rect 31128 12124 32505 12152
rect 19116 12056 26004 12084
rect 19116 12044 19122 12056
rect 26050 12044 26056 12096
rect 26108 12084 26114 12096
rect 26421 12087 26479 12093
rect 26421 12084 26433 12087
rect 26108 12056 26433 12084
rect 26108 12044 26114 12056
rect 26421 12053 26433 12056
rect 26467 12053 26479 12087
rect 27430 12084 27436 12096
rect 27391 12056 27436 12084
rect 26421 12047 26479 12053
rect 27430 12044 27436 12056
rect 27488 12044 27494 12096
rect 30190 12044 30196 12096
rect 30248 12084 30254 12096
rect 31128 12084 31156 12124
rect 32493 12121 32505 12124
rect 32539 12121 32551 12155
rect 32493 12115 32551 12121
rect 32582 12112 32588 12164
rect 32640 12152 32646 12164
rect 32677 12155 32735 12161
rect 32677 12152 32689 12155
rect 32640 12124 32689 12152
rect 32640 12112 32646 12124
rect 32677 12121 32689 12124
rect 32723 12121 32735 12155
rect 32677 12115 32735 12121
rect 30248 12056 31156 12084
rect 31205 12087 31263 12093
rect 30248 12044 30254 12056
rect 31205 12053 31217 12087
rect 31251 12084 31263 12087
rect 31386 12084 31392 12096
rect 31251 12056 31392 12084
rect 31251 12053 31263 12056
rect 31205 12047 31263 12053
rect 31386 12044 31392 12056
rect 31444 12044 31450 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11880 5871 11883
rect 7650 11880 7656 11892
rect 5859 11852 7656 11880
rect 5859 11849 5871 11852
rect 5813 11843 5871 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 14734 11880 14740 11892
rect 14139 11852 14740 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 17126 11880 17132 11892
rect 17087 11852 17132 11880
rect 17126 11840 17132 11852
rect 17184 11840 17190 11892
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 19889 11883 19947 11889
rect 17368 11852 18644 11880
rect 17368 11840 17374 11852
rect 3786 11812 3792 11824
rect 2792 11784 3792 11812
rect 2130 11744 2136 11756
rect 2091 11716 2136 11744
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 2792 11753 2820 11784
rect 3786 11772 3792 11784
rect 3844 11772 3850 11824
rect 6178 11772 6184 11824
rect 6236 11812 6242 11824
rect 6825 11815 6883 11821
rect 6825 11812 6837 11815
rect 6236 11784 6837 11812
rect 6236 11772 6242 11784
rect 6825 11781 6837 11784
rect 6871 11781 6883 11815
rect 6825 11775 6883 11781
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11713 2835 11747
rect 3033 11747 3091 11753
rect 3033 11744 3045 11747
rect 2777 11707 2835 11713
rect 2884 11716 3045 11744
rect 2884 11676 2912 11716
rect 3033 11713 3045 11716
rect 3079 11713 3091 11747
rect 5534 11744 5540 11756
rect 5495 11716 5540 11744
rect 3033 11707 3091 11713
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 2332 11648 2912 11676
rect 5169 11679 5227 11685
rect 2332 11617 2360 11648
rect 5169 11645 5181 11679
rect 5215 11676 5227 11679
rect 5258 11676 5264 11688
rect 5215 11648 5264 11676
rect 5215 11645 5227 11648
rect 5169 11639 5227 11645
rect 5258 11636 5264 11648
rect 5316 11636 5322 11688
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11676 5687 11679
rect 6454 11676 6460 11688
rect 5675 11648 6460 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 6454 11636 6460 11648
rect 6512 11636 6518 11688
rect 6840 11676 6868 11775
rect 7098 11772 7104 11824
rect 7156 11812 7162 11824
rect 8490 11815 8548 11821
rect 8490 11812 8502 11815
rect 7156 11784 8502 11812
rect 7156 11772 7162 11784
rect 8490 11781 8502 11784
rect 8536 11781 8548 11815
rect 8490 11775 8548 11781
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 16850 11812 16856 11824
rect 12584 11784 16856 11812
rect 12584 11772 12590 11784
rect 8754 11744 8760 11756
rect 8715 11716 8760 11744
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 12066 11744 12072 11756
rect 12027 11716 12072 11744
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 13262 11744 13268 11756
rect 13223 11716 13268 11744
rect 13262 11704 13268 11716
rect 13320 11704 13326 11756
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11713 13415 11747
rect 13357 11707 13415 11713
rect 7098 11676 7104 11688
rect 6840 11648 7104 11676
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 12342 11676 12348 11688
rect 12303 11648 12348 11676
rect 12342 11636 12348 11648
rect 12400 11636 12406 11688
rect 13372 11676 13400 11707
rect 13446 11704 13452 11756
rect 13504 11744 13510 11756
rect 13633 11747 13691 11753
rect 13504 11716 13549 11744
rect 13504 11704 13510 11716
rect 13633 11713 13645 11747
rect 13679 11744 13691 11747
rect 13814 11744 13820 11756
rect 13679 11716 13820 11744
rect 13679 11713 13691 11716
rect 13633 11707 13691 11713
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 15488 11753 15516 11784
rect 16850 11772 16856 11784
rect 16908 11812 16914 11824
rect 18616 11812 18644 11852
rect 19889 11849 19901 11883
rect 19935 11880 19947 11883
rect 20806 11880 20812 11892
rect 19935 11852 20812 11880
rect 19935 11849 19947 11852
rect 19889 11843 19947 11849
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 23293 11883 23351 11889
rect 23293 11880 23305 11883
rect 20916 11852 23305 11880
rect 20916 11812 20944 11852
rect 23293 11849 23305 11852
rect 23339 11880 23351 11883
rect 23842 11880 23848 11892
rect 23339 11852 23848 11880
rect 23339 11849 23351 11852
rect 23293 11843 23351 11849
rect 23842 11840 23848 11852
rect 23900 11840 23906 11892
rect 24486 11840 24492 11892
rect 24544 11880 24550 11892
rect 25130 11880 25136 11892
rect 24544 11852 24716 11880
rect 25091 11852 25136 11880
rect 24544 11840 24550 11852
rect 16908 11784 18552 11812
rect 18616 11784 20944 11812
rect 21024 11815 21082 11821
rect 16908 11772 16914 11784
rect 15206 11747 15264 11753
rect 15206 11744 15218 11747
rect 14700 11716 15218 11744
rect 14700 11704 14706 11716
rect 15206 11713 15218 11716
rect 15252 11713 15264 11747
rect 15206 11707 15264 11713
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 18253 11747 18311 11753
rect 18253 11713 18265 11747
rect 18299 11744 18311 11747
rect 18414 11744 18420 11756
rect 18299 11716 18420 11744
rect 18299 11713 18311 11716
rect 18253 11707 18311 11713
rect 18414 11704 18420 11716
rect 18472 11704 18478 11756
rect 18524 11753 18552 11784
rect 21024 11781 21036 11815
rect 21070 11812 21082 11815
rect 21450 11812 21456 11824
rect 21070 11784 21456 11812
rect 21070 11781 21082 11784
rect 21024 11775 21082 11781
rect 21450 11772 21456 11784
rect 21508 11772 21514 11824
rect 23474 11772 23480 11824
rect 23532 11812 23538 11824
rect 24581 11815 24639 11821
rect 24581 11812 24593 11815
rect 23532 11784 24593 11812
rect 23532 11772 23538 11784
rect 24581 11781 24593 11784
rect 24627 11781 24639 11815
rect 24688 11812 24716 11852
rect 25130 11840 25136 11852
rect 25188 11840 25194 11892
rect 27890 11840 27896 11892
rect 27948 11880 27954 11892
rect 28261 11883 28319 11889
rect 28261 11880 28273 11883
rect 27948 11852 28273 11880
rect 27948 11840 27954 11852
rect 28261 11849 28273 11852
rect 28307 11849 28319 11883
rect 28261 11843 28319 11849
rect 30469 11883 30527 11889
rect 30469 11849 30481 11883
rect 30515 11880 30527 11883
rect 30742 11880 30748 11892
rect 30515 11852 30748 11880
rect 30515 11849 30527 11852
rect 30469 11843 30527 11849
rect 30742 11840 30748 11852
rect 30800 11840 30806 11892
rect 30852 11852 32996 11880
rect 26142 11812 26148 11824
rect 24688 11784 26148 11812
rect 24581 11775 24639 11781
rect 18509 11747 18567 11753
rect 18509 11713 18521 11747
rect 18555 11713 18567 11747
rect 19242 11744 19248 11756
rect 19203 11716 19248 11744
rect 18509 11707 18567 11713
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 22002 11744 22008 11756
rect 19352 11716 22008 11744
rect 14458 11676 14464 11688
rect 13372 11648 14464 11676
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 2317 11611 2375 11617
rect 2317 11577 2329 11611
rect 2363 11577 2375 11611
rect 2317 11571 2375 11577
rect 6730 11568 6736 11620
rect 6788 11608 6794 11620
rect 7006 11608 7012 11620
rect 6788 11580 7012 11608
rect 6788 11568 6794 11580
rect 7006 11568 7012 11580
rect 7064 11608 7070 11620
rect 7377 11611 7435 11617
rect 7377 11608 7389 11611
rect 7064 11580 7389 11608
rect 7064 11568 7070 11580
rect 7377 11577 7389 11580
rect 7423 11577 7435 11611
rect 7377 11571 7435 11577
rect 10870 11568 10876 11620
rect 10928 11608 10934 11620
rect 19352 11608 19380 11716
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 22186 11744 22192 11756
rect 22147 11716 22192 11744
rect 22186 11704 22192 11716
rect 22244 11704 22250 11756
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11713 22339 11747
rect 22281 11707 22339 11713
rect 21269 11679 21327 11685
rect 21269 11645 21281 11679
rect 21315 11676 21327 11679
rect 21634 11676 21640 11688
rect 21315 11648 21640 11676
rect 21315 11645 21327 11648
rect 21269 11639 21327 11645
rect 21634 11636 21640 11648
rect 21692 11636 21698 11688
rect 22296 11608 22324 11707
rect 22370 11704 22376 11756
rect 22428 11744 22434 11756
rect 22428 11716 22473 11744
rect 22428 11704 22434 11716
rect 22554 11704 22560 11756
rect 22612 11744 22618 11756
rect 24596 11744 24624 11775
rect 25516 11753 25544 11784
rect 26142 11772 26148 11784
rect 26200 11772 26206 11824
rect 28166 11812 28172 11824
rect 28079 11784 28172 11812
rect 25409 11747 25467 11753
rect 25409 11744 25421 11747
rect 22612 11716 22705 11744
rect 24596 11716 25421 11744
rect 22612 11704 22618 11716
rect 25409 11713 25421 11716
rect 25455 11713 25467 11747
rect 25409 11707 25467 11713
rect 25501 11747 25559 11753
rect 25501 11713 25513 11747
rect 25547 11713 25559 11747
rect 25501 11707 25559 11713
rect 25590 11704 25596 11756
rect 25648 11744 25654 11756
rect 25777 11747 25835 11753
rect 25648 11716 25693 11744
rect 25648 11704 25654 11716
rect 25777 11713 25789 11747
rect 25823 11744 25835 11747
rect 27430 11744 27436 11756
rect 25823 11716 27436 11744
rect 25823 11713 25835 11716
rect 25777 11707 25835 11713
rect 22572 11676 22600 11704
rect 25792 11676 25820 11707
rect 27430 11704 27436 11716
rect 27488 11704 27494 11756
rect 28092 11753 28120 11784
rect 28166 11772 28172 11784
rect 28224 11812 28230 11824
rect 30852 11812 30880 11852
rect 28224 11784 30880 11812
rect 28224 11772 28230 11784
rect 28077 11747 28135 11753
rect 28077 11713 28089 11747
rect 28123 11713 28135 11747
rect 28077 11707 28135 11713
rect 30101 11747 30159 11753
rect 30101 11713 30113 11747
rect 30147 11713 30159 11747
rect 30282 11744 30288 11756
rect 30243 11716 30288 11744
rect 30101 11707 30159 11713
rect 22572 11648 25820 11676
rect 30116 11676 30144 11707
rect 30282 11704 30288 11716
rect 30340 11704 30346 11756
rect 30558 11704 30564 11756
rect 30616 11744 30622 11756
rect 30929 11747 30987 11753
rect 30929 11744 30941 11747
rect 30616 11716 30941 11744
rect 30616 11704 30622 11716
rect 30929 11713 30941 11716
rect 30975 11713 30987 11747
rect 31110 11744 31116 11756
rect 31071 11716 31116 11744
rect 30929 11707 30987 11713
rect 30190 11676 30196 11688
rect 30116 11648 30196 11676
rect 30190 11636 30196 11648
rect 30248 11636 30254 11688
rect 30944 11676 30972 11707
rect 31110 11704 31116 11716
rect 31168 11704 31174 11756
rect 31202 11704 31208 11756
rect 31260 11744 31266 11756
rect 31343 11747 31401 11753
rect 31260 11716 31305 11744
rect 31260 11704 31266 11716
rect 31343 11713 31355 11747
rect 31389 11744 31401 11747
rect 31478 11744 31484 11756
rect 31389 11716 31484 11744
rect 31389 11713 31401 11716
rect 31343 11707 31401 11713
rect 31478 11704 31484 11716
rect 31536 11744 31542 11756
rect 31938 11744 31944 11756
rect 31536 11716 31944 11744
rect 31536 11704 31542 11716
rect 31938 11704 31944 11716
rect 31996 11704 32002 11756
rect 32968 11753 32996 11852
rect 34422 11840 34428 11892
rect 34480 11880 34486 11892
rect 35253 11883 35311 11889
rect 35253 11880 35265 11883
rect 34480 11852 35265 11880
rect 34480 11840 34486 11852
rect 35253 11849 35265 11852
rect 35299 11849 35311 11883
rect 35253 11843 35311 11849
rect 39850 11840 39856 11892
rect 39908 11880 39914 11892
rect 39945 11883 40003 11889
rect 39945 11880 39957 11883
rect 39908 11852 39957 11880
rect 39908 11840 39914 11852
rect 39945 11849 39957 11852
rect 39991 11880 40003 11883
rect 39991 11852 40632 11880
rect 39991 11849 40003 11852
rect 39945 11843 40003 11849
rect 35529 11815 35587 11821
rect 35529 11781 35541 11815
rect 35575 11812 35587 11815
rect 36630 11812 36636 11824
rect 35575 11784 36636 11812
rect 35575 11781 35587 11784
rect 35529 11775 35587 11781
rect 36630 11772 36636 11784
rect 36688 11772 36694 11824
rect 38286 11772 38292 11824
rect 38344 11812 38350 11824
rect 40604 11821 40632 11852
rect 40405 11815 40463 11821
rect 40405 11812 40417 11815
rect 38344 11784 40417 11812
rect 38344 11772 38350 11784
rect 40405 11781 40417 11784
rect 40451 11781 40463 11815
rect 40405 11775 40463 11781
rect 40589 11815 40647 11821
rect 40589 11781 40601 11815
rect 40635 11781 40647 11815
rect 40589 11775 40647 11781
rect 32953 11747 33011 11753
rect 32953 11713 32965 11747
rect 32999 11744 33011 11747
rect 34330 11744 34336 11756
rect 32999 11716 34336 11744
rect 32999 11713 33011 11716
rect 32953 11707 33011 11713
rect 34330 11704 34336 11716
rect 34388 11704 34394 11756
rect 34790 11704 34796 11756
rect 34848 11744 34854 11756
rect 35437 11747 35495 11753
rect 35437 11744 35449 11747
rect 34848 11716 35449 11744
rect 34848 11704 34854 11716
rect 35437 11713 35449 11716
rect 35483 11713 35495 11747
rect 35437 11707 35495 11713
rect 35621 11747 35679 11753
rect 35621 11713 35633 11747
rect 35667 11713 35679 11747
rect 35802 11744 35808 11756
rect 35763 11716 35808 11744
rect 35621 11707 35679 11713
rect 32122 11676 32128 11688
rect 30944 11648 32128 11676
rect 32122 11636 32128 11648
rect 32180 11676 32186 11688
rect 32674 11676 32680 11688
rect 32180 11648 32680 11676
rect 32180 11636 32186 11648
rect 32674 11636 32680 11648
rect 32732 11636 32738 11688
rect 35636 11676 35664 11707
rect 35802 11704 35808 11716
rect 35860 11704 35866 11756
rect 38654 11704 38660 11756
rect 38712 11744 38718 11756
rect 38821 11747 38879 11753
rect 38821 11744 38833 11747
rect 38712 11716 38833 11744
rect 38712 11704 38718 11716
rect 38821 11713 38833 11716
rect 38867 11713 38879 11747
rect 38821 11707 38879 11713
rect 35710 11676 35716 11688
rect 35452 11648 35716 11676
rect 35452 11620 35480 11648
rect 35710 11636 35716 11648
rect 35768 11636 35774 11688
rect 38562 11676 38568 11688
rect 38523 11648 38568 11676
rect 38562 11636 38568 11648
rect 38620 11636 38626 11688
rect 24486 11608 24492 11620
rect 10928 11580 14596 11608
rect 10928 11568 10934 11580
rect 4157 11543 4215 11549
rect 4157 11509 4169 11543
rect 4203 11540 4215 11543
rect 4890 11540 4896 11552
rect 4203 11512 4896 11540
rect 4203 11509 4215 11512
rect 4157 11503 4215 11509
rect 4890 11500 4896 11512
rect 4948 11540 4954 11552
rect 5442 11540 5448 11552
rect 4948 11512 5448 11540
rect 4948 11500 4954 11512
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 12986 11540 12992 11552
rect 12947 11512 12992 11540
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 14568 11540 14596 11580
rect 18524 11580 19380 11608
rect 21744 11580 22232 11608
rect 22296 11580 24492 11608
rect 15470 11540 15476 11552
rect 14568 11512 15476 11540
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 16022 11540 16028 11552
rect 15983 11512 16028 11540
rect 16022 11500 16028 11512
rect 16080 11500 16086 11552
rect 16114 11500 16120 11552
rect 16172 11540 16178 11552
rect 18524 11540 18552 11580
rect 16172 11512 18552 11540
rect 16172 11500 16178 11512
rect 18690 11500 18696 11552
rect 18748 11540 18754 11552
rect 19337 11543 19395 11549
rect 19337 11540 19349 11543
rect 18748 11512 19349 11540
rect 18748 11500 18754 11512
rect 19337 11509 19349 11512
rect 19383 11540 19395 11543
rect 21744 11540 21772 11580
rect 21910 11540 21916 11552
rect 19383 11512 21772 11540
rect 21871 11512 21916 11540
rect 19383 11509 19395 11512
rect 19337 11503 19395 11509
rect 21910 11500 21916 11512
rect 21968 11500 21974 11552
rect 22204 11540 22232 11580
rect 24486 11568 24492 11580
rect 24544 11568 24550 11620
rect 27890 11568 27896 11620
rect 27948 11608 27954 11620
rect 31662 11608 31668 11620
rect 27948 11580 31668 11608
rect 27948 11568 27954 11580
rect 31662 11568 31668 11580
rect 31720 11568 31726 11620
rect 35434 11568 35440 11620
rect 35492 11568 35498 11620
rect 58158 11608 58164 11620
rect 58119 11580 58164 11608
rect 58158 11568 58164 11580
rect 58216 11568 58222 11620
rect 24118 11540 24124 11552
rect 22204 11512 24124 11540
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 31573 11543 31631 11549
rect 31573 11509 31585 11543
rect 31619 11540 31631 11543
rect 33042 11540 33048 11552
rect 31619 11512 33048 11540
rect 31619 11509 31631 11512
rect 31573 11503 31631 11509
rect 33042 11500 33048 11512
rect 33100 11500 33106 11552
rect 40770 11540 40776 11552
rect 40731 11512 40776 11540
rect 40770 11500 40776 11512
rect 40828 11500 40834 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 13446 11296 13452 11348
rect 13504 11336 13510 11348
rect 15933 11339 15991 11345
rect 15933 11336 15945 11339
rect 13504 11308 15945 11336
rect 13504 11296 13510 11308
rect 15933 11305 15945 11308
rect 15979 11305 15991 11339
rect 15933 11299 15991 11305
rect 18138 11296 18144 11348
rect 18196 11336 18202 11348
rect 18690 11336 18696 11348
rect 18196 11308 18696 11336
rect 18196 11296 18202 11308
rect 18690 11296 18696 11308
rect 18748 11296 18754 11348
rect 19058 11296 19064 11348
rect 19116 11336 19122 11348
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 19116 11308 19257 11336
rect 19116 11296 19122 11308
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 20162 11336 20168 11348
rect 20123 11308 20168 11336
rect 19245 11299 19303 11305
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 21634 11296 21640 11348
rect 21692 11336 21698 11348
rect 25038 11336 25044 11348
rect 21692 11308 25044 11336
rect 21692 11296 21698 11308
rect 25038 11296 25044 11308
rect 25096 11296 25102 11348
rect 25590 11296 25596 11348
rect 25648 11336 25654 11348
rect 25869 11339 25927 11345
rect 25869 11336 25881 11339
rect 25648 11308 25881 11336
rect 25648 11296 25654 11308
rect 25869 11305 25881 11308
rect 25915 11305 25927 11339
rect 25869 11299 25927 11305
rect 30282 11296 30288 11348
rect 30340 11336 30346 11348
rect 32493 11339 32551 11345
rect 32493 11336 32505 11339
rect 30340 11308 32505 11336
rect 30340 11296 30346 11308
rect 32493 11305 32505 11308
rect 32539 11336 32551 11339
rect 33410 11336 33416 11348
rect 32539 11308 33416 11336
rect 32539 11305 32551 11308
rect 32493 11299 32551 11305
rect 33410 11296 33416 11308
rect 33468 11296 33474 11348
rect 36998 11296 37004 11348
rect 37056 11336 37062 11348
rect 38102 11336 38108 11348
rect 37056 11308 38108 11336
rect 37056 11296 37062 11308
rect 38102 11296 38108 11308
rect 38160 11296 38166 11348
rect 38654 11336 38660 11348
rect 38615 11308 38660 11336
rect 38654 11296 38660 11308
rect 38712 11296 38718 11348
rect 15470 11268 15476 11280
rect 15431 11240 15476 11268
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 21177 11271 21235 11277
rect 21177 11237 21189 11271
rect 21223 11268 21235 11271
rect 21358 11268 21364 11280
rect 21223 11240 21364 11268
rect 21223 11237 21235 11240
rect 21177 11231 21235 11237
rect 21358 11228 21364 11240
rect 21416 11228 21422 11280
rect 29086 11228 29092 11280
rect 29144 11268 29150 11280
rect 29362 11268 29368 11280
rect 29144 11240 29368 11268
rect 29144 11228 29150 11240
rect 29362 11228 29368 11240
rect 29420 11228 29426 11280
rect 39022 11268 39028 11280
rect 35728 11240 39028 11268
rect 5626 11160 5632 11212
rect 5684 11200 5690 11212
rect 6457 11203 6515 11209
rect 6457 11200 6469 11203
rect 5684 11172 6469 11200
rect 5684 11160 5690 11172
rect 6457 11169 6469 11172
rect 6503 11200 6515 11203
rect 6546 11200 6552 11212
rect 6503 11172 6552 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 6546 11160 6552 11172
rect 6604 11160 6610 11212
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 14093 11203 14151 11209
rect 14093 11200 14105 11203
rect 12584 11172 14105 11200
rect 12584 11160 12590 11172
rect 14093 11169 14105 11172
rect 14139 11169 14151 11203
rect 14093 11163 14151 11169
rect 6178 11132 6184 11144
rect 6139 11104 6184 11132
rect 6178 11092 6184 11104
rect 6236 11092 6242 11144
rect 9766 11092 9772 11144
rect 9824 11132 9830 11144
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 9824 11104 10333 11132
rect 9824 11092 9830 11104
rect 10321 11101 10333 11104
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 14349 11135 14407 11141
rect 14349 11132 14361 11135
rect 13044 11104 14361 11132
rect 13044 11092 13050 11104
rect 14349 11101 14361 11104
rect 14395 11101 14407 11135
rect 15488 11132 15516 11228
rect 21634 11200 21640 11212
rect 21595 11172 21640 11200
rect 21634 11160 21640 11172
rect 21692 11160 21698 11212
rect 23842 11200 23848 11212
rect 23803 11172 23848 11200
rect 23842 11160 23848 11172
rect 23900 11160 23906 11212
rect 24118 11160 24124 11212
rect 24176 11200 24182 11212
rect 31018 11200 31024 11212
rect 24176 11172 31024 11200
rect 24176 11160 24182 11172
rect 16117 11135 16175 11141
rect 16117 11132 16129 11135
rect 15488 11104 16129 11132
rect 14349 11095 14407 11101
rect 16117 11101 16129 11104
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11132 16359 11135
rect 16666 11132 16672 11144
rect 16347 11104 16672 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 16666 11092 16672 11104
rect 16724 11092 16730 11144
rect 20349 11135 20407 11141
rect 20349 11101 20361 11135
rect 20395 11132 20407 11135
rect 21082 11132 21088 11144
rect 20395 11104 21088 11132
rect 20395 11101 20407 11104
rect 20349 11095 20407 11101
rect 21082 11092 21088 11104
rect 21140 11092 21146 11144
rect 21910 11141 21916 11144
rect 21904 11132 21916 11141
rect 21871 11104 21916 11132
rect 21904 11095 21916 11104
rect 21910 11092 21916 11095
rect 21968 11092 21974 11144
rect 23014 11092 23020 11144
rect 23072 11132 23078 11144
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 23072 11104 23673 11132
rect 23072 11092 23078 11104
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 24578 11092 24584 11144
rect 24636 11132 24642 11144
rect 24765 11135 24823 11141
rect 24765 11132 24777 11135
rect 24636 11104 24777 11132
rect 24636 11092 24642 11104
rect 24765 11101 24777 11104
rect 24811 11101 24823 11135
rect 24946 11132 24952 11144
rect 24907 11104 24952 11132
rect 24765 11095 24823 11101
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 25148 11141 25176 11172
rect 31018 11160 31024 11172
rect 31076 11160 31082 11212
rect 25041 11135 25099 11141
rect 25041 11101 25053 11135
rect 25087 11101 25099 11135
rect 25041 11095 25099 11101
rect 25133 11135 25191 11141
rect 25133 11101 25145 11135
rect 25179 11101 25191 11135
rect 26050 11132 26056 11144
rect 26011 11104 26056 11132
rect 25133 11095 25191 11101
rect 10134 11064 10140 11076
rect 10095 11036 10140 11064
rect 10134 11024 10140 11036
rect 10192 11024 10198 11076
rect 11330 11024 11336 11076
rect 11388 11064 11394 11076
rect 12710 11064 12716 11076
rect 11388 11036 12716 11064
rect 11388 11024 11394 11036
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 14918 11064 14924 11076
rect 14240 11036 14924 11064
rect 14240 11024 14246 11036
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 20990 11064 20996 11076
rect 20951 11036 20996 11064
rect 20990 11024 20996 11036
rect 21048 11024 21054 11076
rect 24854 11024 24860 11076
rect 24912 11064 24918 11076
rect 25056 11064 25084 11095
rect 26050 11092 26056 11104
rect 26108 11092 26114 11144
rect 26142 11092 26148 11144
rect 26200 11132 26206 11144
rect 28353 11135 28411 11141
rect 28353 11132 28365 11135
rect 26200 11104 28365 11132
rect 26200 11092 26206 11104
rect 28353 11101 28365 11104
rect 28399 11101 28411 11135
rect 28353 11095 28411 11101
rect 28442 11092 28448 11144
rect 28500 11132 28506 11144
rect 29086 11132 29092 11144
rect 28500 11104 29092 11132
rect 28500 11092 28506 11104
rect 29086 11092 29092 11104
rect 29144 11092 29150 11144
rect 30926 11092 30932 11144
rect 30984 11132 30990 11144
rect 31113 11135 31171 11141
rect 31113 11132 31125 11135
rect 30984 11104 31125 11132
rect 30984 11092 30990 11104
rect 31113 11101 31125 11104
rect 31159 11101 31171 11135
rect 35618 11132 35624 11144
rect 35579 11104 35624 11132
rect 31113 11095 31171 11101
rect 35618 11092 35624 11104
rect 35676 11092 35682 11144
rect 35728 11141 35756 11240
rect 39022 11228 39028 11240
rect 39080 11228 39086 11280
rect 36449 11203 36507 11209
rect 36449 11200 36461 11203
rect 35820 11172 36461 11200
rect 35820 11141 35848 11172
rect 36449 11169 36461 11172
rect 36495 11169 36507 11203
rect 36449 11163 36507 11169
rect 35713 11135 35771 11141
rect 35713 11101 35725 11135
rect 35759 11101 35771 11135
rect 35713 11095 35771 11101
rect 35805 11135 35863 11141
rect 35805 11101 35817 11135
rect 35851 11101 35863 11135
rect 35805 11095 35863 11101
rect 35989 11135 36047 11141
rect 35989 11101 36001 11135
rect 36035 11101 36047 11135
rect 36630 11132 36636 11144
rect 36591 11104 36636 11132
rect 35989 11095 36047 11101
rect 26234 11064 26240 11076
rect 24912 11036 25084 11064
rect 26195 11036 26240 11064
rect 24912 11024 24918 11036
rect 26234 11024 26240 11036
rect 26292 11024 26298 11076
rect 28537 11067 28595 11073
rect 28537 11033 28549 11067
rect 28583 11064 28595 11067
rect 28626 11064 28632 11076
rect 28583 11036 28632 11064
rect 28583 11033 28595 11036
rect 28537 11027 28595 11033
rect 28626 11024 28632 11036
rect 28684 11024 28690 11076
rect 31386 11073 31392 11076
rect 31380 11027 31392 11073
rect 31444 11064 31450 11076
rect 34885 11067 34943 11073
rect 34885 11064 34897 11067
rect 31444 11036 31480 11064
rect 32048 11036 34897 11064
rect 31386 11024 31392 11027
rect 31444 11024 31450 11036
rect 9401 10999 9459 11005
rect 9401 10965 9413 10999
rect 9447 10996 9459 10999
rect 9674 10996 9680 11008
rect 9447 10968 9680 10996
rect 9447 10965 9459 10968
rect 9401 10959 9459 10965
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 15010 10996 15016 11008
rect 11940 10968 15016 10996
rect 11940 10956 11946 10968
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 15654 10956 15660 11008
rect 15712 10996 15718 11008
rect 16482 10996 16488 11008
rect 15712 10968 16488 10996
rect 15712 10956 15718 10968
rect 16482 10956 16488 10968
rect 16540 10996 16546 11008
rect 19426 10996 19432 11008
rect 16540 10968 19432 10996
rect 16540 10956 16546 10968
rect 19426 10956 19432 10968
rect 19484 10956 19490 11008
rect 22462 10956 22468 11008
rect 22520 10996 22526 11008
rect 23017 10999 23075 11005
rect 23017 10996 23029 10999
rect 22520 10968 23029 10996
rect 22520 10956 22526 10968
rect 23017 10965 23029 10968
rect 23063 10965 23075 10999
rect 23474 10996 23480 11008
rect 23387 10968 23480 10996
rect 23017 10959 23075 10965
rect 23474 10956 23480 10968
rect 23532 10996 23538 11008
rect 24670 10996 24676 11008
rect 23532 10968 24676 10996
rect 23532 10956 23538 10968
rect 24670 10956 24676 10968
rect 24728 10956 24734 11008
rect 25406 10996 25412 11008
rect 25367 10968 25412 10996
rect 25406 10956 25412 10968
rect 25464 10956 25470 11008
rect 30653 10999 30711 11005
rect 30653 10965 30665 10999
rect 30699 10996 30711 10999
rect 31478 10996 31484 11008
rect 30699 10968 31484 10996
rect 30699 10965 30711 10968
rect 30653 10959 30711 10965
rect 31478 10956 31484 10968
rect 31536 10956 31542 11008
rect 31662 10956 31668 11008
rect 31720 10996 31726 11008
rect 32048 10996 32076 11036
rect 34885 11033 34897 11036
rect 34931 11064 34943 11067
rect 36004 11064 36032 11095
rect 36630 11092 36636 11104
rect 36688 11092 36694 11144
rect 37645 11135 37703 11141
rect 37645 11101 37657 11135
rect 37691 11132 37703 11135
rect 38470 11132 38476 11144
rect 37691 11104 38476 11132
rect 37691 11101 37703 11104
rect 37645 11095 37703 11101
rect 38470 11092 38476 11104
rect 38528 11132 38534 11144
rect 39040 11141 39068 11228
rect 40770 11200 40776 11212
rect 39132 11172 40776 11200
rect 39132 11141 39160 11172
rect 40770 11160 40776 11172
rect 40828 11160 40834 11212
rect 38933 11135 38991 11141
rect 38933 11132 38945 11135
rect 38528 11104 38945 11132
rect 38528 11092 38534 11104
rect 38933 11101 38945 11104
rect 38979 11101 38991 11135
rect 38933 11095 38991 11101
rect 39025 11135 39083 11141
rect 39025 11101 39037 11135
rect 39071 11101 39083 11135
rect 39025 11095 39083 11101
rect 39117 11135 39175 11141
rect 39117 11101 39129 11135
rect 39163 11101 39175 11135
rect 39117 11095 39175 11101
rect 39301 11135 39359 11141
rect 39301 11101 39313 11135
rect 39347 11101 39359 11135
rect 39301 11095 39359 11101
rect 34931 11036 36032 11064
rect 36817 11067 36875 11073
rect 34931 11033 34943 11036
rect 34885 11027 34943 11033
rect 36817 11033 36829 11067
rect 36863 11064 36875 11067
rect 37550 11064 37556 11076
rect 36863 11036 37556 11064
rect 36863 11033 36875 11036
rect 36817 11027 36875 11033
rect 37550 11024 37556 11036
rect 37608 11064 37614 11076
rect 38286 11064 38292 11076
rect 37608 11036 38292 11064
rect 37608 11024 37614 11036
rect 38286 11024 38292 11036
rect 38344 11024 38350 11076
rect 39316 11064 39344 11095
rect 38672 11036 39344 11064
rect 35342 10996 35348 11008
rect 31720 10968 32076 10996
rect 35303 10968 35348 10996
rect 31720 10956 31726 10968
rect 35342 10956 35348 10968
rect 35400 10956 35406 11008
rect 38102 10956 38108 11008
rect 38160 10996 38166 11008
rect 38672 10996 38700 11036
rect 38160 10968 38700 10996
rect 38160 10956 38166 10968
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 6270 10752 6276 10804
rect 6328 10792 6334 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 6328 10764 6377 10792
rect 6328 10752 6334 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 8849 10795 8907 10801
rect 8849 10761 8861 10795
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 8864 10724 8892 10755
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 12032 10764 12173 10792
rect 12032 10752 12038 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 12161 10755 12219 10761
rect 15010 10752 15016 10804
rect 15068 10792 15074 10804
rect 17586 10792 17592 10804
rect 15068 10764 17592 10792
rect 15068 10752 15074 10764
rect 17586 10752 17592 10764
rect 17644 10752 17650 10804
rect 22189 10795 22247 10801
rect 22189 10761 22201 10795
rect 22235 10792 22247 10795
rect 22370 10792 22376 10804
rect 22235 10764 22376 10792
rect 22235 10761 22247 10764
rect 22189 10755 22247 10761
rect 22370 10752 22376 10764
rect 22428 10752 22434 10804
rect 23658 10752 23664 10804
rect 23716 10792 23722 10804
rect 27433 10795 27491 10801
rect 27433 10792 27445 10795
rect 23716 10764 27445 10792
rect 23716 10752 23722 10764
rect 27433 10761 27445 10764
rect 27479 10792 27491 10795
rect 27479 10764 28672 10792
rect 27479 10761 27491 10764
rect 27433 10755 27491 10761
rect 5460 10696 8892 10724
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 5460 10665 5488 10696
rect 9214 10684 9220 10736
rect 9272 10724 9278 10736
rect 9769 10727 9827 10733
rect 9769 10724 9781 10727
rect 9272 10696 9781 10724
rect 9272 10684 9278 10696
rect 9769 10693 9781 10696
rect 9815 10724 9827 10727
rect 12618 10724 12624 10736
rect 9815 10696 12624 10724
rect 9815 10693 9827 10696
rect 9769 10687 9827 10693
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 17310 10724 17316 10736
rect 17271 10696 17316 10724
rect 17310 10684 17316 10696
rect 17368 10684 17374 10736
rect 22557 10727 22615 10733
rect 22557 10693 22569 10727
rect 22603 10724 22615 10727
rect 23474 10724 23480 10736
rect 22603 10696 23480 10724
rect 22603 10693 22615 10696
rect 22557 10687 22615 10693
rect 23474 10684 23480 10696
rect 23532 10684 23538 10736
rect 24762 10724 24768 10736
rect 23584 10696 24768 10724
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 4672 10628 5457 10656
rect 4672 10616 4678 10628
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 6546 10656 6552 10668
rect 6507 10628 6552 10656
rect 5445 10619 5503 10625
rect 6546 10616 6552 10628
rect 6604 10616 6610 10668
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10656 7067 10659
rect 7282 10656 7288 10668
rect 7055 10628 7288 10656
rect 7055 10625 7067 10628
rect 7009 10619 7067 10625
rect 7282 10616 7288 10628
rect 7340 10656 7346 10668
rect 9950 10656 9956 10668
rect 7340 10628 9956 10656
rect 7340 10616 7346 10628
rect 9950 10616 9956 10628
rect 10008 10656 10014 10668
rect 10134 10656 10140 10668
rect 10008 10628 10140 10656
rect 10008 10616 10014 10628
rect 10134 10616 10140 10628
rect 10192 10616 10198 10668
rect 10410 10616 10416 10668
rect 10468 10656 10474 10668
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 10468 10628 11897 10656
rect 10468 10616 10474 10628
rect 11885 10625 11897 10628
rect 11931 10625 11943 10659
rect 17126 10656 17132 10668
rect 17087 10628 17132 10656
rect 11885 10619 11943 10625
rect 17126 10616 17132 10628
rect 17184 10616 17190 10668
rect 22373 10659 22431 10665
rect 22373 10625 22385 10659
rect 22419 10656 22431 10659
rect 22462 10656 22468 10668
rect 22419 10628 22468 10656
rect 22419 10625 22431 10628
rect 22373 10619 22431 10625
rect 22462 10616 22468 10628
rect 22520 10616 22526 10668
rect 23014 10656 23020 10668
rect 22975 10628 23020 10656
rect 23014 10616 23020 10628
rect 23072 10616 23078 10668
rect 23201 10659 23259 10665
rect 23201 10625 23213 10659
rect 23247 10625 23259 10659
rect 23201 10619 23259 10625
rect 4890 10548 4896 10600
rect 4948 10588 4954 10600
rect 6641 10591 6699 10597
rect 6641 10588 6653 10591
rect 4948 10560 6653 10588
rect 4948 10548 4954 10560
rect 6641 10557 6653 10560
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10557 8723 10591
rect 8665 10551 8723 10557
rect 9033 10591 9091 10597
rect 9033 10557 9045 10591
rect 9079 10588 9091 10591
rect 9674 10588 9680 10600
rect 9079 10560 9680 10588
rect 9079 10557 9091 10560
rect 9033 10551 9091 10557
rect 5626 10520 5632 10532
rect 5587 10492 5632 10520
rect 5626 10480 5632 10492
rect 5684 10520 5690 10532
rect 5994 10520 6000 10532
rect 5684 10492 6000 10520
rect 5684 10480 5690 10492
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 8680 10520 8708 10551
rect 9674 10548 9680 10560
rect 9732 10588 9738 10600
rect 10870 10588 10876 10600
rect 9732 10560 10876 10588
rect 9732 10548 9738 10560
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 11514 10588 11520 10600
rect 11475 10560 11520 10588
rect 11514 10548 11520 10560
rect 11572 10548 11578 10600
rect 11974 10588 11980 10600
rect 11935 10560 11980 10588
rect 11974 10548 11980 10560
rect 12032 10548 12038 10600
rect 21358 10548 21364 10600
rect 21416 10588 21422 10600
rect 22830 10588 22836 10600
rect 21416 10560 22836 10588
rect 21416 10548 21422 10560
rect 22830 10548 22836 10560
rect 22888 10588 22894 10600
rect 23216 10588 23244 10619
rect 23290 10616 23296 10668
rect 23348 10656 23354 10668
rect 23584 10656 23612 10696
rect 24762 10684 24768 10696
rect 24820 10684 24826 10736
rect 25308 10727 25366 10733
rect 25308 10693 25320 10727
rect 25354 10724 25366 10727
rect 25406 10724 25412 10736
rect 25354 10696 25412 10724
rect 25354 10693 25366 10696
rect 25308 10687 25366 10693
rect 25406 10684 25412 10696
rect 25464 10684 25470 10736
rect 28644 10733 28672 10764
rect 31110 10752 31116 10804
rect 31168 10792 31174 10804
rect 31573 10795 31631 10801
rect 31573 10792 31585 10795
rect 31168 10764 31585 10792
rect 31168 10752 31174 10764
rect 31573 10761 31585 10764
rect 31619 10761 31631 10795
rect 36630 10792 36636 10804
rect 36591 10764 36636 10792
rect 31573 10755 31631 10761
rect 36630 10752 36636 10764
rect 36688 10752 36694 10804
rect 38102 10752 38108 10804
rect 38160 10792 38166 10804
rect 38381 10795 38439 10801
rect 38381 10792 38393 10795
rect 38160 10764 38393 10792
rect 38160 10752 38166 10764
rect 38381 10761 38393 10764
rect 38427 10792 38439 10795
rect 38427 10764 39344 10792
rect 38427 10761 38439 10764
rect 38381 10755 38439 10761
rect 28629 10727 28687 10733
rect 28629 10693 28641 10727
rect 28675 10693 28687 10727
rect 28629 10687 28687 10693
rect 33042 10684 33048 10736
rect 33100 10724 33106 10736
rect 33238 10727 33296 10733
rect 33238 10724 33250 10727
rect 33100 10696 33250 10724
rect 33100 10684 33106 10696
rect 33238 10693 33250 10696
rect 33284 10693 33296 10727
rect 38562 10724 38568 10736
rect 33238 10687 33296 10693
rect 35268 10696 38568 10724
rect 23348 10628 23612 10656
rect 23348 10616 23354 10628
rect 24210 10616 24216 10668
rect 24268 10656 24274 10668
rect 24305 10659 24363 10665
rect 24305 10656 24317 10659
rect 24268 10628 24317 10656
rect 24268 10616 24274 10628
rect 24305 10625 24317 10628
rect 24351 10656 24363 10659
rect 24854 10656 24860 10668
rect 24351 10628 24860 10656
rect 24351 10625 24363 10628
rect 24305 10619 24363 10625
rect 24854 10616 24860 10628
rect 24912 10616 24918 10668
rect 25038 10656 25044 10668
rect 24999 10628 25044 10656
rect 25038 10616 25044 10628
rect 25096 10616 25102 10668
rect 26234 10656 26240 10668
rect 25148 10628 26240 10656
rect 22888 10560 23244 10588
rect 22888 10548 22894 10560
rect 24486 10548 24492 10600
rect 24544 10588 24550 10600
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 24544 10560 24593 10588
rect 24544 10548 24550 10560
rect 24581 10557 24593 10560
rect 24627 10557 24639 10591
rect 24581 10551 24639 10557
rect 24670 10548 24676 10600
rect 24728 10588 24734 10600
rect 25148 10588 25176 10628
rect 26234 10616 26240 10628
rect 26292 10656 26298 10668
rect 27985 10659 28043 10665
rect 27985 10656 27997 10659
rect 26292 10628 27997 10656
rect 26292 10616 26298 10628
rect 27985 10625 27997 10628
rect 28031 10625 28043 10659
rect 27985 10619 28043 10625
rect 30282 10616 30288 10668
rect 30340 10656 30346 10668
rect 31205 10659 31263 10665
rect 31205 10656 31217 10659
rect 30340 10628 31217 10656
rect 30340 10616 30346 10628
rect 31205 10625 31217 10628
rect 31251 10625 31263 10659
rect 31205 10619 31263 10625
rect 31389 10659 31447 10665
rect 31389 10625 31401 10659
rect 31435 10656 31447 10659
rect 31938 10656 31944 10668
rect 31435 10628 31944 10656
rect 31435 10625 31447 10628
rect 31389 10619 31447 10625
rect 31938 10616 31944 10628
rect 31996 10616 32002 10668
rect 24728 10560 25176 10588
rect 33505 10591 33563 10597
rect 24728 10548 24734 10560
rect 33505 10557 33517 10591
rect 33551 10588 33563 10591
rect 34698 10588 34704 10600
rect 33551 10560 34704 10588
rect 33551 10557 33563 10560
rect 33505 10551 33563 10557
rect 34698 10548 34704 10560
rect 34756 10588 34762 10600
rect 35268 10597 35296 10696
rect 38562 10684 38568 10696
rect 38620 10684 38626 10736
rect 39316 10724 39344 10764
rect 39316 10696 39620 10724
rect 35342 10616 35348 10668
rect 35400 10656 35406 10668
rect 35509 10659 35567 10665
rect 35509 10656 35521 10659
rect 35400 10628 35521 10656
rect 35400 10616 35406 10628
rect 35509 10625 35521 10628
rect 35555 10625 35567 10659
rect 35509 10619 35567 10625
rect 37734 10616 37740 10668
rect 37792 10656 37798 10668
rect 37921 10659 37979 10665
rect 37921 10656 37933 10659
rect 37792 10628 37933 10656
rect 37792 10616 37798 10628
rect 37921 10625 37933 10628
rect 37967 10656 37979 10659
rect 39209 10659 39267 10665
rect 39209 10656 39221 10659
rect 37967 10628 39221 10656
rect 37967 10625 37979 10628
rect 37921 10619 37979 10625
rect 39209 10625 39221 10628
rect 39255 10625 39267 10659
rect 39209 10619 39267 10625
rect 39301 10659 39359 10665
rect 39301 10625 39313 10659
rect 39347 10625 39359 10659
rect 39301 10619 39359 10625
rect 35253 10591 35311 10597
rect 35253 10588 35265 10591
rect 34756 10560 35265 10588
rect 34756 10548 34762 10560
rect 35253 10557 35265 10560
rect 35299 10557 35311 10591
rect 35253 10551 35311 10557
rect 39022 10548 39028 10600
rect 39080 10588 39086 10600
rect 39316 10588 39344 10619
rect 39390 10616 39396 10668
rect 39448 10656 39454 10668
rect 39592 10665 39620 10696
rect 39577 10659 39635 10665
rect 39448 10628 39493 10656
rect 39448 10616 39454 10628
rect 39577 10625 39589 10659
rect 39623 10625 39635 10659
rect 39577 10619 39635 10625
rect 39080 10560 39344 10588
rect 39080 10548 39086 10560
rect 14090 10520 14096 10532
rect 8680 10492 14096 10520
rect 14090 10480 14096 10492
rect 14148 10480 14154 10532
rect 23109 10523 23167 10529
rect 23109 10489 23121 10523
rect 23155 10520 23167 10523
rect 24504 10520 24532 10548
rect 23155 10492 24532 10520
rect 23155 10489 23167 10492
rect 23109 10483 23167 10489
rect 27062 10480 27068 10532
rect 27120 10520 27126 10532
rect 27120 10492 29960 10520
rect 27120 10480 27126 10492
rect 29932 10464 29960 10492
rect 30374 10480 30380 10532
rect 30432 10520 30438 10532
rect 30432 10492 32628 10520
rect 30432 10480 30438 10492
rect 9214 10452 9220 10464
rect 9175 10424 9220 10452
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 18138 10412 18144 10464
rect 18196 10452 18202 10464
rect 18969 10455 19027 10461
rect 18969 10452 18981 10455
rect 18196 10424 18981 10452
rect 18196 10412 18202 10424
rect 18969 10421 18981 10424
rect 19015 10452 19027 10455
rect 19242 10452 19248 10464
rect 19015 10424 19248 10452
rect 19015 10421 19027 10424
rect 18969 10415 19027 10421
rect 19242 10412 19248 10424
rect 19300 10412 19306 10464
rect 20809 10455 20867 10461
rect 20809 10421 20821 10455
rect 20855 10452 20867 10455
rect 20990 10452 20996 10464
rect 20855 10424 20996 10452
rect 20855 10421 20867 10424
rect 20809 10415 20867 10421
rect 20990 10412 20996 10424
rect 21048 10452 21054 10464
rect 21634 10452 21640 10464
rect 21048 10424 21640 10452
rect 21048 10412 21054 10424
rect 21634 10412 21640 10424
rect 21692 10412 21698 10464
rect 25406 10412 25412 10464
rect 25464 10452 25470 10464
rect 26421 10455 26479 10461
rect 26421 10452 26433 10455
rect 25464 10424 26433 10452
rect 25464 10412 25470 10424
rect 26421 10421 26433 10424
rect 26467 10452 26479 10455
rect 27982 10452 27988 10464
rect 26467 10424 27988 10452
rect 26467 10421 26479 10424
rect 26421 10415 26479 10421
rect 27982 10412 27988 10424
rect 28040 10412 28046 10464
rect 28169 10455 28227 10461
rect 28169 10421 28181 10455
rect 28215 10452 28227 10455
rect 29546 10452 29552 10464
rect 28215 10424 29552 10452
rect 28215 10421 28227 10424
rect 28169 10415 28227 10421
rect 29546 10412 29552 10424
rect 29604 10412 29610 10464
rect 29914 10452 29920 10464
rect 29875 10424 29920 10452
rect 29914 10412 29920 10424
rect 29972 10412 29978 10464
rect 31938 10412 31944 10464
rect 31996 10452 32002 10464
rect 32125 10455 32183 10461
rect 32125 10452 32137 10455
rect 31996 10424 32137 10452
rect 31996 10412 32002 10424
rect 32125 10421 32137 10424
rect 32171 10452 32183 10455
rect 32398 10452 32404 10464
rect 32171 10424 32404 10452
rect 32171 10421 32183 10424
rect 32125 10415 32183 10421
rect 32398 10412 32404 10424
rect 32456 10412 32462 10464
rect 32600 10452 32628 10492
rect 34514 10452 34520 10464
rect 32600 10424 34520 10452
rect 34514 10412 34520 10424
rect 34572 10412 34578 10464
rect 34793 10455 34851 10461
rect 34793 10421 34805 10455
rect 34839 10452 34851 10455
rect 35618 10452 35624 10464
rect 34839 10424 35624 10452
rect 34839 10421 34851 10424
rect 34793 10415 34851 10421
rect 35618 10412 35624 10424
rect 35676 10412 35682 10464
rect 38930 10452 38936 10464
rect 38891 10424 38936 10452
rect 38930 10412 38936 10424
rect 38988 10412 38994 10464
rect 58158 10452 58164 10464
rect 58119 10424 58164 10452
rect 58158 10412 58164 10424
rect 58216 10412 58222 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 16482 10248 16488 10260
rect 16443 10220 16488 10248
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 22830 10248 22836 10260
rect 22791 10220 22836 10248
rect 22830 10208 22836 10220
rect 22888 10208 22894 10260
rect 24946 10208 24952 10260
rect 25004 10248 25010 10260
rect 25225 10251 25283 10257
rect 25225 10248 25237 10251
rect 25004 10220 25237 10248
rect 25004 10208 25010 10220
rect 25225 10217 25237 10220
rect 25271 10217 25283 10251
rect 25225 10211 25283 10217
rect 28261 10251 28319 10257
rect 28261 10217 28273 10251
rect 28307 10248 28319 10251
rect 28534 10248 28540 10260
rect 28307 10220 28540 10248
rect 28307 10217 28319 10220
rect 28261 10211 28319 10217
rect 28534 10208 28540 10220
rect 28592 10208 28598 10260
rect 28997 10251 29055 10257
rect 28997 10217 29009 10251
rect 29043 10248 29055 10251
rect 29270 10248 29276 10260
rect 29043 10220 29276 10248
rect 29043 10217 29055 10220
rect 28997 10211 29055 10217
rect 29270 10208 29276 10220
rect 29328 10208 29334 10260
rect 38562 10248 38568 10260
rect 38523 10220 38568 10248
rect 38562 10208 38568 10220
rect 38620 10208 38626 10260
rect 4985 10183 5043 10189
rect 4985 10180 4997 10183
rect 2746 10152 4997 10180
rect 2746 10112 2774 10152
rect 4985 10149 4997 10152
rect 5031 10149 5043 10183
rect 4985 10143 5043 10149
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 9953 10183 10011 10189
rect 9953 10180 9965 10183
rect 8260 10152 9965 10180
rect 8260 10140 8266 10152
rect 9953 10149 9965 10152
rect 9999 10149 10011 10183
rect 9953 10143 10011 10149
rect 24302 10140 24308 10192
rect 24360 10180 24366 10192
rect 30374 10180 30380 10192
rect 24360 10152 30380 10180
rect 24360 10140 24366 10152
rect 30374 10140 30380 10152
rect 30432 10140 30438 10192
rect 5626 10112 5632 10124
rect 2700 10084 2774 10112
rect 5539 10084 5632 10112
rect 2700 10053 2728 10084
rect 5626 10072 5632 10084
rect 5684 10112 5690 10124
rect 10410 10112 10416 10124
rect 5684 10084 9076 10112
rect 10371 10084 10416 10112
rect 5684 10072 5690 10084
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10013 2743 10047
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2685 10007 2743 10013
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 6178 10004 6184 10056
rect 6236 10044 6242 10056
rect 6273 10047 6331 10053
rect 6273 10044 6285 10047
rect 6236 10016 6285 10044
rect 6236 10004 6242 10016
rect 6273 10013 6285 10016
rect 6319 10013 6331 10047
rect 8938 10044 8944 10056
rect 8899 10016 8944 10044
rect 6273 10007 6331 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9048 10044 9076 10084
rect 10410 10072 10416 10084
rect 10468 10072 10474 10124
rect 10597 10115 10655 10121
rect 10597 10081 10609 10115
rect 10643 10112 10655 10115
rect 13538 10112 13544 10124
rect 10643 10084 13544 10112
rect 10643 10081 10655 10084
rect 10597 10075 10655 10081
rect 10612 10044 10640 10075
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 24486 10072 24492 10124
rect 24544 10112 24550 10124
rect 26602 10112 26608 10124
rect 24544 10084 26608 10112
rect 24544 10072 24550 10084
rect 26602 10072 26608 10084
rect 26660 10072 26666 10124
rect 28626 10072 28632 10124
rect 28684 10112 28690 10124
rect 31202 10112 31208 10124
rect 28684 10084 31208 10112
rect 28684 10072 28690 10084
rect 9048 10016 10640 10044
rect 24581 10047 24639 10053
rect 24581 10013 24593 10047
rect 24627 10044 24639 10047
rect 24670 10044 24676 10056
rect 24627 10016 24676 10044
rect 24627 10013 24639 10016
rect 24581 10007 24639 10013
rect 24670 10004 24676 10016
rect 24728 10004 24734 10056
rect 25406 10044 25412 10056
rect 25367 10016 25412 10044
rect 25406 10004 25412 10016
rect 25464 10004 25470 10056
rect 27706 10044 27712 10056
rect 27667 10016 27712 10044
rect 27706 10004 27712 10016
rect 27764 10004 27770 10056
rect 27982 10044 27988 10056
rect 27943 10016 27988 10044
rect 27982 10004 27988 10016
rect 28040 10004 28046 10056
rect 28077 10047 28135 10053
rect 28077 10013 28089 10047
rect 28123 10044 28135 10047
rect 28534 10044 28540 10056
rect 28123 10016 28540 10044
rect 28123 10013 28135 10016
rect 28077 10007 28135 10013
rect 28534 10004 28540 10016
rect 28592 10004 28598 10056
rect 29270 10004 29276 10056
rect 29328 10044 29334 10056
rect 29932 10053 29960 10084
rect 31202 10072 31208 10084
rect 31260 10072 31266 10124
rect 29825 10047 29883 10053
rect 29825 10044 29837 10047
rect 29328 10016 29837 10044
rect 29328 10004 29334 10016
rect 29825 10013 29837 10016
rect 29871 10013 29883 10047
rect 29825 10007 29883 10013
rect 29917 10047 29975 10053
rect 29917 10013 29929 10047
rect 29963 10013 29975 10047
rect 29917 10007 29975 10013
rect 30006 10004 30012 10056
rect 30064 10044 30070 10056
rect 30193 10047 30251 10053
rect 30064 10016 30109 10044
rect 30064 10004 30070 10016
rect 30193 10013 30205 10047
rect 30239 10044 30251 10047
rect 32122 10044 32128 10056
rect 30239 10016 32128 10044
rect 30239 10013 30251 10016
rect 30193 10007 30251 10013
rect 32122 10004 32128 10016
rect 32180 10004 32186 10056
rect 36633 10047 36691 10053
rect 36633 10013 36645 10047
rect 36679 10044 36691 10047
rect 37093 10047 37151 10053
rect 37093 10044 37105 10047
rect 36679 10016 37105 10044
rect 36679 10013 36691 10016
rect 36633 10007 36691 10013
rect 37093 10013 37105 10016
rect 37139 10044 37151 10047
rect 37182 10044 37188 10056
rect 37139 10016 37188 10044
rect 37139 10013 37151 10016
rect 37093 10007 37151 10013
rect 37182 10004 37188 10016
rect 37240 10004 37246 10056
rect 5353 9979 5411 9985
rect 5353 9945 5365 9979
rect 5399 9976 5411 9979
rect 6454 9976 6460 9988
rect 5399 9948 6316 9976
rect 6367 9948 6460 9976
rect 5399 9945 5411 9948
rect 5353 9939 5411 9945
rect 1670 9868 1676 9920
rect 1728 9908 1734 9920
rect 2501 9911 2559 9917
rect 2501 9908 2513 9911
rect 1728 9880 2513 9908
rect 1728 9868 1734 9880
rect 2501 9877 2513 9880
rect 2547 9877 2559 9911
rect 2501 9871 2559 9877
rect 5442 9868 5448 9920
rect 5500 9908 5506 9920
rect 6288 9908 6316 9948
rect 6454 9936 6460 9948
rect 6512 9976 6518 9988
rect 11974 9976 11980 9988
rect 6512 9948 11980 9976
rect 6512 9936 6518 9948
rect 11974 9936 11980 9948
rect 12032 9936 12038 9988
rect 14090 9936 14096 9988
rect 14148 9976 14154 9988
rect 16577 9979 16635 9985
rect 16577 9976 16589 9979
rect 14148 9948 16589 9976
rect 14148 9936 14154 9948
rect 16577 9945 16589 9948
rect 16623 9976 16635 9979
rect 17126 9976 17132 9988
rect 16623 9948 17132 9976
rect 16623 9945 16635 9948
rect 16577 9939 16635 9945
rect 17126 9936 17132 9948
rect 17184 9936 17190 9988
rect 25593 9979 25651 9985
rect 25593 9945 25605 9979
rect 25639 9945 25651 9979
rect 25593 9939 25651 9945
rect 27893 9979 27951 9985
rect 27893 9945 27905 9979
rect 27939 9976 27951 9979
rect 28442 9976 28448 9988
rect 27939 9948 28448 9976
rect 27939 9945 27951 9948
rect 27893 9939 27951 9945
rect 6362 9908 6368 9920
rect 5500 9880 5545 9908
rect 6288 9880 6368 9908
rect 5500 9868 5506 9880
rect 6362 9868 6368 9880
rect 6420 9868 6426 9920
rect 6822 9868 6828 9920
rect 6880 9908 6886 9920
rect 8386 9908 8392 9920
rect 6880 9880 8392 9908
rect 6880 9868 6886 9880
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 9122 9908 9128 9920
rect 9083 9880 9128 9908
rect 9122 9868 9128 9880
rect 9180 9868 9186 9920
rect 10318 9908 10324 9920
rect 10279 9880 10324 9908
rect 10318 9868 10324 9880
rect 10376 9908 10382 9920
rect 11149 9911 11207 9917
rect 11149 9908 11161 9911
rect 10376 9880 11161 9908
rect 10376 9868 10382 9880
rect 11149 9877 11161 9880
rect 11195 9877 11207 9911
rect 11149 9871 11207 9877
rect 24670 9868 24676 9920
rect 24728 9908 24734 9920
rect 24765 9911 24823 9917
rect 24765 9908 24777 9911
rect 24728 9880 24777 9908
rect 24728 9868 24734 9880
rect 24765 9877 24777 9880
rect 24811 9908 24823 9911
rect 25608 9908 25636 9939
rect 28442 9936 28448 9948
rect 28500 9936 28506 9988
rect 24811 9880 25636 9908
rect 29549 9911 29607 9917
rect 24811 9877 24823 9880
rect 24765 9871 24823 9877
rect 29549 9877 29561 9911
rect 29595 9908 29607 9911
rect 30650 9908 30656 9920
rect 29595 9880 30656 9908
rect 29595 9877 29607 9880
rect 29549 9871 29607 9877
rect 30650 9868 30656 9880
rect 30708 9868 30714 9920
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 1857 9707 1915 9713
rect 1857 9673 1869 9707
rect 1903 9673 1915 9707
rect 1857 9667 1915 9673
rect 8389 9707 8447 9713
rect 8389 9673 8401 9707
rect 8435 9704 8447 9707
rect 8938 9704 8944 9716
rect 8435 9676 8944 9704
rect 8435 9673 8447 9676
rect 8389 9667 8447 9673
rect 1872 9636 1900 9667
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 10229 9707 10287 9713
rect 10229 9673 10241 9707
rect 10275 9704 10287 9707
rect 10410 9704 10416 9716
rect 10275 9676 10416 9704
rect 10275 9673 10287 9676
rect 10229 9667 10287 9673
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 19978 9664 19984 9716
rect 20036 9704 20042 9716
rect 21358 9704 21364 9716
rect 20036 9676 21364 9704
rect 20036 9664 20042 9676
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 22462 9664 22468 9716
rect 22520 9664 22526 9716
rect 29917 9707 29975 9713
rect 25608 9676 26188 9704
rect 2562 9639 2620 9645
rect 2562 9636 2574 9639
rect 1872 9608 2574 9636
rect 2562 9605 2574 9608
rect 2608 9605 2620 9639
rect 2562 9599 2620 9605
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 5534 9636 5540 9648
rect 4571 9608 5540 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 7282 9636 7288 9648
rect 7243 9608 7288 9636
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 9122 9645 9128 9648
rect 9116 9636 9128 9645
rect 9083 9608 9128 9636
rect 9116 9599 9128 9608
rect 9122 9596 9128 9599
rect 9180 9596 9186 9648
rect 9582 9596 9588 9648
rect 9640 9636 9646 9648
rect 16758 9636 16764 9648
rect 9640 9608 16764 9636
rect 9640 9596 9646 9608
rect 16758 9596 16764 9608
rect 16816 9596 16822 9648
rect 20714 9636 20720 9648
rect 20675 9608 20720 9636
rect 20714 9596 20720 9608
rect 20772 9596 20778 9648
rect 22480 9636 22508 9664
rect 25608 9645 25636 9676
rect 22741 9639 22799 9645
rect 22741 9636 22753 9639
rect 22480 9608 22753 9636
rect 22741 9605 22753 9608
rect 22787 9605 22799 9639
rect 25593 9639 25651 9645
rect 25593 9636 25605 9639
rect 22741 9599 22799 9605
rect 22940 9608 25605 9636
rect 22940 9580 22968 9608
rect 25593 9605 25605 9608
rect 25639 9605 25651 9639
rect 25593 9599 25651 9605
rect 25685 9639 25743 9645
rect 25685 9605 25697 9639
rect 25731 9636 25743 9639
rect 26050 9636 26056 9648
rect 25731 9608 26056 9636
rect 25731 9605 25743 9608
rect 25685 9599 25743 9605
rect 26050 9596 26056 9608
rect 26108 9596 26114 9648
rect 26160 9636 26188 9676
rect 29917 9673 29929 9707
rect 29963 9704 29975 9707
rect 30006 9704 30012 9716
rect 29963 9676 30012 9704
rect 29963 9673 29975 9676
rect 29917 9667 29975 9673
rect 30006 9664 30012 9676
rect 30064 9664 30070 9716
rect 39390 9704 39396 9716
rect 38580 9676 39396 9704
rect 28166 9636 28172 9648
rect 26160 9608 28172 9636
rect 28166 9596 28172 9608
rect 28224 9596 28230 9648
rect 29546 9636 29552 9648
rect 29459 9608 29552 9636
rect 29546 9596 29552 9608
rect 29604 9636 29610 9648
rect 30282 9636 30288 9648
rect 29604 9608 30288 9636
rect 29604 9596 29610 9608
rect 30282 9596 30288 9608
rect 30340 9596 30346 9648
rect 31573 9639 31631 9645
rect 31573 9605 31585 9639
rect 31619 9636 31631 9639
rect 35437 9639 35495 9645
rect 31619 9608 32536 9636
rect 31619 9605 31631 9608
rect 31573 9599 31631 9605
rect 32508 9580 32536 9608
rect 35437 9605 35449 9639
rect 35483 9636 35495 9639
rect 35802 9636 35808 9648
rect 35483 9608 35808 9636
rect 35483 9605 35495 9608
rect 35437 9599 35495 9605
rect 35802 9596 35808 9608
rect 35860 9596 35866 9648
rect 36354 9596 36360 9648
rect 36412 9636 36418 9648
rect 37550 9636 37556 9648
rect 36412 9608 37412 9636
rect 37511 9608 37556 9636
rect 36412 9596 36418 9608
rect 1670 9568 1676 9580
rect 1631 9540 1676 9568
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9568 4951 9571
rect 5442 9568 5448 9580
rect 4939 9540 5448 9568
rect 4939 9537 4951 9540
rect 4893 9531 4951 9537
rect 1854 9460 1860 9512
rect 1912 9500 1918 9512
rect 2317 9503 2375 9509
rect 2317 9500 2329 9503
rect 1912 9472 2329 9500
rect 1912 9460 1918 9472
rect 2317 9469 2329 9472
rect 2363 9469 2375 9503
rect 2317 9463 2375 9469
rect 3697 9435 3755 9441
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 4908 9432 4936 9531
rect 5442 9528 5448 9540
rect 5500 9528 5506 9580
rect 8202 9568 8208 9580
rect 8163 9540 8208 9568
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 13357 9571 13415 9577
rect 13357 9568 13369 9571
rect 12584 9540 13369 9568
rect 12584 9528 12590 9540
rect 13357 9537 13369 9540
rect 13403 9537 13415 9571
rect 14182 9568 14188 9580
rect 14143 9540 14188 9568
rect 13357 9531 13415 9537
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 14274 9528 14280 9580
rect 14332 9568 14338 9580
rect 14458 9568 14464 9580
rect 14332 9540 14464 9568
rect 14332 9528 14338 9540
rect 14458 9528 14464 9540
rect 14516 9528 14522 9580
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 18325 9571 18383 9577
rect 18325 9568 18337 9571
rect 17920 9540 18337 9568
rect 17920 9528 17926 9540
rect 18325 9537 18337 9540
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 18690 9528 18696 9580
rect 18748 9568 18754 9580
rect 22465 9571 22523 9577
rect 22465 9568 22477 9571
rect 18748 9540 22477 9568
rect 18748 9528 18754 9540
rect 22465 9537 22477 9540
rect 22511 9537 22523 9571
rect 22646 9568 22652 9580
rect 22607 9540 22652 9568
rect 22465 9531 22523 9537
rect 22646 9528 22652 9540
rect 22704 9528 22710 9580
rect 22833 9571 22891 9577
rect 22833 9537 22845 9571
rect 22879 9537 22891 9571
rect 22833 9531 22891 9537
rect 4985 9503 5043 9509
rect 4985 9469 4997 9503
rect 5031 9500 5043 9503
rect 5626 9500 5632 9512
rect 5031 9472 5632 9500
rect 5031 9469 5043 9472
rect 4985 9463 5043 9469
rect 5626 9460 5632 9472
rect 5684 9500 5690 9512
rect 6454 9500 6460 9512
rect 5684 9472 6460 9500
rect 5684 9460 5690 9472
rect 6454 9460 6460 9472
rect 6512 9460 6518 9512
rect 8021 9503 8079 9509
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8846 9500 8852 9512
rect 8067 9472 8248 9500
rect 8807 9472 8852 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8220 9432 8248 9472
rect 8846 9460 8852 9472
rect 8904 9460 8910 9512
rect 13449 9503 13507 9509
rect 13449 9469 13461 9503
rect 13495 9469 13507 9503
rect 13449 9463 13507 9469
rect 3743 9404 4936 9432
rect 5000 9404 8248 9432
rect 13464 9432 13492 9463
rect 13538 9460 13544 9512
rect 13596 9500 13602 9512
rect 13596 9472 13641 9500
rect 13596 9460 13602 9472
rect 22186 9460 22192 9512
rect 22244 9500 22250 9512
rect 22848 9500 22876 9531
rect 22922 9528 22928 9580
rect 22980 9528 22986 9580
rect 25406 9568 25412 9580
rect 25367 9540 25412 9568
rect 25406 9528 25412 9540
rect 25464 9528 25470 9580
rect 25777 9571 25835 9577
rect 25777 9537 25789 9571
rect 25823 9537 25835 9571
rect 29730 9568 29736 9580
rect 29691 9540 29736 9568
rect 25777 9531 25835 9537
rect 25792 9500 25820 9531
rect 29730 9528 29736 9540
rect 29788 9528 29794 9580
rect 32122 9568 32128 9580
rect 32083 9540 32128 9568
rect 32122 9528 32128 9540
rect 32180 9528 32186 9580
rect 32306 9568 32312 9580
rect 32267 9540 32312 9568
rect 32306 9528 32312 9540
rect 32364 9528 32370 9580
rect 32401 9571 32459 9577
rect 32401 9537 32413 9571
rect 32447 9537 32459 9571
rect 32401 9531 32459 9537
rect 28261 9503 28319 9509
rect 28261 9500 28273 9503
rect 22244 9472 28273 9500
rect 22244 9460 22250 9472
rect 28261 9469 28273 9472
rect 28307 9469 28319 9503
rect 28534 9500 28540 9512
rect 28495 9472 28540 9500
rect 28261 9463 28319 9469
rect 13906 9432 13912 9444
rect 13464 9404 13912 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 5000 9364 5028 9404
rect 4028 9336 5028 9364
rect 5169 9367 5227 9373
rect 4028 9324 4034 9336
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 6270 9364 6276 9376
rect 5215 9336 6276 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6362 9324 6368 9376
rect 6420 9364 6426 9376
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 6420 9336 6469 9364
rect 6420 9324 6426 9336
rect 6457 9333 6469 9336
rect 6503 9364 6515 9367
rect 6914 9364 6920 9376
rect 6503 9336 6920 9364
rect 6503 9333 6515 9336
rect 6457 9327 6515 9333
rect 6914 9324 6920 9336
rect 6972 9324 6978 9376
rect 7374 9364 7380 9376
rect 7335 9336 7380 9364
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 8220 9364 8248 9404
rect 13906 9392 13912 9404
rect 13964 9392 13970 9444
rect 23017 9435 23075 9441
rect 23017 9401 23029 9435
rect 23063 9432 23075 9435
rect 23382 9432 23388 9444
rect 23063 9404 23388 9432
rect 23063 9401 23075 9404
rect 23017 9395 23075 9401
rect 23382 9392 23388 9404
rect 23440 9392 23446 9444
rect 25961 9435 26019 9441
rect 25961 9401 25973 9435
rect 26007 9432 26019 9435
rect 26694 9432 26700 9444
rect 26007 9404 26700 9432
rect 26007 9401 26019 9404
rect 25961 9395 26019 9401
rect 26694 9392 26700 9404
rect 26752 9392 26758 9444
rect 28276 9432 28304 9463
rect 28534 9460 28540 9472
rect 28592 9460 28598 9512
rect 29914 9460 29920 9512
rect 29972 9500 29978 9512
rect 30377 9503 30435 9509
rect 30377 9500 30389 9503
rect 29972 9472 30389 9500
rect 29972 9460 29978 9472
rect 30377 9469 30389 9472
rect 30423 9469 30435 9503
rect 32416 9500 32444 9531
rect 32490 9528 32496 9580
rect 32548 9568 32554 9580
rect 35621 9571 35679 9577
rect 32548 9540 32593 9568
rect 32548 9528 32554 9540
rect 35621 9537 35633 9571
rect 35667 9568 35679 9571
rect 36446 9568 36452 9580
rect 35667 9540 36452 9568
rect 35667 9537 35679 9540
rect 35621 9531 35679 9537
rect 36446 9528 36452 9540
rect 36504 9528 36510 9580
rect 37384 9568 37412 9608
rect 37550 9596 37556 9608
rect 37608 9596 37614 9648
rect 37921 9639 37979 9645
rect 37921 9605 37933 9639
rect 37967 9636 37979 9639
rect 38580 9636 38608 9676
rect 39390 9664 39396 9676
rect 39448 9664 39454 9716
rect 37967 9608 38608 9636
rect 38648 9639 38706 9645
rect 37967 9605 37979 9608
rect 37921 9599 37979 9605
rect 38648 9605 38660 9639
rect 38694 9636 38706 9639
rect 38930 9636 38936 9648
rect 38694 9608 38936 9636
rect 38694 9605 38706 9608
rect 38648 9599 38706 9605
rect 38930 9596 38936 9608
rect 38988 9596 38994 9648
rect 37737 9571 37795 9577
rect 37737 9568 37749 9571
rect 37384 9540 37749 9568
rect 37737 9537 37749 9540
rect 37783 9568 37795 9571
rect 37783 9540 39804 9568
rect 37783 9537 37795 9540
rect 37737 9531 37795 9537
rect 32950 9500 32956 9512
rect 32416 9472 32956 9500
rect 30377 9463 30435 9469
rect 32950 9460 32956 9472
rect 33008 9460 33014 9512
rect 37918 9460 37924 9512
rect 37976 9500 37982 9512
rect 38381 9503 38439 9509
rect 38381 9500 38393 9503
rect 37976 9472 38393 9500
rect 37976 9460 37982 9472
rect 38381 9469 38393 9472
rect 38427 9469 38439 9503
rect 38381 9463 38439 9469
rect 28718 9432 28724 9444
rect 28276 9404 28724 9432
rect 28718 9392 28724 9404
rect 28776 9392 28782 9444
rect 39776 9441 39804 9540
rect 39761 9435 39819 9441
rect 39761 9401 39773 9435
rect 39807 9401 39819 9435
rect 39761 9395 39819 9401
rect 10318 9364 10324 9376
rect 8220 9336 10324 9364
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 10689 9367 10747 9373
rect 10689 9364 10701 9367
rect 10468 9336 10701 9364
rect 10468 9324 10474 9336
rect 10689 9333 10701 9336
rect 10735 9333 10747 9367
rect 12526 9364 12532 9376
rect 12487 9336 12532 9364
rect 10689 9327 10747 9333
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 12989 9367 13047 9373
rect 12989 9333 13001 9367
rect 13035 9364 13047 9367
rect 13170 9364 13176 9376
rect 13035 9336 13176 9364
rect 13035 9333 13047 9336
rect 12989 9327 13047 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 14366 9364 14372 9376
rect 14327 9336 14372 9364
rect 14366 9324 14372 9336
rect 14424 9324 14430 9376
rect 15289 9367 15347 9373
rect 15289 9333 15301 9367
rect 15335 9364 15347 9367
rect 15562 9364 15568 9376
rect 15335 9336 15568 9364
rect 15335 9333 15347 9336
rect 15289 9327 15347 9333
rect 15562 9324 15568 9336
rect 15620 9324 15626 9376
rect 15841 9367 15899 9373
rect 15841 9333 15853 9367
rect 15887 9364 15899 9367
rect 15930 9364 15936 9376
rect 15887 9336 15936 9364
rect 15887 9333 15899 9336
rect 15841 9327 15899 9333
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16761 9367 16819 9373
rect 16761 9333 16773 9367
rect 16807 9364 16819 9367
rect 17218 9364 17224 9376
rect 16807 9336 17224 9364
rect 16807 9333 16819 9336
rect 16761 9327 16819 9333
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 17862 9364 17868 9376
rect 17823 9336 17868 9364
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 18506 9364 18512 9376
rect 18467 9336 18512 9364
rect 18506 9324 18512 9336
rect 18564 9324 18570 9376
rect 32769 9367 32827 9373
rect 32769 9333 32781 9367
rect 32815 9364 32827 9367
rect 33594 9364 33600 9376
rect 32815 9336 33600 9364
rect 32815 9333 32827 9336
rect 32769 9327 32827 9333
rect 33594 9324 33600 9336
rect 33652 9324 33658 9376
rect 35253 9367 35311 9373
rect 35253 9333 35265 9367
rect 35299 9364 35311 9367
rect 35342 9364 35348 9376
rect 35299 9336 35348 9364
rect 35299 9333 35311 9336
rect 35253 9327 35311 9333
rect 35342 9324 35348 9336
rect 35400 9324 35406 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 6638 9120 6644 9172
rect 6696 9160 6702 9172
rect 7469 9163 7527 9169
rect 7469 9160 7481 9163
rect 6696 9132 7481 9160
rect 6696 9120 6702 9132
rect 7469 9129 7481 9132
rect 7515 9160 7527 9163
rect 10226 9160 10232 9172
rect 7515 9132 9996 9160
rect 10139 9132 10232 9160
rect 7515 9129 7527 9132
rect 7469 9123 7527 9129
rect 4706 9092 4712 9104
rect 4667 9064 4712 9092
rect 4706 9052 4712 9064
rect 4764 9052 4770 9104
rect 9858 9092 9864 9104
rect 8956 9064 9864 9092
rect 2501 9027 2559 9033
rect 2501 8993 2513 9027
rect 2547 9024 2559 9027
rect 2866 9024 2872 9036
rect 2547 8996 2872 9024
rect 2547 8993 2559 8996
rect 2501 8987 2559 8993
rect 2866 8984 2872 8996
rect 2924 9024 2930 9036
rect 3970 9024 3976 9036
rect 2924 8996 3976 9024
rect 2924 8984 2930 8996
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 5258 8984 5264 9036
rect 5316 9024 5322 9036
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 5316 8996 5457 9024
rect 5316 8984 5322 8996
rect 5445 8993 5457 8996
rect 5491 8993 5503 9027
rect 5445 8987 5503 8993
rect 2314 8956 2320 8968
rect 2275 8928 2320 8956
rect 2314 8916 2320 8928
rect 2372 8916 2378 8968
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 5040 8928 5181 8956
rect 5040 8916 5046 8928
rect 5169 8925 5181 8928
rect 5215 8925 5227 8959
rect 5169 8919 5227 8925
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8956 6975 8959
rect 7006 8956 7012 8968
rect 6963 8928 7012 8956
rect 6963 8925 6975 8928
rect 6917 8919 6975 8925
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 8956 8965 8984 9064
rect 9858 9052 9864 9064
rect 9916 9052 9922 9104
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 9048 8996 9229 9024
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 4525 8891 4583 8897
rect 4525 8857 4537 8891
rect 4571 8888 4583 8891
rect 4614 8888 4620 8900
rect 4571 8860 4620 8888
rect 4571 8857 4583 8860
rect 4525 8851 4583 8857
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 6270 8848 6276 8900
rect 6328 8888 6334 8900
rect 9048 8888 9076 8996
rect 9217 8993 9229 8996
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 9309 9027 9367 9033
rect 9309 8993 9321 9027
rect 9355 9024 9367 9027
rect 9766 9024 9772 9036
rect 9355 8996 9772 9024
rect 9355 8993 9367 8996
rect 9309 8987 9367 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 9968 9024 9996 9132
rect 10226 9120 10232 9132
rect 10284 9160 10290 9172
rect 20622 9160 20628 9172
rect 10284 9132 20208 9160
rect 20535 9132 20628 9160
rect 10284 9120 10290 9132
rect 10318 9052 10324 9104
rect 10376 9092 10382 9104
rect 13357 9095 13415 9101
rect 10376 9064 12434 9092
rect 10376 9052 10382 9064
rect 11238 9024 11244 9036
rect 9968 8996 11244 9024
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 11882 9024 11888 9036
rect 11348 8996 11888 9024
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9490 8956 9496 8968
rect 9451 8928 9496 8956
rect 9125 8919 9183 8925
rect 6328 8860 9076 8888
rect 9140 8888 9168 8919
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 9858 8916 9864 8968
rect 9916 8956 9922 8968
rect 11348 8965 11376 8996
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 12406 9024 12434 9064
rect 13357 9061 13369 9095
rect 13403 9092 13415 9095
rect 14182 9092 14188 9104
rect 13403 9064 14188 9092
rect 13403 9061 13415 9064
rect 13357 9055 13415 9061
rect 14182 9052 14188 9064
rect 14240 9052 14246 9104
rect 16114 9092 16120 9104
rect 16027 9064 16120 9092
rect 16114 9052 16120 9064
rect 16172 9092 16178 9104
rect 17034 9092 17040 9104
rect 16172 9064 17040 9092
rect 16172 9052 16178 9064
rect 17034 9052 17040 9064
rect 17092 9052 17098 9104
rect 18690 9092 18696 9104
rect 18651 9064 18696 9092
rect 18690 9052 18696 9064
rect 18748 9052 18754 9104
rect 20180 9092 20208 9132
rect 20622 9120 20628 9132
rect 20680 9160 20686 9172
rect 25406 9160 25412 9172
rect 20680 9132 25412 9160
rect 20680 9120 20686 9132
rect 25406 9120 25412 9132
rect 25464 9120 25470 9172
rect 28905 9163 28963 9169
rect 28905 9129 28917 9163
rect 28951 9160 28963 9163
rect 30466 9160 30472 9172
rect 28951 9132 30472 9160
rect 28951 9129 28963 9132
rect 28905 9123 28963 9129
rect 30466 9120 30472 9132
rect 30524 9120 30530 9172
rect 31846 9120 31852 9172
rect 31904 9160 31910 9172
rect 32677 9163 32735 9169
rect 32677 9160 32689 9163
rect 31904 9132 32689 9160
rect 31904 9120 31910 9132
rect 32677 9129 32689 9132
rect 32723 9129 32735 9163
rect 33686 9160 33692 9172
rect 33647 9132 33692 9160
rect 32677 9123 32735 9129
rect 33686 9120 33692 9132
rect 33744 9120 33750 9172
rect 35802 9120 35808 9172
rect 35860 9160 35866 9172
rect 36081 9163 36139 9169
rect 36081 9160 36093 9163
rect 35860 9132 36093 9160
rect 35860 9120 35866 9132
rect 36081 9129 36093 9132
rect 36127 9129 36139 9163
rect 36081 9123 36139 9129
rect 22554 9092 22560 9104
rect 20180 9064 22560 9092
rect 22554 9052 22560 9064
rect 22612 9052 22618 9104
rect 28534 9052 28540 9104
rect 28592 9092 28598 9104
rect 28592 9064 32444 9092
rect 28592 9052 28598 9064
rect 12989 9027 13047 9033
rect 12989 9024 13001 9027
rect 12406 8996 13001 9024
rect 12989 8993 13001 8996
rect 13035 8993 13047 9027
rect 12989 8987 13047 8993
rect 15473 9027 15531 9033
rect 15473 8993 15485 9027
rect 15519 9024 15531 9027
rect 16850 9024 16856 9036
rect 15519 8996 16856 9024
rect 15519 8993 15531 8996
rect 15473 8987 15531 8993
rect 16850 8984 16856 8996
rect 16908 9024 16914 9036
rect 17313 9027 17371 9033
rect 17313 9024 17325 9027
rect 16908 8996 17325 9024
rect 16908 8984 16914 8996
rect 17313 8993 17325 8996
rect 17359 8993 17371 9027
rect 17313 8987 17371 8993
rect 21177 9027 21235 9033
rect 21177 8993 21189 9027
rect 21223 9024 21235 9027
rect 21818 9024 21824 9036
rect 21223 8996 21824 9024
rect 21223 8993 21235 8996
rect 21177 8987 21235 8993
rect 21818 8984 21824 8996
rect 21876 9024 21882 9036
rect 21913 9027 21971 9033
rect 21913 9024 21925 9027
rect 21876 8996 21925 9024
rect 21876 8984 21882 8996
rect 21913 8993 21925 8996
rect 21959 8993 21971 9027
rect 22186 9024 22192 9036
rect 22147 8996 22192 9024
rect 21913 8987 21971 8993
rect 22186 8984 22192 8996
rect 22244 8984 22250 9036
rect 32416 9024 32444 9064
rect 34698 9024 34704 9036
rect 32416 8996 33548 9024
rect 34659 8996 34704 9024
rect 11149 8959 11207 8965
rect 11149 8956 11161 8959
rect 9916 8928 11161 8956
rect 9916 8916 9922 8928
rect 11149 8925 11161 8928
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 11333 8959 11391 8965
rect 11333 8925 11345 8959
rect 11379 8925 11391 8959
rect 11333 8919 11391 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8925 11575 8959
rect 11517 8919 11575 8925
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8956 11759 8959
rect 13170 8956 13176 8968
rect 11747 8928 12434 8956
rect 13131 8928 13176 8956
rect 11747 8925 11759 8928
rect 11701 8919 11759 8925
rect 10226 8888 10232 8900
rect 9140 8860 10232 8888
rect 6328 8848 6334 8860
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 11238 8848 11244 8900
rect 11296 8888 11302 8900
rect 11440 8888 11468 8919
rect 11296 8860 11468 8888
rect 11296 8848 11302 8860
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 1670 8780 1676 8832
rect 1728 8820 1734 8832
rect 2133 8823 2191 8829
rect 2133 8820 2145 8823
rect 1728 8792 2145 8820
rect 1728 8780 1734 8792
rect 2133 8789 2145 8792
rect 2179 8789 2191 8823
rect 2133 8783 2191 8789
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 3053 8823 3111 8829
rect 3053 8820 3065 8823
rect 2832 8792 3065 8820
rect 2832 8780 2838 8792
rect 3053 8789 3065 8792
rect 3099 8789 3111 8823
rect 3878 8820 3884 8832
rect 3839 8792 3884 8820
rect 3053 8783 3111 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 6733 8823 6791 8829
rect 6733 8820 6745 8823
rect 6604 8792 6745 8820
rect 6604 8780 6610 8792
rect 6733 8789 6745 8792
rect 6779 8789 6791 8823
rect 6733 8783 6791 8789
rect 8021 8823 8079 8829
rect 8021 8789 8033 8823
rect 8067 8820 8079 8823
rect 8110 8820 8116 8832
rect 8067 8792 8116 8820
rect 8067 8789 8079 8792
rect 8021 8783 8079 8789
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 9674 8820 9680 8832
rect 9635 8792 9680 8820
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 11532 8820 11560 8919
rect 12406 8888 12434 8928
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 15206 8959 15264 8965
rect 15206 8956 15218 8959
rect 14424 8928 15218 8956
rect 14424 8916 14430 8928
rect 15206 8925 15218 8928
rect 15252 8925 15264 8959
rect 15930 8956 15936 8968
rect 15891 8928 15936 8956
rect 15206 8919 15264 8925
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 18966 8956 18972 8968
rect 16040 8928 18972 8956
rect 13446 8888 13452 8900
rect 12406 8860 13452 8888
rect 13446 8848 13452 8860
rect 13504 8848 13510 8900
rect 11882 8820 11888 8832
rect 9824 8792 11560 8820
rect 11843 8792 11888 8820
rect 9824 8780 9830 8792
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 13964 8792 14105 8820
rect 13964 8780 13970 8792
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14093 8783 14151 8789
rect 14182 8780 14188 8832
rect 14240 8820 14246 8832
rect 14458 8820 14464 8832
rect 14240 8792 14464 8820
rect 14240 8780 14246 8792
rect 14458 8780 14464 8792
rect 14516 8820 14522 8832
rect 16040 8820 16068 8928
rect 18966 8916 18972 8928
rect 19024 8916 19030 8968
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 19116 8928 19257 8956
rect 19116 8916 19122 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 20714 8916 20720 8968
rect 20772 8956 20778 8968
rect 21085 8959 21143 8965
rect 21085 8956 21097 8959
rect 20772 8928 21097 8956
rect 20772 8916 20778 8928
rect 21085 8925 21097 8928
rect 21131 8925 21143 8959
rect 21269 8959 21327 8965
rect 21269 8956 21281 8959
rect 21085 8919 21143 8925
rect 21192 8928 21281 8956
rect 21192 8900 21220 8928
rect 21269 8925 21281 8928
rect 21315 8925 21327 8959
rect 28350 8956 28356 8968
rect 28311 8928 28356 8956
rect 21269 8919 21327 8925
rect 28350 8916 28356 8928
rect 28408 8916 28414 8968
rect 28718 8956 28724 8968
rect 28679 8928 28724 8956
rect 28718 8916 28724 8928
rect 28776 8916 28782 8968
rect 31294 8916 31300 8968
rect 31352 8956 31358 8968
rect 32125 8959 32183 8965
rect 32125 8956 32137 8959
rect 31352 8928 32137 8956
rect 31352 8916 31358 8928
rect 32125 8925 32137 8928
rect 32171 8925 32183 8959
rect 32398 8956 32404 8968
rect 32359 8928 32404 8956
rect 32125 8919 32183 8925
rect 32398 8916 32404 8928
rect 32456 8916 32462 8968
rect 32508 8965 32536 8996
rect 32493 8959 32551 8965
rect 32493 8925 32505 8959
rect 32539 8956 32551 8959
rect 32674 8956 32680 8968
rect 32539 8928 32680 8956
rect 32539 8925 32551 8928
rect 32493 8919 32551 8925
rect 32674 8916 32680 8928
rect 32732 8916 32738 8968
rect 33134 8956 33140 8968
rect 33095 8928 33140 8956
rect 33134 8916 33140 8928
rect 33192 8916 33198 8968
rect 33410 8956 33416 8968
rect 33371 8928 33416 8956
rect 33410 8916 33416 8928
rect 33468 8916 33474 8968
rect 33520 8965 33548 8996
rect 34698 8984 34704 8996
rect 34756 8984 34762 9036
rect 33505 8959 33563 8965
rect 33505 8925 33517 8959
rect 33551 8925 33563 8959
rect 34716 8956 34744 8984
rect 37918 8956 37924 8968
rect 34716 8928 37924 8956
rect 33505 8919 33563 8925
rect 37918 8916 37924 8928
rect 37976 8916 37982 8968
rect 58158 8956 58164 8968
rect 58119 8928 58164 8956
rect 58158 8916 58164 8928
rect 58216 8916 58222 8968
rect 17310 8848 17316 8900
rect 17368 8888 17374 8900
rect 17558 8891 17616 8897
rect 17558 8888 17570 8891
rect 17368 8860 17570 8888
rect 17368 8848 17374 8860
rect 17558 8857 17570 8860
rect 17604 8857 17616 8891
rect 17558 8851 17616 8857
rect 19150 8848 19156 8900
rect 19208 8888 19214 8900
rect 19490 8891 19548 8897
rect 19490 8888 19502 8891
rect 19208 8860 19502 8888
rect 19208 8848 19214 8860
rect 19490 8857 19502 8860
rect 19536 8857 19548 8891
rect 19490 8851 19548 8857
rect 21174 8848 21180 8900
rect 21232 8848 21238 8900
rect 28166 8848 28172 8900
rect 28224 8888 28230 8900
rect 28537 8891 28595 8897
rect 28537 8888 28549 8891
rect 28224 8860 28549 8888
rect 28224 8848 28230 8860
rect 28537 8857 28549 8860
rect 28583 8857 28595 8891
rect 28537 8851 28595 8857
rect 28629 8891 28687 8897
rect 28629 8857 28641 8891
rect 28675 8888 28687 8891
rect 29730 8888 29736 8900
rect 28675 8860 29736 8888
rect 28675 8857 28687 8860
rect 28629 8851 28687 8857
rect 29730 8848 29736 8860
rect 29788 8848 29794 8900
rect 29914 8888 29920 8900
rect 29875 8860 29920 8888
rect 29914 8848 29920 8860
rect 29972 8848 29978 8900
rect 34974 8897 34980 8900
rect 32309 8891 32367 8897
rect 32309 8888 32321 8891
rect 30024 8860 32321 8888
rect 16666 8820 16672 8832
rect 14516 8792 16068 8820
rect 16627 8792 16672 8820
rect 14516 8780 14522 8792
rect 16666 8780 16672 8792
rect 16724 8780 16730 8832
rect 17034 8780 17040 8832
rect 17092 8820 17098 8832
rect 23382 8820 23388 8832
rect 17092 8792 23388 8820
rect 17092 8780 17098 8792
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 28442 8780 28448 8832
rect 28500 8820 28506 8832
rect 30024 8820 30052 8860
rect 32309 8857 32321 8860
rect 32355 8888 32367 8891
rect 33321 8891 33379 8897
rect 33321 8888 33333 8891
rect 32355 8860 33333 8888
rect 32355 8857 32367 8860
rect 32309 8851 32367 8857
rect 33321 8857 33333 8860
rect 33367 8857 33379 8891
rect 33321 8851 33379 8857
rect 34968 8851 34980 8897
rect 35032 8888 35038 8900
rect 35032 8860 35068 8888
rect 28500 8792 30052 8820
rect 28500 8780 28506 8792
rect 30926 8780 30932 8832
rect 30984 8820 30990 8832
rect 31205 8823 31263 8829
rect 31205 8820 31217 8823
rect 30984 8792 31217 8820
rect 30984 8780 30990 8792
rect 31205 8789 31217 8792
rect 31251 8789 31263 8823
rect 32324 8820 32352 8851
rect 34974 8848 34980 8851
rect 35032 8848 35038 8860
rect 36446 8848 36452 8900
rect 36504 8888 36510 8900
rect 37093 8891 37151 8897
rect 37093 8888 37105 8891
rect 36504 8860 37105 8888
rect 36504 8848 36510 8860
rect 37093 8857 37105 8860
rect 37139 8857 37151 8891
rect 37093 8851 37151 8857
rect 37277 8891 37335 8897
rect 37277 8857 37289 8891
rect 37323 8888 37335 8891
rect 37323 8860 37780 8888
rect 37323 8857 37335 8860
rect 37277 8851 37335 8857
rect 32490 8820 32496 8832
rect 32324 8792 32496 8820
rect 31205 8783 31263 8789
rect 32490 8780 32496 8792
rect 32548 8780 32554 8832
rect 36722 8780 36728 8832
rect 36780 8820 36786 8832
rect 37292 8820 37320 8851
rect 36780 8792 37320 8820
rect 37461 8823 37519 8829
rect 36780 8780 36786 8792
rect 37461 8789 37473 8823
rect 37507 8820 37519 8823
rect 37550 8820 37556 8832
rect 37507 8792 37556 8820
rect 37507 8789 37519 8792
rect 37461 8783 37519 8789
rect 37550 8780 37556 8792
rect 37608 8780 37614 8832
rect 37752 8820 37780 8860
rect 38010 8848 38016 8900
rect 38068 8888 38074 8900
rect 38166 8891 38224 8897
rect 38166 8888 38178 8891
rect 38068 8860 38178 8888
rect 38068 8848 38074 8860
rect 38166 8857 38178 8860
rect 38212 8857 38224 8891
rect 38166 8851 38224 8857
rect 39301 8823 39359 8829
rect 39301 8820 39313 8823
rect 37752 8792 39313 8820
rect 39301 8789 39313 8792
rect 39347 8789 39359 8823
rect 39301 8783 39359 8789
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 1673 8619 1731 8625
rect 1673 8585 1685 8619
rect 1719 8585 1731 8619
rect 7006 8616 7012 8628
rect 6967 8588 7012 8616
rect 1673 8579 1731 8585
rect 1688 8548 1716 8579
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 7558 8576 7564 8628
rect 7616 8616 7622 8628
rect 7616 8588 9812 8616
rect 7616 8576 7622 8588
rect 2378 8551 2436 8557
rect 2378 8548 2390 8551
rect 1688 8520 2390 8548
rect 2378 8517 2390 8520
rect 2424 8517 2436 8551
rect 2378 8511 2436 8517
rect 4614 8508 4620 8560
rect 4672 8548 4678 8560
rect 9674 8557 9680 8560
rect 9668 8548 9680 8557
rect 4672 8520 8064 8548
rect 9635 8520 9680 8548
rect 4672 8508 4678 8520
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8480 1547 8483
rect 1670 8480 1676 8492
rect 1535 8452 1676 8480
rect 1535 8449 1547 8452
rect 1489 8443 1547 8449
rect 1670 8440 1676 8452
rect 1728 8440 1734 8492
rect 5166 8440 5172 8492
rect 5224 8480 5230 8492
rect 6638 8480 6644 8492
rect 5224 8452 6644 8480
rect 5224 8440 5230 8452
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 7837 8483 7895 8489
rect 7837 8480 7849 8483
rect 6871 8452 7512 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 1854 8372 1860 8424
rect 1912 8412 1918 8424
rect 2133 8415 2191 8421
rect 2133 8412 2145 8415
rect 1912 8384 2145 8412
rect 1912 8372 1918 8384
rect 2133 8381 2145 8384
rect 2179 8381 2191 8415
rect 4982 8412 4988 8424
rect 4943 8384 4988 8412
rect 2133 8375 2191 8381
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 5261 8415 5319 8421
rect 5261 8381 5273 8415
rect 5307 8381 5319 8415
rect 5261 8375 5319 8381
rect 2866 8236 2872 8288
rect 2924 8276 2930 8288
rect 3513 8279 3571 8285
rect 3513 8276 3525 8279
rect 2924 8248 3525 8276
rect 2924 8236 2930 8248
rect 3513 8245 3525 8248
rect 3559 8245 3571 8279
rect 3970 8276 3976 8288
rect 3931 8248 3976 8276
rect 3513 8239 3571 8245
rect 3970 8236 3976 8248
rect 4028 8236 4034 8288
rect 5276 8276 5304 8375
rect 7484 8353 7512 8452
rect 7760 8452 7849 8480
rect 7469 8347 7527 8353
rect 7469 8313 7481 8347
rect 7515 8313 7527 8347
rect 7760 8344 7788 8452
rect 7837 8449 7849 8452
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 7926 8412 7932 8424
rect 7887 8384 7932 8412
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 8036 8421 8064 8520
rect 9668 8511 9680 8520
rect 9674 8508 9680 8511
rect 9732 8508 9738 8560
rect 9784 8548 9812 8588
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11296 8588 12173 8616
rect 11296 8576 11302 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 16850 8616 16856 8628
rect 13780 8588 16856 8616
rect 13780 8576 13786 8588
rect 16850 8576 16856 8588
rect 16908 8576 16914 8628
rect 17310 8616 17316 8628
rect 17271 8588 17316 8616
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 19061 8619 19119 8625
rect 17420 8588 18920 8616
rect 11514 8548 11520 8560
rect 9784 8520 11520 8548
rect 11514 8508 11520 8520
rect 11572 8508 11578 8560
rect 12989 8551 13047 8557
rect 12989 8517 13001 8551
rect 13035 8548 13047 8551
rect 13814 8548 13820 8560
rect 13035 8520 13820 8548
rect 13035 8517 13047 8520
rect 12989 8511 13047 8517
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 16758 8548 16764 8560
rect 16719 8520 16764 8548
rect 16758 8508 16764 8520
rect 16816 8548 16822 8560
rect 17420 8548 17448 8588
rect 16816 8520 17448 8548
rect 17696 8520 18736 8548
rect 16816 8508 16822 8520
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 9398 8480 9404 8492
rect 8904 8452 9404 8480
rect 8904 8440 8910 8452
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 11885 8483 11943 8489
rect 9548 8452 10824 8480
rect 9548 8440 9554 8452
rect 8021 8415 8079 8421
rect 8021 8381 8033 8415
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 10796 8353 10824 8452
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 13906 8480 13912 8492
rect 11931 8452 13912 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 13906 8440 13912 8452
rect 13964 8440 13970 8492
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8449 14059 8483
rect 14734 8480 14740 8492
rect 14695 8452 14740 8480
rect 14001 8443 14059 8449
rect 11974 8412 11980 8424
rect 11935 8384 11980 8412
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 14016 8412 14044 8443
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 17494 8480 17500 8492
rect 16040 8452 17500 8480
rect 16040 8421 16068 8452
rect 17494 8440 17500 8452
rect 17552 8489 17558 8492
rect 17696 8489 17724 8520
rect 17552 8483 17601 8489
rect 17552 8449 17555 8483
rect 17589 8449 17601 8483
rect 17552 8443 17601 8449
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 17773 8483 17831 8489
rect 17773 8449 17785 8483
rect 17819 8449 17831 8483
rect 17954 8480 17960 8492
rect 17915 8452 17960 8480
rect 17773 8443 17831 8449
rect 17552 8440 17558 8443
rect 16025 8415 16083 8421
rect 16025 8412 16037 8415
rect 13556 8384 14044 8412
rect 14200 8384 16037 8412
rect 13556 8356 13584 8384
rect 8757 8347 8815 8353
rect 8757 8344 8769 8347
rect 7760 8316 8769 8344
rect 7469 8307 7527 8313
rect 8757 8313 8769 8316
rect 8803 8344 8815 8347
rect 10781 8347 10839 8353
rect 8803 8316 9444 8344
rect 8803 8313 8815 8316
rect 8757 8307 8815 8313
rect 5534 8276 5540 8288
rect 5276 8248 5540 8276
rect 5534 8236 5540 8248
rect 5592 8276 5598 8288
rect 7558 8276 7564 8288
rect 5592 8248 7564 8276
rect 5592 8236 5598 8248
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 9416 8276 9444 8316
rect 10781 8313 10793 8347
rect 10827 8344 10839 8347
rect 11698 8344 11704 8356
rect 10827 8316 11704 8344
rect 10827 8313 10839 8316
rect 10781 8307 10839 8313
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 13538 8344 13544 8356
rect 13499 8316 13544 8344
rect 13538 8304 13544 8316
rect 13596 8304 13602 8356
rect 14200 8344 14228 8384
rect 16025 8381 16037 8384
rect 16071 8381 16083 8415
rect 17788 8412 17816 8443
rect 17954 8440 17960 8452
rect 18012 8480 18018 8492
rect 18417 8483 18475 8489
rect 18417 8480 18429 8483
rect 18012 8452 18429 8480
rect 18012 8440 18018 8452
rect 18417 8449 18429 8452
rect 18463 8449 18475 8483
rect 18598 8480 18604 8492
rect 18559 8452 18604 8480
rect 18417 8443 18475 8449
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 18708 8489 18736 8520
rect 18693 8483 18751 8489
rect 18693 8449 18705 8483
rect 18739 8449 18751 8483
rect 18693 8443 18751 8449
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8480 18843 8483
rect 18892 8480 18920 8588
rect 19061 8585 19073 8619
rect 19107 8616 19119 8619
rect 19150 8616 19156 8628
rect 19107 8588 19156 8616
rect 19107 8585 19119 8588
rect 19061 8579 19119 8585
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 27709 8619 27767 8625
rect 27709 8585 27721 8619
rect 27755 8616 27767 8619
rect 29549 8619 29607 8625
rect 27755 8588 29224 8616
rect 27755 8585 27767 8588
rect 27709 8579 27767 8585
rect 19521 8551 19579 8557
rect 19521 8548 19533 8551
rect 19306 8520 19533 8548
rect 18831 8452 19012 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 18322 8412 18328 8424
rect 17788 8384 18328 8412
rect 16025 8375 16083 8381
rect 18322 8372 18328 8384
rect 18380 8372 18386 8424
rect 18708 8412 18736 8443
rect 18874 8412 18880 8424
rect 18708 8384 18880 8412
rect 18874 8372 18880 8384
rect 18932 8372 18938 8424
rect 18984 8412 19012 8452
rect 19150 8440 19156 8492
rect 19208 8480 19214 8492
rect 19306 8480 19334 8520
rect 19521 8517 19533 8520
rect 19567 8517 19579 8551
rect 19521 8511 19579 8517
rect 19705 8551 19763 8557
rect 19705 8517 19717 8551
rect 19751 8548 19763 8551
rect 20622 8548 20628 8560
rect 19751 8520 20628 8548
rect 19751 8517 19763 8520
rect 19705 8511 19763 8517
rect 20622 8508 20628 8520
rect 20680 8508 20686 8560
rect 24210 8548 24216 8560
rect 23860 8520 24216 8548
rect 19208 8452 19334 8480
rect 19208 8440 19214 8452
rect 19426 8440 19432 8492
rect 19484 8480 19490 8492
rect 19889 8483 19947 8489
rect 19889 8480 19901 8483
rect 19484 8452 19901 8480
rect 19484 8440 19490 8452
rect 19889 8449 19901 8452
rect 19935 8449 19947 8483
rect 21818 8480 21824 8492
rect 21779 8452 21824 8480
rect 19889 8443 19947 8449
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 22097 8483 22155 8489
rect 22097 8449 22109 8483
rect 22143 8480 22155 8483
rect 22830 8480 22836 8492
rect 22143 8452 22836 8480
rect 22143 8449 22155 8452
rect 22097 8443 22155 8449
rect 22830 8440 22836 8452
rect 22888 8480 22894 8492
rect 23014 8480 23020 8492
rect 22888 8452 23020 8480
rect 22888 8440 22894 8452
rect 23014 8440 23020 8452
rect 23072 8440 23078 8492
rect 23382 8440 23388 8492
rect 23440 8480 23446 8492
rect 23860 8489 23888 8520
rect 24210 8508 24216 8520
rect 24268 8508 24274 8560
rect 27341 8551 27399 8557
rect 27341 8517 27353 8551
rect 27387 8548 27399 8551
rect 29196 8548 29224 8588
rect 29549 8585 29561 8619
rect 29595 8616 29607 8619
rect 29730 8616 29736 8628
rect 29595 8588 29736 8616
rect 29595 8585 29607 8588
rect 29549 8579 29607 8585
rect 29730 8576 29736 8588
rect 29788 8576 29794 8628
rect 32766 8576 32772 8628
rect 32824 8616 32830 8628
rect 32861 8619 32919 8625
rect 32861 8616 32873 8619
rect 32824 8588 32873 8616
rect 32824 8576 32830 8588
rect 32861 8585 32873 8588
rect 32907 8585 32919 8619
rect 32861 8579 32919 8585
rect 34885 8619 34943 8625
rect 34885 8585 34897 8619
rect 34931 8616 34943 8619
rect 34974 8616 34980 8628
rect 34931 8588 34980 8616
rect 34931 8585 34943 8588
rect 34885 8579 34943 8585
rect 34974 8576 34980 8588
rect 35032 8576 35038 8628
rect 38010 8616 38016 8628
rect 37971 8588 38016 8616
rect 38010 8576 38016 8588
rect 38068 8576 38074 8628
rect 30558 8548 30564 8560
rect 27387 8520 28488 8548
rect 29196 8520 30564 8548
rect 27387 8517 27399 8520
rect 27341 8511 27399 8517
rect 28460 8492 28488 8520
rect 30558 8508 30564 8520
rect 30616 8508 30622 8560
rect 30650 8508 30656 8560
rect 30708 8557 30714 8560
rect 30708 8548 30720 8557
rect 32582 8548 32588 8560
rect 30708 8520 30753 8548
rect 32543 8520 32588 8548
rect 30708 8511 30720 8520
rect 30708 8508 30714 8511
rect 32582 8508 32588 8520
rect 32640 8508 32646 8560
rect 35802 8548 35808 8560
rect 35268 8520 35808 8548
rect 23753 8483 23811 8489
rect 23753 8480 23765 8483
rect 23440 8452 23765 8480
rect 23440 8440 23446 8452
rect 23753 8449 23765 8452
rect 23799 8449 23811 8483
rect 23753 8443 23811 8449
rect 23845 8483 23903 8489
rect 23845 8449 23857 8483
rect 23891 8449 23903 8483
rect 23845 8443 23903 8449
rect 20070 8412 20076 8424
rect 18984 8384 20076 8412
rect 20070 8372 20076 8384
rect 20128 8372 20134 8424
rect 20993 8415 21051 8421
rect 20993 8381 21005 8415
rect 21039 8412 21051 8415
rect 21082 8412 21088 8424
rect 21039 8384 21088 8412
rect 21039 8381 21051 8384
rect 20993 8375 21051 8381
rect 21082 8372 21088 8384
rect 21140 8372 21146 8424
rect 14016 8316 14228 8344
rect 9582 8276 9588 8288
rect 9416 8248 9588 8276
rect 9582 8236 9588 8248
rect 9640 8236 9646 8288
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 14016 8276 14044 8316
rect 15010 8304 15016 8356
rect 15068 8344 15074 8356
rect 15473 8347 15531 8353
rect 15473 8344 15485 8347
rect 15068 8316 15485 8344
rect 15068 8304 15074 8316
rect 15473 8313 15485 8316
rect 15519 8313 15531 8347
rect 15473 8307 15531 8313
rect 18966 8304 18972 8356
rect 19024 8344 19030 8356
rect 23382 8344 23388 8356
rect 19024 8316 23388 8344
rect 19024 8304 19030 8316
rect 23382 8304 23388 8316
rect 23440 8304 23446 8356
rect 23768 8344 23796 8443
rect 23934 8440 23940 8492
rect 23992 8480 23998 8492
rect 24121 8483 24179 8489
rect 23992 8452 24037 8480
rect 23992 8440 23998 8452
rect 24121 8449 24133 8483
rect 24167 8480 24179 8483
rect 24578 8480 24584 8492
rect 24167 8452 24584 8480
rect 24167 8449 24179 8452
rect 24121 8443 24179 8449
rect 24578 8440 24584 8452
rect 24636 8440 24642 8492
rect 26326 8440 26332 8492
rect 26384 8480 26390 8492
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 26384 8452 27169 8480
rect 26384 8440 26390 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 27430 8480 27436 8492
rect 27391 8452 27436 8480
rect 27157 8443 27215 8449
rect 27430 8440 27436 8452
rect 27488 8440 27494 8492
rect 27525 8483 27583 8489
rect 27525 8449 27537 8483
rect 27571 8480 27583 8483
rect 28442 8480 28448 8492
rect 27571 8452 28304 8480
rect 28403 8452 28448 8480
rect 27571 8449 27583 8452
rect 27525 8443 27583 8449
rect 28166 8412 28172 8424
rect 28127 8384 28172 8412
rect 28166 8372 28172 8384
rect 28224 8372 28230 8424
rect 28276 8412 28304 8452
rect 28442 8440 28448 8452
rect 28500 8440 28506 8492
rect 32309 8483 32367 8489
rect 28644 8452 31754 8480
rect 28534 8412 28540 8424
rect 28276 8384 28540 8412
rect 28534 8372 28540 8384
rect 28592 8372 28598 8424
rect 26786 8344 26792 8356
rect 23768 8316 26792 8344
rect 26786 8304 26792 8316
rect 26844 8344 26850 8356
rect 28644 8344 28672 8452
rect 30926 8412 30932 8424
rect 30887 8384 30932 8412
rect 30926 8372 30932 8384
rect 30984 8372 30990 8424
rect 31726 8412 31754 8452
rect 32309 8449 32321 8483
rect 32355 8480 32367 8483
rect 32398 8480 32404 8492
rect 32355 8452 32404 8480
rect 32355 8449 32367 8452
rect 32309 8443 32367 8449
rect 32398 8440 32404 8452
rect 32456 8440 32462 8492
rect 32490 8440 32496 8492
rect 32548 8480 32554 8492
rect 32548 8452 32593 8480
rect 32548 8440 32554 8452
rect 32674 8440 32680 8492
rect 32732 8480 32738 8492
rect 35268 8489 35296 8520
rect 35802 8508 35808 8520
rect 35860 8548 35866 8560
rect 38378 8548 38384 8560
rect 35860 8520 38384 8548
rect 35860 8508 35866 8520
rect 35161 8483 35219 8489
rect 32732 8452 32777 8480
rect 32732 8440 32738 8452
rect 35161 8449 35173 8483
rect 35207 8449 35219 8483
rect 35161 8443 35219 8449
rect 35253 8483 35311 8489
rect 35253 8449 35265 8483
rect 35299 8449 35311 8483
rect 35253 8443 35311 8449
rect 34333 8415 34391 8421
rect 34333 8412 34345 8415
rect 31726 8384 34345 8412
rect 34333 8381 34345 8384
rect 34379 8412 34391 8415
rect 35176 8412 35204 8443
rect 35342 8440 35348 8492
rect 35400 8480 35406 8492
rect 35400 8452 35445 8480
rect 35400 8440 35406 8452
rect 35526 8440 35532 8492
rect 35584 8480 35590 8492
rect 37369 8483 37427 8489
rect 37369 8480 37381 8483
rect 35584 8452 37381 8480
rect 35584 8440 35590 8452
rect 37369 8449 37381 8452
rect 37415 8449 37427 8483
rect 37550 8480 37556 8492
rect 37511 8452 37556 8480
rect 37369 8443 37427 8449
rect 37550 8440 37556 8452
rect 37608 8440 37614 8492
rect 37660 8489 37688 8520
rect 38378 8508 38384 8520
rect 38436 8508 38442 8560
rect 37645 8483 37703 8489
rect 37645 8449 37657 8483
rect 37691 8449 37703 8483
rect 37645 8443 37703 8449
rect 37734 8440 37740 8492
rect 37792 8480 37798 8492
rect 37792 8452 37837 8480
rect 37792 8440 37798 8452
rect 35618 8412 35624 8424
rect 34379 8384 35624 8412
rect 34379 8381 34391 8384
rect 34333 8375 34391 8381
rect 35618 8372 35624 8384
rect 35676 8372 35682 8424
rect 26844 8316 28672 8344
rect 26844 8304 26850 8316
rect 14182 8276 14188 8288
rect 9824 8248 14044 8276
rect 14143 8248 14188 8276
rect 9824 8236 9830 8248
rect 14182 8236 14188 8248
rect 14240 8236 14246 8288
rect 14918 8276 14924 8288
rect 14831 8248 14924 8276
rect 14918 8236 14924 8248
rect 14976 8276 14982 8288
rect 18230 8276 18236 8288
rect 14976 8248 18236 8276
rect 14976 8236 14982 8248
rect 18230 8236 18236 8248
rect 18288 8236 18294 8288
rect 18598 8236 18604 8288
rect 18656 8276 18662 8288
rect 19150 8276 19156 8288
rect 18656 8248 19156 8276
rect 18656 8236 18662 8248
rect 19150 8236 19156 8248
rect 19208 8236 19214 8288
rect 23477 8279 23535 8285
rect 23477 8245 23489 8279
rect 23523 8276 23535 8279
rect 23566 8276 23572 8288
rect 23523 8248 23572 8276
rect 23523 8245 23535 8248
rect 23477 8239 23535 8245
rect 23566 8236 23572 8248
rect 23624 8236 23630 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 2314 8032 2320 8084
rect 2372 8072 2378 8084
rect 2409 8075 2467 8081
rect 2409 8072 2421 8075
rect 2372 8044 2421 8072
rect 2372 8032 2378 8044
rect 2409 8041 2421 8044
rect 2455 8041 2467 8075
rect 5350 8072 5356 8084
rect 5263 8044 5356 8072
rect 2409 8035 2467 8041
rect 5350 8032 5356 8044
rect 5408 8072 5414 8084
rect 7282 8072 7288 8084
rect 5408 8044 7288 8072
rect 5408 8032 5414 8044
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7653 8075 7711 8081
rect 7653 8041 7665 8075
rect 7699 8072 7711 8075
rect 7926 8072 7932 8084
rect 7699 8044 7932 8072
rect 7699 8041 7711 8044
rect 7653 8035 7711 8041
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9490 8072 9496 8084
rect 8352 8044 9496 8072
rect 8352 8032 8358 8044
rect 9490 8032 9496 8044
rect 9548 8072 9554 8084
rect 16574 8072 16580 8084
rect 9548 8044 16580 8072
rect 9548 8032 9554 8044
rect 16574 8032 16580 8044
rect 16632 8032 16638 8084
rect 18322 8072 18328 8084
rect 18283 8044 18328 8072
rect 18322 8032 18328 8044
rect 18380 8032 18386 8084
rect 23934 8032 23940 8084
rect 23992 8072 23998 8084
rect 24397 8075 24455 8081
rect 24397 8072 24409 8075
rect 23992 8044 24409 8072
rect 23992 8032 23998 8044
rect 24397 8041 24409 8044
rect 24443 8041 24455 8075
rect 24397 8035 24455 8041
rect 26234 8032 26240 8084
rect 26292 8072 26298 8084
rect 26697 8075 26755 8081
rect 26697 8072 26709 8075
rect 26292 8044 26709 8072
rect 26292 8032 26298 8044
rect 26697 8041 26709 8044
rect 26743 8072 26755 8075
rect 27430 8072 27436 8084
rect 26743 8044 27436 8072
rect 26743 8041 26755 8044
rect 26697 8035 26755 8041
rect 27430 8032 27436 8044
rect 27488 8032 27494 8084
rect 28994 8072 29000 8084
rect 28955 8044 29000 8072
rect 28994 8032 29000 8044
rect 29052 8032 29058 8084
rect 31573 8075 31631 8081
rect 31573 8041 31585 8075
rect 31619 8072 31631 8075
rect 32306 8072 32312 8084
rect 31619 8044 32312 8072
rect 31619 8041 31631 8044
rect 31573 8035 31631 8041
rect 32306 8032 32312 8044
rect 32364 8032 32370 8084
rect 37277 8075 37335 8081
rect 37277 8041 37289 8075
rect 37323 8072 37335 8075
rect 37734 8072 37740 8084
rect 37323 8044 37740 8072
rect 37323 8041 37335 8044
rect 37277 8035 37335 8041
rect 2884 7976 4200 8004
rect 2884 7948 2912 7976
rect 2866 7936 2872 7948
rect 2827 7908 2872 7936
rect 2866 7896 2872 7908
rect 2924 7896 2930 7948
rect 4172 7945 4200 7976
rect 9398 7964 9404 8016
rect 9456 8004 9462 8016
rect 11517 8007 11575 8013
rect 11517 8004 11529 8007
rect 9456 7976 11529 8004
rect 9456 7964 9462 7976
rect 11517 7973 11529 7976
rect 11563 8004 11575 8007
rect 12066 8004 12072 8016
rect 11563 7976 12072 8004
rect 11563 7973 11575 7976
rect 11517 7967 11575 7973
rect 12066 7964 12072 7976
rect 12124 7964 12130 8016
rect 26344 7976 28948 8004
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 4157 7939 4215 7945
rect 4157 7905 4169 7939
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 4525 7939 4583 7945
rect 4525 7905 4537 7939
rect 4571 7936 4583 7939
rect 5534 7936 5540 7948
rect 4571 7908 5540 7936
rect 4571 7905 4583 7908
rect 4525 7899 4583 7905
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2958 7868 2964 7880
rect 2823 7840 2964 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 3068 7800 3096 7899
rect 5534 7896 5540 7908
rect 5592 7896 5598 7948
rect 18046 7896 18052 7948
rect 18104 7936 18110 7948
rect 19797 7939 19855 7945
rect 19797 7936 19809 7939
rect 18104 7908 19809 7936
rect 18104 7896 18110 7908
rect 19797 7905 19809 7908
rect 19843 7905 19855 7939
rect 19797 7899 19855 7905
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 5626 7868 5632 7880
rect 4111 7840 5632 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 6270 7868 6276 7880
rect 6231 7840 6276 7868
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6546 7877 6552 7880
rect 6540 7868 6552 7877
rect 6507 7840 6552 7868
rect 6540 7831 6552 7840
rect 6546 7828 6552 7831
rect 6604 7828 6610 7880
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 8205 7871 8263 7877
rect 8205 7868 8217 7871
rect 7156 7840 8217 7868
rect 7156 7828 7162 7840
rect 8205 7837 8217 7840
rect 8251 7868 8263 7871
rect 12989 7871 13047 7877
rect 8251 7840 12434 7868
rect 8251 7837 8263 7840
rect 8205 7831 8263 7837
rect 4614 7800 4620 7812
rect 3068 7772 4620 7800
rect 4614 7760 4620 7772
rect 4672 7760 4678 7812
rect 4982 7760 4988 7812
rect 5040 7800 5046 7812
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 5040 7772 5273 7800
rect 5040 7760 5046 7772
rect 5261 7769 5273 7772
rect 5307 7769 5319 7803
rect 10229 7803 10287 7809
rect 10229 7800 10241 7803
rect 5261 7763 5319 7769
rect 9692 7772 10241 7800
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 1857 7735 1915 7741
rect 1857 7732 1869 7735
rect 1820 7704 1869 7732
rect 1820 7692 1826 7704
rect 1857 7701 1869 7704
rect 1903 7701 1915 7735
rect 1857 7695 1915 7701
rect 3881 7735 3939 7741
rect 3881 7701 3893 7735
rect 3927 7732 3939 7735
rect 3970 7732 3976 7744
rect 3927 7704 3976 7732
rect 3927 7701 3939 7704
rect 3881 7695 3939 7701
rect 3970 7692 3976 7704
rect 4028 7692 4034 7744
rect 9214 7732 9220 7744
rect 9175 7704 9220 7732
rect 9214 7692 9220 7704
rect 9272 7692 9278 7744
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 9692 7741 9720 7772
rect 10229 7769 10241 7772
rect 10275 7769 10287 7803
rect 12406 7800 12434 7840
rect 12989 7837 13001 7871
rect 13035 7868 13047 7871
rect 15102 7868 15108 7880
rect 13035 7840 15108 7868
rect 13035 7837 13047 7840
rect 12989 7831 13047 7837
rect 15102 7828 15108 7840
rect 15160 7828 15166 7880
rect 15381 7871 15439 7877
rect 15381 7837 15393 7871
rect 15427 7868 15439 7871
rect 19058 7868 19064 7880
rect 15427 7840 19064 7868
rect 15427 7837 15439 7840
rect 15381 7831 15439 7837
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 23566 7828 23572 7880
rect 23624 7877 23630 7880
rect 23624 7868 23636 7877
rect 23845 7871 23903 7877
rect 23624 7840 23669 7868
rect 23624 7831 23636 7840
rect 23845 7837 23857 7871
rect 23891 7868 23903 7871
rect 25130 7868 25136 7880
rect 23891 7840 25136 7868
rect 23891 7837 23903 7840
rect 23845 7831 23903 7837
rect 23624 7828 23630 7831
rect 25130 7828 25136 7840
rect 25188 7868 25194 7880
rect 25317 7871 25375 7877
rect 25317 7868 25329 7871
rect 25188 7840 25329 7868
rect 25188 7828 25194 7840
rect 25317 7837 25329 7840
rect 25363 7837 25375 7871
rect 25317 7831 25375 7837
rect 25866 7828 25872 7880
rect 25924 7868 25930 7880
rect 26344 7868 26372 7976
rect 28718 7896 28724 7948
rect 28776 7936 28782 7948
rect 28920 7936 28948 7976
rect 29638 7964 29644 8016
rect 29696 8004 29702 8016
rect 29696 7976 35894 8004
rect 29696 7964 29702 7976
rect 35866 7936 35894 7976
rect 37292 7936 37320 8035
rect 37734 8032 37740 8044
rect 37792 8032 37798 8084
rect 28776 7908 28856 7936
rect 28920 7908 32628 7936
rect 35866 7908 37320 7936
rect 28776 7896 28782 7908
rect 28442 7868 28448 7880
rect 25924 7840 26372 7868
rect 28403 7840 28448 7868
rect 25924 7828 25930 7840
rect 28442 7828 28448 7840
rect 28500 7828 28506 7880
rect 28828 7877 28856 7908
rect 28813 7871 28871 7877
rect 28813 7837 28825 7871
rect 28859 7837 28871 7871
rect 31386 7868 31392 7880
rect 28813 7831 28871 7837
rect 28966 7840 31392 7868
rect 15654 7809 15660 7812
rect 12406 7772 15608 7800
rect 10229 7763 10287 7769
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 9548 7704 9689 7732
rect 9548 7692 9554 7704
rect 9677 7701 9689 7704
rect 9723 7701 9735 7735
rect 9677 7695 9735 7701
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 12710 7732 12716 7744
rect 10928 7704 12716 7732
rect 10928 7692 10934 7704
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 13541 7735 13599 7741
rect 13541 7701 13553 7735
rect 13587 7732 13599 7735
rect 13722 7732 13728 7744
rect 13587 7704 13728 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 14645 7735 14703 7741
rect 14645 7701 14657 7735
rect 14691 7732 14703 7735
rect 14734 7732 14740 7744
rect 14691 7704 14740 7732
rect 14691 7701 14703 7704
rect 14645 7695 14703 7701
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 15580 7732 15608 7772
rect 15648 7763 15660 7809
rect 15712 7800 15718 7812
rect 17221 7803 17279 7809
rect 17221 7800 17233 7803
rect 15712 7772 15748 7800
rect 16592 7772 17233 7800
rect 15654 7760 15660 7763
rect 15712 7760 15718 7772
rect 16592 7732 16620 7772
rect 17221 7769 17233 7772
rect 17267 7800 17279 7803
rect 17773 7803 17831 7809
rect 17773 7800 17785 7803
rect 17267 7772 17785 7800
rect 17267 7769 17279 7772
rect 17221 7763 17279 7769
rect 17773 7769 17785 7772
rect 17819 7800 17831 7803
rect 17954 7800 17960 7812
rect 17819 7772 17960 7800
rect 17819 7769 17831 7772
rect 17773 7763 17831 7769
rect 17954 7760 17960 7772
rect 18012 7760 18018 7812
rect 18509 7803 18567 7809
rect 18509 7769 18521 7803
rect 18555 7800 18567 7803
rect 18598 7800 18604 7812
rect 18555 7772 18604 7800
rect 18555 7769 18567 7772
rect 18509 7763 18567 7769
rect 18598 7760 18604 7772
rect 18656 7760 18662 7812
rect 18693 7803 18751 7809
rect 18693 7769 18705 7803
rect 18739 7769 18751 7803
rect 18693 7763 18751 7769
rect 19337 7803 19395 7809
rect 19337 7769 19349 7803
rect 19383 7800 19395 7803
rect 20530 7800 20536 7812
rect 19383 7772 20536 7800
rect 19383 7769 19395 7772
rect 19337 7763 19395 7769
rect 16758 7732 16764 7744
rect 15580 7704 16620 7732
rect 16719 7704 16764 7732
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 18708 7732 18736 7763
rect 20530 7760 20536 7772
rect 20588 7760 20594 7812
rect 24581 7803 24639 7809
rect 24581 7769 24593 7803
rect 24627 7769 24639 7803
rect 24581 7763 24639 7769
rect 19426 7732 19432 7744
rect 18708 7704 19432 7732
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 20346 7732 20352 7744
rect 20307 7704 20352 7732
rect 20346 7692 20352 7704
rect 20404 7692 20410 7744
rect 21634 7732 21640 7744
rect 21595 7704 21640 7732
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 22465 7735 22523 7741
rect 22465 7701 22477 7735
rect 22511 7732 22523 7735
rect 22738 7732 22744 7744
rect 22511 7704 22744 7732
rect 22511 7701 22523 7704
rect 22465 7695 22523 7701
rect 22738 7692 22744 7704
rect 22796 7732 22802 7744
rect 24596 7732 24624 7763
rect 24670 7760 24676 7812
rect 24728 7800 24734 7812
rect 25590 7809 25596 7812
rect 24765 7803 24823 7809
rect 24765 7800 24777 7803
rect 24728 7772 24777 7800
rect 24728 7760 24734 7772
rect 24765 7769 24777 7772
rect 24811 7769 24823 7803
rect 24765 7763 24823 7769
rect 25584 7763 25596 7809
rect 25648 7800 25654 7812
rect 25648 7772 25684 7800
rect 25590 7760 25596 7763
rect 25648 7760 25654 7772
rect 28166 7760 28172 7812
rect 28224 7800 28230 7812
rect 28629 7803 28687 7809
rect 28629 7800 28641 7803
rect 28224 7772 28641 7800
rect 28224 7760 28230 7772
rect 28629 7769 28641 7772
rect 28675 7769 28687 7803
rect 28629 7763 28687 7769
rect 28721 7803 28779 7809
rect 28721 7769 28733 7803
rect 28767 7800 28779 7803
rect 28966 7800 28994 7840
rect 31386 7828 31392 7840
rect 31444 7828 31450 7880
rect 28767 7772 28994 7800
rect 31205 7803 31263 7809
rect 28767 7769 28779 7772
rect 28721 7763 28779 7769
rect 31205 7769 31217 7803
rect 31251 7769 31263 7803
rect 32600 7800 32628 7908
rect 34790 7828 34796 7880
rect 34848 7868 34854 7880
rect 35250 7868 35256 7880
rect 34848 7840 35256 7868
rect 34848 7828 34854 7840
rect 35250 7828 35256 7840
rect 35308 7828 35314 7880
rect 35621 7871 35679 7877
rect 35621 7837 35633 7871
rect 35667 7868 35679 7871
rect 36262 7868 36268 7880
rect 35667 7840 36268 7868
rect 35667 7837 35679 7840
rect 35621 7831 35679 7837
rect 36262 7828 36268 7840
rect 36320 7828 36326 7880
rect 58158 7868 58164 7880
rect 58119 7840 58164 7868
rect 58158 7828 58164 7840
rect 58216 7828 58222 7880
rect 35345 7803 35403 7809
rect 32600 7772 35112 7800
rect 31205 7763 31263 7769
rect 22796 7704 24624 7732
rect 22796 7692 22802 7704
rect 30282 7692 30288 7744
rect 30340 7732 30346 7744
rect 31220 7732 31248 7763
rect 35084 7741 35112 7772
rect 35345 7769 35357 7803
rect 35391 7769 35403 7803
rect 35345 7763 35403 7769
rect 30340 7704 31248 7732
rect 35069 7735 35127 7741
rect 30340 7692 30346 7704
rect 35069 7701 35081 7735
rect 35115 7701 35127 7735
rect 35360 7732 35388 7763
rect 35434 7760 35440 7812
rect 35492 7800 35498 7812
rect 35492 7772 35537 7800
rect 35492 7760 35498 7772
rect 37090 7732 37096 7744
rect 35360 7704 37096 7732
rect 35069 7695 35127 7701
rect 37090 7692 37096 7704
rect 37148 7692 37154 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 6178 7488 6184 7540
rect 6236 7528 6242 7540
rect 6546 7528 6552 7540
rect 6236 7500 6552 7528
rect 6236 7488 6242 7500
rect 6546 7488 6552 7500
rect 6604 7528 6610 7540
rect 10413 7531 10471 7537
rect 6604 7500 7972 7528
rect 6604 7488 6610 7500
rect 3418 7420 3424 7472
rect 3476 7460 3482 7472
rect 7374 7460 7380 7472
rect 3476 7432 6592 7460
rect 3476 7420 3482 7432
rect 3694 7392 3700 7404
rect 3655 7364 3700 7392
rect 3694 7352 3700 7364
rect 3752 7352 3758 7404
rect 3970 7392 3976 7404
rect 3931 7364 3976 7392
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 4120 7364 4165 7392
rect 4120 7352 4126 7364
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 5261 7395 5319 7401
rect 4304 7364 4349 7392
rect 4304 7352 4310 7364
rect 5261 7361 5273 7395
rect 5307 7392 5319 7395
rect 6362 7392 6368 7404
rect 5307 7364 6368 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 6564 7401 6592 7432
rect 6748 7432 7380 7460
rect 6748 7401 6776 7432
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 7558 7460 7564 7472
rect 7519 7432 7564 7460
rect 7558 7420 7564 7432
rect 7616 7420 7622 7472
rect 7944 7460 7972 7500
rect 10413 7497 10425 7531
rect 10459 7528 10471 7531
rect 12526 7528 12532 7540
rect 10459 7500 12532 7528
rect 10459 7497 10471 7500
rect 10413 7491 10471 7497
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 15565 7531 15623 7537
rect 15028 7500 15516 7528
rect 7944 7432 8064 7460
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 6914 7392 6920 7404
rect 6875 7364 6920 7392
rect 6733 7355 6791 7361
rect 6914 7352 6920 7364
rect 6972 7352 6978 7404
rect 7098 7392 7104 7404
rect 7059 7364 7104 7392
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7926 7392 7932 7404
rect 7887 7364 7932 7392
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 8036 7401 8064 7432
rect 11882 7420 11888 7472
rect 11940 7460 11946 7472
rect 12314 7463 12372 7469
rect 12314 7460 12326 7463
rect 11940 7432 12326 7460
rect 11940 7420 11946 7432
rect 12314 7429 12326 7432
rect 12360 7429 12372 7463
rect 12314 7423 12372 7429
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 12066 7392 12072 7404
rect 12027 7364 12072 7392
rect 8021 7355 8079 7361
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 12176 7364 14136 7392
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7324 3939 7327
rect 5350 7324 5356 7336
rect 3927 7296 5356 7324
rect 3927 7293 3939 7296
rect 3881 7287 3939 7293
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 6822 7324 6828 7336
rect 5960 7296 6684 7324
rect 6783 7296 6828 7324
rect 5960 7284 5966 7296
rect 6656 7268 6684 7296
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 12176 7324 12204 7364
rect 6932 7296 12204 7324
rect 1949 7259 2007 7265
rect 1949 7225 1961 7259
rect 1995 7256 2007 7259
rect 3053 7259 3111 7265
rect 1995 7228 2774 7256
rect 1995 7225 2007 7228
rect 1949 7219 2007 7225
rect 2501 7191 2559 7197
rect 2501 7157 2513 7191
rect 2547 7188 2559 7191
rect 2590 7188 2596 7200
rect 2547 7160 2596 7188
rect 2547 7157 2559 7160
rect 2501 7151 2559 7157
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 2746 7188 2774 7228
rect 3053 7225 3065 7259
rect 3099 7256 3111 7259
rect 4890 7256 4896 7268
rect 3099 7228 4896 7256
rect 3099 7225 3111 7228
rect 3053 7219 3111 7225
rect 4890 7216 4896 7228
rect 4948 7216 4954 7268
rect 5258 7216 5264 7268
rect 5316 7256 5322 7268
rect 6365 7259 6423 7265
rect 6365 7256 6377 7259
rect 5316 7228 6377 7256
rect 5316 7216 5322 7228
rect 6365 7225 6377 7228
rect 6411 7225 6423 7259
rect 6365 7219 6423 7225
rect 6638 7216 6644 7268
rect 6696 7256 6702 7268
rect 6932 7256 6960 7296
rect 6696 7228 6960 7256
rect 8205 7259 8263 7265
rect 6696 7216 6702 7228
rect 8205 7225 8217 7259
rect 8251 7256 8263 7259
rect 10042 7256 10048 7268
rect 8251 7228 10048 7256
rect 8251 7225 8263 7228
rect 8205 7219 8263 7225
rect 10042 7216 10048 7228
rect 10100 7216 10106 7268
rect 10965 7259 11023 7265
rect 10965 7225 10977 7259
rect 11011 7256 11023 7259
rect 14108 7256 14136 7364
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 14918 7392 14924 7404
rect 14240 7364 14285 7392
rect 14879 7364 14924 7392
rect 14240 7352 14246 7364
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15028 7392 15056 7500
rect 15488 7460 15516 7500
rect 15565 7497 15577 7531
rect 15611 7528 15623 7531
rect 15654 7528 15660 7540
rect 15611 7500 15660 7528
rect 15611 7497 15623 7500
rect 15565 7491 15623 7497
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 17586 7488 17592 7540
rect 17644 7528 17650 7540
rect 18138 7528 18144 7540
rect 17644 7500 18144 7528
rect 17644 7488 17650 7500
rect 18138 7488 18144 7500
rect 18196 7488 18202 7540
rect 18506 7488 18512 7540
rect 18564 7528 18570 7540
rect 23017 7531 23075 7537
rect 18564 7500 22968 7528
rect 18564 7488 18570 7500
rect 16669 7463 16727 7469
rect 16669 7460 16681 7463
rect 15488 7432 16681 7460
rect 16669 7429 16681 7432
rect 16715 7429 16727 7463
rect 16669 7423 16727 7429
rect 16758 7420 16764 7472
rect 16816 7460 16822 7472
rect 16853 7463 16911 7469
rect 16853 7460 16865 7463
rect 16816 7432 16865 7460
rect 16816 7420 16822 7432
rect 16853 7429 16865 7432
rect 16899 7460 16911 7463
rect 22186 7460 22192 7472
rect 16899 7432 21036 7460
rect 16899 7429 16911 7432
rect 16853 7423 16911 7429
rect 15084 7395 15142 7401
rect 15084 7392 15096 7395
rect 15028 7364 15096 7392
rect 15084 7361 15096 7364
rect 15130 7361 15142 7395
rect 15084 7355 15142 7361
rect 15200 7395 15258 7401
rect 15200 7361 15212 7395
rect 15246 7361 15258 7395
rect 15309 7395 15367 7401
rect 15309 7392 15321 7395
rect 15200 7355 15258 7361
rect 15304 7361 15321 7392
rect 15355 7361 15367 7395
rect 17034 7392 17040 7404
rect 16947 7364 17040 7392
rect 15304 7355 15367 7361
rect 14550 7284 14556 7336
rect 14608 7324 14614 7336
rect 15215 7324 15243 7355
rect 14608 7296 15243 7324
rect 14608 7284 14614 7296
rect 15304 7256 15332 7355
rect 17034 7352 17040 7364
rect 17092 7392 17098 7404
rect 17865 7395 17923 7401
rect 17092 7364 17816 7392
rect 17092 7352 17098 7364
rect 15930 7256 15936 7268
rect 11011 7228 11652 7256
rect 14108 7228 15936 7256
rect 11011 7225 11023 7228
rect 10965 7219 11023 7225
rect 3142 7188 3148 7200
rect 2746 7160 3148 7188
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3510 7188 3516 7200
rect 3471 7160 3516 7188
rect 3510 7148 3516 7160
rect 3568 7148 3574 7200
rect 3970 7148 3976 7200
rect 4028 7188 4034 7200
rect 4246 7188 4252 7200
rect 4028 7160 4252 7188
rect 4028 7148 4034 7160
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 5813 7191 5871 7197
rect 5813 7157 5825 7191
rect 5859 7188 5871 7191
rect 7742 7188 7748 7200
rect 5859 7160 7748 7188
rect 5859 7157 5871 7160
rect 5813 7151 5871 7157
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 8757 7191 8815 7197
rect 8757 7188 8769 7191
rect 8628 7160 8769 7188
rect 8628 7148 8634 7160
rect 8757 7157 8769 7160
rect 8803 7157 8815 7191
rect 8757 7151 8815 7157
rect 9861 7191 9919 7197
rect 9861 7157 9873 7191
rect 9907 7188 9919 7191
rect 10318 7188 10324 7200
rect 9907 7160 10324 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 10928 7160 11529 7188
rect 10928 7148 10934 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 11624 7188 11652 7228
rect 15930 7216 15936 7228
rect 15988 7256 15994 7268
rect 16025 7259 16083 7265
rect 16025 7256 16037 7259
rect 15988 7228 16037 7256
rect 15988 7216 15994 7228
rect 16025 7225 16037 7228
rect 16071 7225 16083 7259
rect 16025 7219 16083 7225
rect 13170 7188 13176 7200
rect 11624 7160 13176 7188
rect 11517 7151 11575 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13446 7188 13452 7200
rect 13407 7160 13452 7188
rect 13446 7148 13452 7160
rect 13504 7148 13510 7200
rect 14090 7188 14096 7200
rect 14051 7160 14096 7188
rect 14090 7148 14096 7160
rect 14148 7148 14154 7200
rect 17788 7188 17816 7364
rect 17865 7361 17877 7395
rect 17911 7392 17923 7395
rect 19337 7395 19395 7401
rect 17911 7364 18460 7392
rect 17911 7361 17923 7364
rect 17865 7355 17923 7361
rect 18138 7324 18144 7336
rect 18099 7296 18144 7324
rect 18138 7284 18144 7296
rect 18196 7284 18202 7336
rect 18432 7324 18460 7364
rect 19337 7361 19349 7395
rect 19383 7392 19395 7395
rect 19426 7392 19432 7404
rect 19383 7364 19432 7392
rect 19383 7361 19395 7364
rect 19337 7355 19395 7361
rect 19426 7352 19432 7364
rect 19484 7352 19490 7404
rect 20162 7352 20168 7404
rect 20220 7392 20226 7404
rect 20438 7392 20444 7404
rect 20220 7364 20444 7392
rect 20220 7352 20226 7364
rect 20438 7352 20444 7364
rect 20496 7392 20502 7404
rect 20901 7395 20959 7401
rect 20901 7392 20913 7395
rect 20496 7364 20913 7392
rect 20496 7352 20502 7364
rect 20901 7361 20913 7364
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 18874 7324 18880 7336
rect 18432 7296 18880 7324
rect 18874 7284 18880 7296
rect 18932 7324 18938 7336
rect 21008 7324 21036 7432
rect 21100 7432 22192 7460
rect 21100 7401 21128 7432
rect 21085 7395 21143 7401
rect 21085 7361 21097 7395
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 21174 7352 21180 7404
rect 21232 7392 21238 7404
rect 21634 7392 21640 7404
rect 21232 7364 21640 7392
rect 21232 7352 21238 7364
rect 21634 7352 21640 7364
rect 21692 7392 21698 7404
rect 22020 7401 22048 7432
rect 22186 7420 22192 7432
rect 22244 7460 22250 7472
rect 22738 7460 22744 7472
rect 22244 7432 22600 7460
rect 22699 7432 22744 7460
rect 22244 7420 22250 7432
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 21692 7364 21833 7392
rect 21692 7352 21698 7364
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22465 7395 22523 7401
rect 22465 7361 22477 7395
rect 22511 7361 22523 7395
rect 22572 7392 22600 7432
rect 22738 7420 22744 7432
rect 22796 7420 22802 7472
rect 22940 7460 22968 7500
rect 23017 7497 23029 7531
rect 23063 7528 23075 7531
rect 24118 7528 24124 7540
rect 23063 7500 24124 7528
rect 23063 7497 23075 7500
rect 23017 7491 23075 7497
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 24670 7488 24676 7540
rect 24728 7528 24734 7540
rect 25590 7528 25596 7540
rect 24728 7500 25360 7528
rect 25551 7500 25596 7528
rect 24728 7488 24734 7500
rect 22940 7432 23796 7460
rect 22649 7395 22707 7401
rect 22649 7392 22661 7395
rect 22572 7364 22661 7392
rect 22465 7355 22523 7361
rect 22649 7361 22661 7364
rect 22695 7361 22707 7395
rect 22830 7392 22836 7404
rect 22791 7364 22836 7392
rect 22649 7355 22707 7361
rect 22480 7324 22508 7355
rect 22830 7352 22836 7364
rect 22888 7352 22894 7404
rect 22922 7352 22928 7404
rect 22980 7392 22986 7404
rect 23661 7395 23719 7401
rect 23661 7392 23673 7395
rect 22980 7364 23673 7392
rect 22980 7352 22986 7364
rect 23661 7361 23673 7364
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 18932 7296 20944 7324
rect 21008 7296 22508 7324
rect 23768 7324 23796 7432
rect 24210 7420 24216 7472
rect 24268 7460 24274 7472
rect 25332 7460 25360 7500
rect 25590 7488 25596 7500
rect 25648 7488 25654 7540
rect 28350 7488 28356 7540
rect 28408 7528 28414 7540
rect 28629 7531 28687 7537
rect 28629 7528 28641 7531
rect 28408 7500 28641 7528
rect 28408 7488 28414 7500
rect 28629 7497 28641 7500
rect 28675 7497 28687 7531
rect 28629 7491 28687 7497
rect 31386 7488 31392 7540
rect 31444 7528 31450 7540
rect 32493 7531 32551 7537
rect 32493 7528 32505 7531
rect 31444 7500 32505 7528
rect 31444 7488 31450 7500
rect 32493 7497 32505 7500
rect 32539 7497 32551 7531
rect 32493 7491 32551 7497
rect 34514 7488 34520 7540
rect 34572 7528 34578 7540
rect 35069 7531 35127 7537
rect 35069 7528 35081 7531
rect 34572 7500 35081 7528
rect 34572 7488 34578 7500
rect 35069 7497 35081 7500
rect 35115 7497 35127 7531
rect 35069 7491 35127 7497
rect 36357 7531 36415 7537
rect 36357 7497 36369 7531
rect 36403 7528 36415 7531
rect 38102 7528 38108 7540
rect 36403 7500 38108 7528
rect 36403 7497 36415 7500
rect 36357 7491 36415 7497
rect 38102 7488 38108 7500
rect 38160 7488 38166 7540
rect 26053 7463 26111 7469
rect 26053 7460 26065 7463
rect 24268 7432 25268 7460
rect 25332 7432 26065 7460
rect 24268 7420 24274 7432
rect 23845 7395 23903 7401
rect 23845 7361 23857 7395
rect 23891 7392 23903 7395
rect 24394 7392 24400 7404
rect 23891 7364 24400 7392
rect 23891 7361 23903 7364
rect 23845 7355 23903 7361
rect 24394 7352 24400 7364
rect 24452 7352 24458 7404
rect 24578 7352 24584 7404
rect 24636 7392 24642 7404
rect 25240 7401 25268 7432
rect 26053 7429 26065 7432
rect 26099 7429 26111 7463
rect 26234 7460 26240 7472
rect 26195 7432 26240 7460
rect 26053 7423 26111 7429
rect 26234 7420 26240 7432
rect 26292 7420 26298 7472
rect 29638 7460 29644 7472
rect 26344 7432 29644 7460
rect 24949 7395 25007 7401
rect 24949 7392 24961 7395
rect 24636 7364 24961 7392
rect 24636 7352 24642 7364
rect 24949 7361 24961 7364
rect 24995 7361 25007 7395
rect 24949 7355 25007 7361
rect 25133 7395 25191 7401
rect 25133 7361 25145 7395
rect 25179 7361 25191 7395
rect 25133 7355 25191 7361
rect 25225 7395 25283 7401
rect 25225 7361 25237 7395
rect 25271 7361 25283 7395
rect 25225 7355 25283 7361
rect 24412 7324 24440 7352
rect 24670 7324 24676 7336
rect 23768 7296 24348 7324
rect 24412 7296 24676 7324
rect 18932 7284 18938 7296
rect 19889 7259 19947 7265
rect 19889 7225 19901 7259
rect 19935 7256 19947 7259
rect 20438 7256 20444 7268
rect 19935 7228 20444 7256
rect 19935 7225 19947 7228
rect 19889 7219 19947 7225
rect 20438 7216 20444 7228
rect 20496 7216 20502 7268
rect 20916 7256 20944 7296
rect 24320 7256 24348 7296
rect 24670 7284 24676 7296
rect 24728 7284 24734 7336
rect 25148 7324 25176 7355
rect 25314 7352 25320 7404
rect 25372 7392 25378 7404
rect 26344 7392 26372 7432
rect 29638 7420 29644 7432
rect 29696 7420 29702 7472
rect 30377 7463 30435 7469
rect 30377 7429 30389 7463
rect 30423 7460 30435 7463
rect 31294 7460 31300 7472
rect 30423 7432 31300 7460
rect 30423 7429 30435 7432
rect 30377 7423 30435 7429
rect 31294 7420 31300 7432
rect 31352 7420 31358 7472
rect 33594 7420 33600 7472
rect 33652 7469 33658 7472
rect 33652 7460 33664 7469
rect 35434 7460 35440 7472
rect 33652 7432 33697 7460
rect 35395 7432 35440 7460
rect 33652 7423 33664 7432
rect 33652 7420 33658 7423
rect 35434 7420 35440 7432
rect 35492 7420 35498 7472
rect 37642 7420 37648 7472
rect 37700 7460 37706 7472
rect 38657 7463 38715 7469
rect 38657 7460 38669 7463
rect 37700 7432 38669 7460
rect 37700 7420 37706 7432
rect 38657 7429 38669 7432
rect 38703 7429 38715 7463
rect 38657 7423 38715 7429
rect 25372 7364 26372 7392
rect 25372 7352 25378 7364
rect 27338 7352 27344 7404
rect 27396 7392 27402 7404
rect 27505 7395 27563 7401
rect 27505 7392 27517 7395
rect 27396 7364 27517 7392
rect 27396 7352 27402 7364
rect 27505 7361 27517 7364
rect 27551 7361 27563 7395
rect 27505 7355 27563 7361
rect 30561 7395 30619 7401
rect 30561 7361 30573 7395
rect 30607 7392 30619 7395
rect 31110 7392 31116 7404
rect 30607 7364 31116 7392
rect 30607 7361 30619 7364
rect 30561 7355 30619 7361
rect 31110 7352 31116 7364
rect 31168 7352 31174 7404
rect 35250 7392 35256 7404
rect 35211 7364 35256 7392
rect 35250 7352 35256 7364
rect 35308 7352 35314 7404
rect 35345 7395 35403 7401
rect 35345 7361 35357 7395
rect 35391 7361 35403 7395
rect 35618 7392 35624 7404
rect 35579 7364 35624 7392
rect 35345 7355 35403 7361
rect 26421 7327 26479 7333
rect 26421 7324 26433 7327
rect 25148 7296 26433 7324
rect 26421 7293 26433 7296
rect 26467 7293 26479 7327
rect 27246 7324 27252 7336
rect 27207 7296 27252 7324
rect 26421 7287 26479 7293
rect 27246 7284 27252 7296
rect 27304 7284 27310 7336
rect 33873 7327 33931 7333
rect 33873 7293 33885 7327
rect 33919 7324 33931 7327
rect 34790 7324 34796 7336
rect 33919 7296 34796 7324
rect 33919 7293 33931 7296
rect 33873 7287 33931 7293
rect 34790 7284 34796 7296
rect 34848 7284 34854 7336
rect 35360 7324 35388 7355
rect 35618 7352 35624 7364
rect 35676 7352 35682 7404
rect 38841 7395 38899 7401
rect 38841 7361 38853 7395
rect 38887 7361 38899 7395
rect 38841 7355 38899 7361
rect 38856 7324 38884 7355
rect 39666 7324 39672 7336
rect 35360 7296 39672 7324
rect 39666 7284 39672 7296
rect 39724 7284 39730 7336
rect 24397 7259 24455 7265
rect 24397 7256 24409 7259
rect 20916 7228 21956 7256
rect 24320 7228 24409 7256
rect 21928 7200 21956 7228
rect 24397 7225 24409 7228
rect 24443 7256 24455 7259
rect 25314 7256 25320 7268
rect 24443 7228 25320 7256
rect 24443 7225 24455 7228
rect 24397 7219 24455 7225
rect 25314 7216 25320 7228
rect 25372 7216 25378 7268
rect 19153 7191 19211 7197
rect 19153 7188 19165 7191
rect 17788 7160 19165 7188
rect 19153 7157 19165 7160
rect 19199 7188 19211 7191
rect 19242 7188 19248 7200
rect 19199 7160 19248 7188
rect 19199 7157 19211 7160
rect 19153 7151 19211 7157
rect 19242 7148 19248 7160
rect 19300 7148 19306 7200
rect 20162 7148 20168 7200
rect 20220 7188 20226 7200
rect 20349 7191 20407 7197
rect 20349 7188 20361 7191
rect 20220 7160 20361 7188
rect 20220 7148 20226 7160
rect 20349 7157 20361 7160
rect 20395 7157 20407 7191
rect 21266 7188 21272 7200
rect 21227 7160 21272 7188
rect 20349 7151 20407 7157
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 21910 7188 21916 7200
rect 21871 7160 21916 7188
rect 21910 7148 21916 7160
rect 21968 7148 21974 7200
rect 23477 7191 23535 7197
rect 23477 7157 23489 7191
rect 23523 7188 23535 7191
rect 23658 7188 23664 7200
rect 23523 7160 23664 7188
rect 23523 7157 23535 7160
rect 23477 7151 23535 7157
rect 23658 7148 23664 7160
rect 23716 7148 23722 7200
rect 29638 7148 29644 7200
rect 29696 7188 29702 7200
rect 30193 7191 30251 7197
rect 30193 7188 30205 7191
rect 29696 7160 30205 7188
rect 29696 7148 29702 7160
rect 30193 7157 30205 7160
rect 30239 7157 30251 7191
rect 30193 7151 30251 7157
rect 38838 7148 38844 7200
rect 38896 7188 38902 7200
rect 39025 7191 39083 7197
rect 39025 7188 39037 7191
rect 38896 7160 39037 7188
rect 38896 7148 38902 7160
rect 39025 7157 39037 7160
rect 39071 7157 39083 7191
rect 39025 7151 39083 7157
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 4341 6987 4399 6993
rect 4341 6984 4353 6987
rect 4120 6956 4353 6984
rect 4120 6944 4126 6956
rect 4341 6953 4353 6956
rect 4387 6953 4399 6987
rect 4341 6947 4399 6953
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 21174 6984 21180 6996
rect 14148 6956 21180 6984
rect 14148 6944 14154 6956
rect 21174 6944 21180 6956
rect 21232 6944 21238 6996
rect 21266 6944 21272 6996
rect 21324 6984 21330 6996
rect 26970 6984 26976 6996
rect 21324 6956 26976 6984
rect 21324 6944 21330 6956
rect 26970 6944 26976 6956
rect 27028 6944 27034 6996
rect 30926 6984 30932 6996
rect 29932 6956 30932 6984
rect 9858 6916 9864 6928
rect 7852 6888 8800 6916
rect 9771 6888 9864 6916
rect 2685 6851 2743 6857
rect 2685 6817 2697 6851
rect 2731 6848 2743 6851
rect 2731 6820 3924 6848
rect 2731 6817 2743 6820
rect 2685 6811 2743 6817
rect 2133 6783 2191 6789
rect 2133 6749 2145 6783
rect 2179 6780 2191 6783
rect 3326 6780 3332 6792
rect 2179 6752 3332 6780
rect 2179 6749 2191 6752
rect 2133 6743 2191 6749
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3896 6780 3924 6820
rect 3970 6808 3976 6860
rect 4028 6848 4034 6860
rect 6733 6851 6791 6857
rect 6733 6848 6745 6851
rect 4028 6820 6745 6848
rect 4028 6808 4034 6820
rect 6733 6817 6745 6820
rect 6779 6848 6791 6851
rect 7852 6848 7880 6888
rect 8662 6848 8668 6860
rect 6779 6820 7880 6848
rect 7944 6820 8668 6848
rect 6779 6817 6791 6820
rect 6733 6811 6791 6817
rect 4522 6780 4528 6792
rect 3896 6752 4528 6780
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 4985 6783 5043 6789
rect 4985 6780 4997 6783
rect 4672 6752 4997 6780
rect 4672 6740 4678 6752
rect 4985 6749 4997 6752
rect 5031 6749 5043 6783
rect 4985 6743 5043 6749
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 6454 6780 6460 6792
rect 5123 6752 6460 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 6454 6740 6460 6752
rect 6512 6740 6518 6792
rect 7944 6789 7972 6820
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 8772 6848 8800 6888
rect 9858 6876 9864 6888
rect 9916 6916 9922 6928
rect 13265 6919 13323 6925
rect 9916 6888 10180 6916
rect 9916 6876 9922 6888
rect 9876 6848 9904 6876
rect 10042 6848 10048 6860
rect 8772 6820 9904 6848
rect 10003 6820 10048 6848
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 10152 6848 10180 6888
rect 13265 6885 13277 6919
rect 13311 6916 13323 6919
rect 13311 6888 19334 6916
rect 13311 6885 13323 6888
rect 13265 6879 13323 6885
rect 11517 6851 11575 6857
rect 10152 6820 10364 6848
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6749 7987 6783
rect 7929 6743 7987 6749
rect 8570 6740 8576 6792
rect 8628 6780 8634 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8628 6752 8953 6780
rect 8628 6740 8634 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6749 9827 6783
rect 9950 6780 9956 6792
rect 9911 6752 9956 6780
rect 9769 6743 9827 6749
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 3050 6712 3056 6724
rect 1627 6684 3056 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 3050 6672 3056 6684
rect 3108 6672 3114 6724
rect 9490 6712 9496 6724
rect 3804 6684 9496 6712
rect 3804 6656 3832 6684
rect 9490 6672 9496 6684
rect 9548 6672 9554 6724
rect 9784 6712 9812 6743
rect 9950 6740 9956 6752
rect 10008 6740 10014 6792
rect 10134 6740 10140 6792
rect 10192 6780 10198 6792
rect 10336 6789 10364 6820
rect 11517 6817 11529 6851
rect 11563 6848 11575 6851
rect 13354 6848 13360 6860
rect 11563 6820 13360 6848
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 13354 6808 13360 6820
rect 13412 6808 13418 6860
rect 15470 6848 15476 6860
rect 15383 6820 15476 6848
rect 15470 6808 15476 6820
rect 15528 6848 15534 6860
rect 19306 6848 19334 6888
rect 19426 6876 19432 6928
rect 19484 6916 19490 6928
rect 21284 6916 21312 6944
rect 19484 6888 21312 6916
rect 19484 6876 19490 6888
rect 23934 6876 23940 6928
rect 23992 6916 23998 6928
rect 24578 6916 24584 6928
rect 23992 6888 24584 6916
rect 23992 6876 23998 6888
rect 24578 6876 24584 6888
rect 24636 6916 24642 6928
rect 24636 6888 25084 6916
rect 24636 6876 24642 6888
rect 20162 6848 20168 6860
rect 15528 6820 16068 6848
rect 19306 6820 20168 6848
rect 15528 6808 15534 6820
rect 16040 6792 16068 6820
rect 20162 6808 20168 6820
rect 20220 6808 20226 6860
rect 21913 6851 21971 6857
rect 21913 6817 21925 6851
rect 21959 6848 21971 6851
rect 22646 6848 22652 6860
rect 21959 6820 22652 6848
rect 21959 6817 21971 6820
rect 21913 6811 21971 6817
rect 22646 6808 22652 6820
rect 22704 6808 22710 6860
rect 24397 6851 24455 6857
rect 23124 6820 24072 6848
rect 10321 6783 10379 6789
rect 10192 6752 10237 6780
rect 10192 6740 10198 6752
rect 10321 6749 10333 6783
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 10502 6740 10508 6792
rect 10560 6780 10566 6792
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 10560 6752 10793 6780
rect 10560 6740 10566 6752
rect 10781 6749 10793 6752
rect 10827 6749 10839 6783
rect 11974 6780 11980 6792
rect 11935 6752 11980 6780
rect 10781 6743 10839 6749
rect 11974 6740 11980 6752
rect 12032 6780 12038 6792
rect 12342 6780 12348 6792
rect 12032 6752 12348 6780
rect 12032 6740 12038 6752
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 12492 6752 12725 6780
rect 12492 6740 12498 6752
rect 12713 6749 12725 6752
rect 12759 6780 12771 6783
rect 13538 6780 13544 6792
rect 12759 6752 13544 6780
rect 12759 6749 12771 6752
rect 12713 6743 12771 6749
rect 13538 6740 13544 6752
rect 13596 6780 13602 6792
rect 14415 6783 14473 6789
rect 14415 6780 14427 6783
rect 13596 6752 14427 6780
rect 13596 6740 13602 6752
rect 14415 6749 14427 6752
rect 14461 6749 14473 6783
rect 14550 6780 14556 6792
rect 14511 6752 14556 6780
rect 14415 6743 14473 6749
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 14642 6740 14648 6792
rect 14700 6789 14706 6792
rect 14700 6780 14708 6789
rect 14829 6783 14887 6789
rect 14700 6752 14745 6780
rect 14700 6743 14708 6752
rect 14829 6749 14841 6783
rect 14875 6780 14887 6783
rect 14918 6780 14924 6792
rect 14875 6752 14924 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 14700 6740 14706 6743
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 16022 6740 16028 6792
rect 16080 6780 16086 6792
rect 16301 6783 16359 6789
rect 16080 6752 16125 6780
rect 16080 6740 16086 6752
rect 16301 6749 16313 6783
rect 16347 6780 16359 6783
rect 17770 6780 17776 6792
rect 16347 6752 17776 6780
rect 16347 6749 16359 6752
rect 16301 6743 16359 6749
rect 11054 6712 11060 6724
rect 9784 6684 11060 6712
rect 11054 6672 11060 6684
rect 11112 6672 11118 6724
rect 12406 6684 12848 6712
rect 3234 6644 3240 6656
rect 3195 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3786 6644 3792 6656
rect 3747 6616 3792 6644
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 5166 6644 5172 6656
rect 4580 6616 5172 6644
rect 4580 6604 4586 6616
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 5997 6647 6055 6653
rect 5997 6613 6009 6647
rect 6043 6644 6055 6647
rect 7006 6644 7012 6656
rect 6043 6616 7012 6644
rect 6043 6613 6055 6616
rect 5997 6607 6055 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 8113 6647 8171 6653
rect 8113 6613 8125 6647
rect 8159 6644 8171 6647
rect 8202 6644 8208 6656
rect 8159 6616 8208 6644
rect 8159 6613 8171 6616
rect 8113 6607 8171 6613
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8478 6604 8484 6656
rect 8536 6644 8542 6656
rect 9122 6644 9128 6656
rect 8536 6616 9128 6644
rect 8536 6604 8542 6616
rect 9122 6604 9128 6616
rect 9180 6604 9186 6656
rect 9585 6647 9643 6653
rect 9585 6613 9597 6647
rect 9631 6644 9643 6647
rect 9858 6644 9864 6656
rect 9631 6616 9864 6644
rect 9631 6613 9643 6616
rect 9585 6607 9643 6613
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 12161 6647 12219 6653
rect 12161 6613 12173 6647
rect 12207 6644 12219 6647
rect 12406 6644 12434 6684
rect 12207 6616 12434 6644
rect 12820 6644 12848 6684
rect 12894 6672 12900 6724
rect 12952 6712 12958 6724
rect 13449 6715 13507 6721
rect 13449 6712 13461 6715
rect 12952 6684 13461 6712
rect 12952 6672 12958 6684
rect 13449 6681 13461 6684
rect 13495 6712 13507 6715
rect 14090 6712 14096 6724
rect 13495 6684 14096 6712
rect 13495 6681 13507 6684
rect 13449 6675 13507 6681
rect 14090 6672 14096 6684
rect 14148 6672 14154 6724
rect 13906 6644 13912 6656
rect 12820 6616 13912 6644
rect 12207 6613 12219 6616
rect 12161 6607 12219 6613
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 13998 6604 14004 6656
rect 14056 6644 14062 6656
rect 14185 6647 14243 6653
rect 14185 6644 14197 6647
rect 14056 6616 14197 6644
rect 14056 6604 14062 6616
rect 14185 6613 14197 6616
rect 14231 6613 14243 6647
rect 14185 6607 14243 6613
rect 14918 6604 14924 6656
rect 14976 6644 14982 6656
rect 16316 6644 16344 6743
rect 17770 6740 17776 6752
rect 17828 6740 17834 6792
rect 18230 6740 18236 6792
rect 18288 6780 18294 6792
rect 21634 6780 21640 6792
rect 18288 6752 20300 6780
rect 21595 6752 21640 6780
rect 18288 6740 18294 6752
rect 19337 6715 19395 6721
rect 19337 6681 19349 6715
rect 19383 6712 19395 6715
rect 20162 6712 20168 6724
rect 19383 6684 20168 6712
rect 19383 6681 19395 6684
rect 19337 6675 19395 6681
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 20272 6712 20300 6752
rect 21634 6740 21640 6752
rect 21692 6740 21698 6792
rect 23124 6712 23152 6820
rect 23382 6740 23388 6792
rect 23440 6780 23446 6792
rect 23477 6783 23535 6789
rect 23477 6780 23489 6783
rect 23440 6752 23489 6780
rect 23440 6740 23446 6752
rect 23477 6749 23489 6752
rect 23523 6749 23535 6783
rect 23477 6743 23535 6749
rect 23569 6783 23627 6789
rect 23569 6749 23581 6783
rect 23615 6749 23627 6783
rect 23569 6743 23627 6749
rect 20272 6684 23152 6712
rect 23584 6712 23612 6743
rect 23658 6740 23664 6792
rect 23716 6780 23722 6792
rect 23845 6783 23903 6789
rect 23716 6752 23761 6780
rect 23716 6740 23722 6752
rect 23845 6749 23857 6783
rect 23891 6780 23903 6783
rect 23934 6780 23940 6792
rect 23891 6752 23940 6780
rect 23891 6749 23903 6752
rect 23845 6743 23903 6749
rect 23934 6740 23940 6752
rect 23992 6740 23998 6792
rect 24044 6780 24072 6820
rect 24397 6817 24409 6851
rect 24443 6848 24455 6851
rect 24946 6848 24952 6860
rect 24443 6820 24952 6848
rect 24443 6817 24455 6820
rect 24397 6811 24455 6817
rect 24946 6808 24952 6820
rect 25004 6808 25010 6860
rect 24578 6780 24584 6792
rect 24044 6752 24584 6780
rect 24578 6740 24584 6752
rect 24636 6780 24642 6792
rect 25056 6789 25084 6888
rect 27246 6876 27252 6928
rect 27304 6916 27310 6928
rect 29932 6916 29960 6956
rect 30926 6944 30932 6956
rect 30984 6944 30990 6996
rect 31294 6984 31300 6996
rect 31255 6956 31300 6984
rect 31294 6944 31300 6956
rect 31352 6944 31358 6996
rect 35989 6987 36047 6993
rect 35989 6984 36001 6987
rect 35176 6956 36001 6984
rect 27304 6888 29960 6916
rect 27304 6876 27310 6888
rect 25958 6848 25964 6860
rect 25919 6820 25964 6848
rect 25958 6808 25964 6820
rect 26016 6808 26022 6860
rect 26237 6851 26295 6857
rect 26237 6817 26249 6851
rect 26283 6848 26295 6851
rect 27062 6848 27068 6860
rect 26283 6820 27068 6848
rect 26283 6817 26295 6820
rect 26237 6811 26295 6817
rect 27062 6808 27068 6820
rect 27120 6848 27126 6860
rect 29932 6857 29960 6888
rect 28353 6851 28411 6857
rect 28353 6848 28365 6851
rect 27120 6820 27660 6848
rect 27120 6808 27126 6820
rect 24673 6783 24731 6789
rect 24673 6780 24685 6783
rect 24636 6752 24685 6780
rect 24636 6740 24642 6752
rect 24673 6749 24685 6752
rect 24719 6749 24731 6783
rect 24673 6743 24731 6749
rect 24765 6783 24823 6789
rect 24765 6749 24777 6783
rect 24811 6749 24823 6783
rect 24765 6743 24823 6749
rect 24857 6783 24915 6789
rect 24857 6749 24869 6783
rect 24903 6749 24915 6783
rect 24857 6743 24915 6749
rect 25041 6783 25099 6789
rect 25041 6749 25053 6783
rect 25087 6749 25099 6783
rect 27522 6780 27528 6792
rect 27483 6752 27528 6780
rect 25041 6743 25099 6749
rect 24210 6712 24216 6724
rect 23584 6684 24216 6712
rect 24210 6672 24216 6684
rect 24268 6712 24274 6724
rect 24780 6712 24808 6743
rect 24268 6684 24808 6712
rect 24268 6672 24274 6684
rect 17586 6644 17592 6656
rect 14976 6616 16344 6644
rect 17547 6616 17592 6644
rect 14976 6604 14982 6616
rect 17586 6604 17592 6616
rect 17644 6604 17650 6656
rect 18322 6644 18328 6656
rect 18283 6616 18328 6644
rect 18322 6604 18328 6616
rect 18380 6604 18386 6656
rect 19978 6644 19984 6656
rect 19939 6616 19984 6644
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 20714 6644 20720 6656
rect 20675 6616 20720 6644
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 23201 6647 23259 6653
rect 23201 6613 23213 6647
rect 23247 6644 23259 6647
rect 23566 6644 23572 6656
rect 23247 6616 23572 6644
rect 23247 6613 23259 6616
rect 23201 6607 23259 6613
rect 23566 6604 23572 6616
rect 23624 6604 23630 6656
rect 24762 6604 24768 6656
rect 24820 6644 24826 6656
rect 24872 6644 24900 6743
rect 27522 6740 27528 6752
rect 27580 6740 27586 6792
rect 27632 6789 27660 6820
rect 27724 6820 28365 6848
rect 27724 6789 27752 6820
rect 28353 6817 28365 6820
rect 28399 6817 28411 6851
rect 28353 6811 28411 6817
rect 29917 6851 29975 6857
rect 29917 6817 29929 6851
rect 29963 6817 29975 6851
rect 35176 6848 35204 6956
rect 35989 6953 36001 6956
rect 36035 6984 36047 6987
rect 38562 6984 38568 6996
rect 36035 6956 38568 6984
rect 36035 6953 36047 6956
rect 35989 6947 36047 6953
rect 38562 6944 38568 6956
rect 38620 6944 38626 6996
rect 38746 6944 38752 6996
rect 38804 6984 38810 6996
rect 39853 6987 39911 6993
rect 39853 6984 39865 6987
rect 38804 6956 39865 6984
rect 38804 6944 38810 6956
rect 39853 6953 39865 6956
rect 39899 6953 39911 6987
rect 39853 6947 39911 6953
rect 35802 6916 35808 6928
rect 29917 6811 29975 6817
rect 33704 6820 35204 6848
rect 27617 6783 27675 6789
rect 27617 6749 27629 6783
rect 27663 6749 27675 6783
rect 27617 6743 27675 6749
rect 27709 6783 27767 6789
rect 27709 6749 27721 6783
rect 27755 6749 27767 6783
rect 27709 6743 27767 6749
rect 27893 6783 27951 6789
rect 27893 6749 27905 6783
rect 27939 6749 27951 6783
rect 27893 6743 27951 6749
rect 27249 6715 27307 6721
rect 27249 6681 27261 6715
rect 27295 6712 27307 6715
rect 27338 6712 27344 6724
rect 27295 6684 27344 6712
rect 27295 6681 27307 6684
rect 27249 6675 27307 6681
rect 27338 6672 27344 6684
rect 27396 6672 27402 6724
rect 27908 6712 27936 6743
rect 28166 6740 28172 6792
rect 28224 6780 28230 6792
rect 28721 6783 28779 6789
rect 28721 6780 28733 6783
rect 28224 6752 28733 6780
rect 28224 6740 28230 6752
rect 28721 6749 28733 6752
rect 28767 6780 28779 6783
rect 31110 6780 31116 6792
rect 28767 6752 31116 6780
rect 28767 6749 28779 6752
rect 28721 6743 28779 6749
rect 31110 6740 31116 6752
rect 31168 6740 31174 6792
rect 27540 6684 27936 6712
rect 27540 6656 27568 6684
rect 28350 6672 28356 6724
rect 28408 6712 28414 6724
rect 30190 6721 30196 6724
rect 28537 6715 28595 6721
rect 28537 6712 28549 6715
rect 28408 6684 28549 6712
rect 28408 6672 28414 6684
rect 28537 6681 28549 6684
rect 28583 6681 28595 6715
rect 28537 6675 28595 6681
rect 30184 6675 30196 6721
rect 30248 6712 30254 6724
rect 30248 6684 30284 6712
rect 30190 6672 30196 6675
rect 30248 6672 30254 6684
rect 24820 6616 24900 6644
rect 24820 6604 24826 6616
rect 27522 6604 27528 6656
rect 27580 6604 27586 6656
rect 28718 6604 28724 6656
rect 28776 6644 28782 6656
rect 33704 6644 33732 6820
rect 35176 6789 35204 6820
rect 35268 6888 35808 6916
rect 33781 6783 33839 6789
rect 33781 6749 33793 6783
rect 33827 6780 33839 6783
rect 35161 6783 35219 6789
rect 35268 6786 35296 6888
rect 35802 6876 35808 6888
rect 35860 6876 35866 6928
rect 39022 6916 39028 6928
rect 36924 6888 39028 6916
rect 33827 6752 35081 6780
rect 33827 6749 33839 6752
rect 33781 6743 33839 6749
rect 33965 6715 34023 6721
rect 33965 6681 33977 6715
rect 34011 6681 34023 6715
rect 34146 6712 34152 6724
rect 34107 6684 34152 6712
rect 33965 6675 34023 6681
rect 28776 6616 33732 6644
rect 33980 6644 34008 6675
rect 34146 6672 34152 6684
rect 34204 6672 34210 6724
rect 35053 6712 35081 6752
rect 35161 6749 35173 6783
rect 35207 6749 35219 6783
rect 35161 6743 35219 6749
rect 35253 6780 35311 6786
rect 35253 6746 35265 6780
rect 35299 6746 35311 6780
rect 35253 6740 35311 6746
rect 35345 6783 35403 6789
rect 35345 6749 35357 6783
rect 35391 6749 35403 6783
rect 35526 6780 35532 6792
rect 35487 6752 35532 6780
rect 35345 6743 35403 6749
rect 35360 6712 35388 6743
rect 35526 6740 35532 6752
rect 35584 6740 35590 6792
rect 36633 6783 36691 6789
rect 36633 6749 36645 6783
rect 36679 6749 36691 6783
rect 36814 6780 36820 6792
rect 36775 6752 36820 6780
rect 36633 6743 36691 6749
rect 35053 6684 35388 6712
rect 36648 6712 36676 6743
rect 36814 6740 36820 6752
rect 36872 6740 36878 6792
rect 36924 6789 36952 6888
rect 39022 6876 39028 6888
rect 39080 6876 39086 6928
rect 36909 6783 36967 6789
rect 36909 6749 36921 6783
rect 36955 6749 36967 6783
rect 36909 6743 36967 6749
rect 36998 6740 37004 6792
rect 37056 6780 37062 6792
rect 37737 6783 37795 6789
rect 37737 6780 37749 6783
rect 37056 6752 37749 6780
rect 37056 6740 37062 6752
rect 37737 6749 37749 6752
rect 37783 6749 37795 6783
rect 37737 6743 37795 6749
rect 38562 6740 38568 6792
rect 38620 6789 38626 6792
rect 38620 6783 38669 6789
rect 38620 6749 38623 6783
rect 38657 6749 38669 6783
rect 38620 6743 38669 6749
rect 38749 6783 38807 6789
rect 38749 6749 38761 6783
rect 38795 6749 38807 6783
rect 38749 6743 38807 6749
rect 38620 6740 38626 6743
rect 38102 6712 38108 6724
rect 36648 6684 38108 6712
rect 38102 6672 38108 6684
rect 38160 6712 38166 6724
rect 38764 6712 38792 6743
rect 38838 6740 38844 6792
rect 38896 6789 38902 6792
rect 38896 6780 38904 6789
rect 39025 6783 39083 6789
rect 38896 6752 38941 6780
rect 38896 6743 38904 6752
rect 39025 6749 39037 6783
rect 39071 6749 39083 6783
rect 39025 6743 39083 6749
rect 38896 6740 38902 6743
rect 38930 6712 38936 6724
rect 38160 6684 38654 6712
rect 38764 6684 38936 6712
rect 38160 6672 38166 6684
rect 34514 6644 34520 6656
rect 33980 6616 34520 6644
rect 28776 6604 28782 6616
rect 34514 6604 34520 6616
rect 34572 6604 34578 6656
rect 34885 6647 34943 6653
rect 34885 6613 34897 6647
rect 34931 6644 34943 6647
rect 35434 6644 35440 6656
rect 34931 6616 35440 6644
rect 34931 6613 34943 6616
rect 34885 6607 34943 6613
rect 35434 6604 35440 6616
rect 35492 6604 35498 6656
rect 37277 6647 37335 6653
rect 37277 6613 37289 6647
rect 37323 6644 37335 6647
rect 37550 6644 37556 6656
rect 37323 6616 37556 6644
rect 37323 6613 37335 6616
rect 37277 6607 37335 6613
rect 37550 6604 37556 6616
rect 37608 6604 37614 6656
rect 38378 6644 38384 6656
rect 38339 6616 38384 6644
rect 38378 6604 38384 6616
rect 38436 6604 38442 6656
rect 38626 6644 38654 6684
rect 38930 6672 38936 6684
rect 38988 6672 38994 6724
rect 39040 6644 39068 6743
rect 38626 6616 39068 6644
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 11514 6440 11520 6452
rect 6512 6412 11520 6440
rect 6512 6400 6518 6412
rect 11514 6400 11520 6412
rect 11572 6440 11578 6452
rect 11974 6440 11980 6452
rect 11572 6412 11980 6440
rect 11572 6400 11578 6412
rect 11974 6400 11980 6412
rect 12032 6400 12038 6452
rect 14642 6400 14648 6452
rect 14700 6440 14706 6452
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 14700 6412 15577 6440
rect 14700 6400 14706 6412
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15565 6403 15623 6409
rect 16022 6400 16028 6452
rect 16080 6440 16086 6452
rect 22002 6440 22008 6452
rect 16080 6412 22008 6440
rect 16080 6400 16086 6412
rect 22002 6400 22008 6412
rect 22060 6400 22066 6452
rect 23474 6400 23480 6452
rect 23532 6440 23538 6452
rect 23661 6443 23719 6449
rect 23661 6440 23673 6443
rect 23532 6412 23673 6440
rect 23532 6400 23538 6412
rect 23661 6409 23673 6412
rect 23707 6409 23719 6443
rect 23661 6403 23719 6409
rect 27430 6400 27436 6452
rect 27488 6440 27494 6452
rect 27617 6443 27675 6449
rect 27617 6440 27629 6443
rect 27488 6412 27629 6440
rect 27488 6400 27494 6412
rect 27617 6409 27629 6412
rect 27663 6409 27675 6443
rect 27617 6403 27675 6409
rect 29086 6400 29092 6452
rect 29144 6440 29150 6452
rect 30006 6440 30012 6452
rect 29144 6412 30012 6440
rect 29144 6400 29150 6412
rect 30006 6400 30012 6412
rect 30064 6400 30070 6452
rect 30190 6440 30196 6452
rect 30151 6412 30196 6440
rect 30190 6400 30196 6412
rect 30248 6400 30254 6452
rect 34146 6400 34152 6452
rect 34204 6440 34210 6452
rect 34204 6412 36492 6440
rect 34204 6400 34210 6412
rect 36464 6384 36492 6412
rect 36814 6400 36820 6452
rect 36872 6440 36878 6452
rect 37277 6443 37335 6449
rect 37277 6440 37289 6443
rect 36872 6412 37289 6440
rect 36872 6400 36878 6412
rect 37277 6409 37289 6412
rect 37323 6409 37335 6443
rect 39666 6440 39672 6452
rect 39627 6412 39672 6440
rect 37277 6403 37335 6409
rect 39666 6400 39672 6412
rect 39724 6400 39730 6452
rect 3237 6375 3295 6381
rect 3237 6341 3249 6375
rect 3283 6372 3295 6375
rect 3786 6372 3792 6384
rect 3283 6344 3792 6372
rect 3283 6341 3295 6344
rect 3237 6335 3295 6341
rect 3786 6332 3792 6344
rect 3844 6332 3850 6384
rect 4985 6375 5043 6381
rect 4985 6341 4997 6375
rect 5031 6372 5043 6375
rect 5534 6372 5540 6384
rect 5031 6344 5540 6372
rect 5031 6341 5043 6344
rect 4985 6335 5043 6341
rect 5534 6332 5540 6344
rect 5592 6372 5598 6384
rect 6270 6372 6276 6384
rect 5592 6344 6276 6372
rect 5592 6332 5598 6344
rect 6270 6332 6276 6344
rect 6328 6332 6334 6384
rect 9858 6381 9864 6384
rect 9852 6372 9864 6381
rect 9819 6344 9864 6372
rect 9852 6335 9864 6344
rect 9858 6332 9864 6335
rect 9916 6332 9922 6384
rect 19058 6372 19064 6384
rect 13740 6344 19064 6372
rect 2498 6304 2504 6316
rect 2459 6276 2504 6304
rect 2498 6264 2504 6276
rect 2556 6264 2562 6316
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5408 6276 5641 6304
rect 5408 6264 5414 6276
rect 5629 6273 5641 6276
rect 5675 6273 5687 6307
rect 5629 6267 5687 6273
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6273 5871 6307
rect 5813 6267 5871 6273
rect 6457 6307 6515 6313
rect 6457 6273 6469 6307
rect 6503 6304 6515 6307
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 6503 6276 6929 6304
rect 6503 6273 6515 6276
rect 6457 6267 6515 6273
rect 6917 6273 6929 6276
rect 6963 6304 6975 6307
rect 7374 6304 7380 6316
rect 6963 6276 7380 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 5828 6236 5856 6267
rect 7374 6264 7380 6276
rect 7432 6264 7438 6316
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7650 6304 7656 6316
rect 7607 6276 7656 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6304 8447 6307
rect 8478 6304 8484 6316
rect 8435 6276 8484 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 9030 6304 9036 6316
rect 8991 6276 9036 6304
rect 9030 6264 9036 6276
rect 9088 6264 9094 6316
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 13740 6313 13768 6344
rect 19058 6332 19064 6344
rect 19116 6332 19122 6384
rect 19334 6332 19340 6384
rect 19392 6372 19398 6384
rect 19518 6372 19524 6384
rect 19392 6344 19524 6372
rect 19392 6332 19398 6344
rect 19518 6332 19524 6344
rect 19576 6332 19582 6384
rect 22186 6332 22192 6384
rect 22244 6372 22250 6384
rect 23293 6375 23351 6381
rect 23293 6372 23305 6375
rect 22244 6344 23305 6372
rect 22244 6332 22250 6344
rect 23293 6341 23305 6344
rect 23339 6341 23351 6375
rect 23293 6335 23351 6341
rect 23385 6375 23443 6381
rect 23385 6341 23397 6375
rect 23431 6372 23443 6375
rect 23750 6372 23756 6384
rect 23431 6344 23756 6372
rect 23431 6341 23443 6344
rect 23385 6335 23443 6341
rect 23750 6332 23756 6344
rect 23808 6332 23814 6384
rect 30837 6375 30895 6381
rect 30837 6341 30849 6375
rect 30883 6372 30895 6375
rect 33134 6372 33140 6384
rect 30883 6344 33140 6372
rect 30883 6341 30895 6344
rect 30837 6335 30895 6341
rect 33134 6332 33140 6344
rect 33192 6332 33198 6384
rect 34422 6372 34428 6384
rect 34383 6344 34428 6372
rect 34422 6332 34428 6344
rect 34480 6372 34486 6384
rect 35802 6372 35808 6384
rect 34480 6344 35296 6372
rect 34480 6332 34486 6344
rect 13998 6313 14004 6316
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 9456 6276 9597 6304
rect 9456 6264 9462 6276
rect 9585 6273 9597 6276
rect 9631 6273 9643 6307
rect 13725 6307 13783 6313
rect 9585 6267 9643 6273
rect 9692 6276 12434 6304
rect 6822 6236 6828 6248
rect 5828 6208 6828 6236
rect 6822 6196 6828 6208
rect 6880 6196 6886 6248
rect 8018 6236 8024 6248
rect 7024 6208 8024 6236
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 7024 6168 7052 6208
rect 8018 6196 8024 6208
rect 8076 6236 8082 6248
rect 9692 6236 9720 6276
rect 8076 6208 9720 6236
rect 8076 6196 8082 6208
rect 6052 6140 7052 6168
rect 7101 6171 7159 6177
rect 6052 6128 6058 6140
rect 7101 6137 7113 6171
rect 7147 6168 7159 6171
rect 8662 6168 8668 6180
rect 7147 6140 8668 6168
rect 7147 6137 7159 6140
rect 7101 6131 7159 6137
rect 8662 6128 8668 6140
rect 8720 6128 8726 6180
rect 10965 6171 11023 6177
rect 10965 6137 10977 6171
rect 11011 6168 11023 6171
rect 11054 6168 11060 6180
rect 11011 6140 11060 6168
rect 11011 6137 11023 6140
rect 10965 6131 11023 6137
rect 11054 6128 11060 6140
rect 11112 6168 11118 6180
rect 11974 6168 11980 6180
rect 11112 6140 11980 6168
rect 11112 6128 11118 6140
rect 11974 6128 11980 6140
rect 12032 6128 12038 6180
rect 12406 6168 12434 6276
rect 13725 6273 13737 6307
rect 13771 6273 13783 6307
rect 13992 6304 14004 6313
rect 13959 6276 14004 6304
rect 13725 6267 13783 6273
rect 13992 6267 14004 6276
rect 13998 6264 14004 6267
rect 14056 6264 14062 6316
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6304 15807 6307
rect 15933 6307 15991 6313
rect 15795 6276 15884 6304
rect 15795 6273 15807 6276
rect 15749 6267 15807 6273
rect 15746 6168 15752 6180
rect 12406 6140 13768 6168
rect 1857 6103 1915 6109
rect 1857 6069 1869 6103
rect 1903 6100 1915 6103
rect 2038 6100 2044 6112
rect 1903 6072 2044 6100
rect 1903 6069 1915 6072
rect 1857 6063 1915 6069
rect 2038 6060 2044 6072
rect 2096 6060 2102 6112
rect 2130 6060 2136 6112
rect 2188 6100 2194 6112
rect 2317 6103 2375 6109
rect 2317 6100 2329 6103
rect 2188 6072 2329 6100
rect 2188 6060 2194 6072
rect 2317 6069 2329 6072
rect 2363 6069 2375 6103
rect 5626 6100 5632 6112
rect 5587 6072 5632 6100
rect 2317 6063 2375 6069
rect 5626 6060 5632 6072
rect 5684 6060 5690 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 7616 6072 7757 6100
rect 7616 6060 7622 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 7892 6072 8217 6100
rect 7892 6060 7898 6072
rect 8205 6069 8217 6072
rect 8251 6069 8263 6103
rect 8846 6100 8852 6112
rect 8807 6072 8852 6100
rect 8205 6063 8263 6069
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 11606 6100 11612 6112
rect 11567 6072 11612 6100
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 12158 6060 12164 6112
rect 12216 6100 12222 6112
rect 12253 6103 12311 6109
rect 12253 6100 12265 6103
rect 12216 6072 12265 6100
rect 12216 6060 12222 6072
rect 12253 6069 12265 6072
rect 12299 6069 12311 6103
rect 12253 6063 12311 6069
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 13081 6103 13139 6109
rect 13081 6100 13093 6103
rect 13044 6072 13093 6100
rect 13044 6060 13050 6072
rect 13081 6069 13093 6072
rect 13127 6069 13139 6103
rect 13740 6100 13768 6140
rect 15028 6140 15752 6168
rect 15028 6100 15056 6140
rect 15746 6128 15752 6140
rect 15804 6128 15810 6180
rect 13740 6072 15056 6100
rect 15105 6103 15163 6109
rect 13081 6063 13139 6069
rect 15105 6069 15117 6103
rect 15151 6100 15163 6103
rect 15856 6100 15884 6276
rect 15933 6273 15945 6307
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 15948 6236 15976 6267
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16632 6276 16865 6304
rect 16632 6264 16638 6276
rect 16853 6273 16865 6276
rect 16899 6304 16911 6307
rect 17313 6307 17371 6313
rect 17313 6304 17325 6307
rect 16899 6276 17325 6304
rect 16899 6273 16911 6276
rect 16853 6267 16911 6273
rect 17313 6273 17325 6276
rect 17359 6273 17371 6307
rect 17313 6267 17371 6273
rect 19705 6307 19763 6313
rect 19705 6273 19717 6307
rect 19751 6304 19763 6307
rect 20622 6304 20628 6316
rect 19751 6276 20628 6304
rect 19751 6273 19763 6276
rect 19705 6267 19763 6273
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 23106 6304 23112 6316
rect 23067 6276 23112 6304
rect 23106 6264 23112 6276
rect 23164 6264 23170 6316
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6273 23535 6307
rect 23477 6267 23535 6273
rect 24673 6307 24731 6313
rect 24673 6273 24685 6307
rect 24719 6304 24731 6307
rect 24854 6304 24860 6316
rect 24719 6276 24860 6304
rect 24719 6273 24731 6276
rect 24673 6267 24731 6273
rect 17034 6236 17040 6248
rect 15948 6208 17040 6236
rect 17034 6196 17040 6208
rect 17092 6196 17098 6248
rect 18598 6196 18604 6248
rect 18656 6236 18662 6248
rect 21634 6236 21640 6248
rect 18656 6208 21640 6236
rect 18656 6196 18662 6208
rect 21634 6196 21640 6208
rect 21692 6236 21698 6248
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 21692 6208 21833 6236
rect 21692 6196 21698 6208
rect 21821 6205 21833 6208
rect 21867 6205 21879 6239
rect 21821 6199 21879 6205
rect 22097 6239 22155 6245
rect 22097 6205 22109 6239
rect 22143 6236 22155 6239
rect 22186 6236 22192 6248
rect 22143 6208 22192 6236
rect 22143 6205 22155 6208
rect 22097 6199 22155 6205
rect 22186 6196 22192 6208
rect 22244 6196 22250 6248
rect 22830 6196 22836 6248
rect 22888 6236 22894 6248
rect 23492 6236 23520 6267
rect 24854 6264 24860 6276
rect 24912 6264 24918 6316
rect 26970 6304 26976 6316
rect 26931 6276 26976 6304
rect 26970 6264 26976 6276
rect 27028 6264 27034 6316
rect 27522 6264 27528 6316
rect 27580 6304 27586 6316
rect 29546 6304 29552 6316
rect 27580 6276 29552 6304
rect 27580 6264 27586 6276
rect 29546 6264 29552 6276
rect 29604 6264 29610 6316
rect 29638 6264 29644 6316
rect 29696 6304 29702 6316
rect 30006 6313 30012 6316
rect 29733 6307 29791 6313
rect 29733 6304 29745 6307
rect 29696 6276 29745 6304
rect 29696 6264 29702 6276
rect 29733 6273 29745 6276
rect 29779 6273 29791 6307
rect 29733 6267 29791 6273
rect 29825 6307 29883 6313
rect 29825 6273 29837 6307
rect 29871 6273 29883 6307
rect 29825 6267 29883 6273
rect 29963 6307 30012 6313
rect 29963 6273 29975 6307
rect 30009 6273 30012 6307
rect 29963 6267 30012 6273
rect 22888 6208 23520 6236
rect 24213 6239 24271 6245
rect 22888 6196 22894 6208
rect 24213 6205 24225 6239
rect 24259 6236 24271 6239
rect 24578 6236 24584 6248
rect 24259 6208 24584 6236
rect 24259 6205 24271 6208
rect 24213 6199 24271 6205
rect 24578 6196 24584 6208
rect 24636 6236 24642 6248
rect 28718 6236 28724 6248
rect 24636 6208 28724 6236
rect 24636 6196 24642 6208
rect 28718 6196 28724 6208
rect 28776 6196 28782 6248
rect 28810 6196 28816 6248
rect 28868 6236 28874 6248
rect 28997 6239 29055 6245
rect 28997 6236 29009 6239
rect 28868 6208 29009 6236
rect 28868 6196 28874 6208
rect 28997 6205 29009 6208
rect 29043 6236 29055 6239
rect 29086 6236 29092 6248
rect 29043 6208 29092 6236
rect 29043 6205 29055 6208
rect 28997 6199 29055 6205
rect 29086 6196 29092 6208
rect 29144 6196 29150 6248
rect 29843 6180 29871 6267
rect 30006 6264 30012 6267
rect 30064 6264 30070 6316
rect 31021 6307 31079 6313
rect 31021 6273 31033 6307
rect 31067 6304 31079 6307
rect 31110 6304 31116 6316
rect 31067 6276 31116 6304
rect 31067 6273 31079 6276
rect 31021 6267 31079 6273
rect 31110 6264 31116 6276
rect 31168 6264 31174 6316
rect 35268 6313 35296 6344
rect 35360 6344 35808 6372
rect 35360 6313 35388 6344
rect 35802 6332 35808 6344
rect 35860 6332 35866 6384
rect 36262 6372 36268 6384
rect 36223 6344 36268 6372
rect 36262 6332 36268 6344
rect 36320 6332 36326 6384
rect 36446 6372 36452 6384
rect 36407 6344 36452 6372
rect 36446 6332 36452 6344
rect 36504 6332 36510 6384
rect 37642 6372 37648 6384
rect 37603 6344 37648 6372
rect 37642 6332 37648 6344
rect 37700 6332 37706 6384
rect 38378 6332 38384 6384
rect 38436 6372 38442 6384
rect 38534 6375 38592 6381
rect 38534 6372 38546 6375
rect 38436 6344 38546 6372
rect 38436 6332 38442 6344
rect 38534 6341 38546 6344
rect 38580 6341 38592 6375
rect 38534 6335 38592 6341
rect 35253 6307 35311 6313
rect 35253 6273 35265 6307
rect 35299 6273 35311 6307
rect 35253 6267 35311 6273
rect 35345 6307 35403 6313
rect 35345 6273 35357 6307
rect 35391 6273 35403 6307
rect 35345 6267 35403 6273
rect 35437 6307 35495 6313
rect 35437 6273 35449 6307
rect 35483 6273 35495 6307
rect 35437 6267 35495 6273
rect 18506 6128 18512 6180
rect 18564 6168 18570 6180
rect 18564 6140 21312 6168
rect 18564 6128 18570 6140
rect 18690 6100 18696 6112
rect 15151 6072 18696 6100
rect 15151 6069 15163 6072
rect 15105 6063 15163 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 19889 6103 19947 6109
rect 19889 6069 19901 6103
rect 19935 6100 19947 6103
rect 20070 6100 20076 6112
rect 19935 6072 20076 6100
rect 19935 6069 19947 6072
rect 19889 6063 19947 6069
rect 20070 6060 20076 6072
rect 20128 6060 20134 6112
rect 20717 6103 20775 6109
rect 20717 6069 20729 6103
rect 20763 6100 20775 6103
rect 20806 6100 20812 6112
rect 20763 6072 20812 6100
rect 20763 6069 20775 6072
rect 20717 6063 20775 6069
rect 20806 6060 20812 6072
rect 20864 6060 20870 6112
rect 21174 6100 21180 6112
rect 21135 6072 21180 6100
rect 21174 6060 21180 6072
rect 21232 6060 21238 6112
rect 21284 6100 21312 6140
rect 22002 6128 22008 6180
rect 22060 6168 22066 6180
rect 25590 6168 25596 6180
rect 22060 6140 25596 6168
rect 22060 6128 22066 6140
rect 25590 6128 25596 6140
rect 25648 6128 25654 6180
rect 27157 6171 27215 6177
rect 25700 6140 26280 6168
rect 23106 6100 23112 6112
rect 21284 6072 23112 6100
rect 23106 6060 23112 6072
rect 23164 6060 23170 6112
rect 23382 6060 23388 6112
rect 23440 6100 23446 6112
rect 25700 6100 25728 6140
rect 26142 6100 26148 6112
rect 23440 6072 25728 6100
rect 26103 6072 26148 6100
rect 23440 6060 23446 6072
rect 26142 6060 26148 6072
rect 26200 6060 26206 6112
rect 26252 6100 26280 6140
rect 27157 6137 27169 6171
rect 27203 6168 27215 6171
rect 28166 6168 28172 6180
rect 27203 6140 28172 6168
rect 27203 6137 27215 6140
rect 27157 6131 27215 6137
rect 28166 6128 28172 6140
rect 28224 6128 28230 6180
rect 29822 6128 29828 6180
rect 29880 6128 29886 6180
rect 35268 6168 35296 6267
rect 35452 6236 35480 6267
rect 35526 6264 35532 6316
rect 35584 6304 35590 6316
rect 35621 6307 35679 6313
rect 35621 6304 35633 6307
rect 35584 6276 35633 6304
rect 35584 6264 35590 6276
rect 35621 6273 35633 6276
rect 35667 6273 35679 6307
rect 35621 6267 35679 6273
rect 37182 6264 37188 6316
rect 37240 6304 37246 6316
rect 37461 6307 37519 6313
rect 37461 6304 37473 6307
rect 37240 6276 37473 6304
rect 37240 6264 37246 6276
rect 37461 6273 37473 6276
rect 37507 6273 37519 6307
rect 37461 6267 37519 6273
rect 37918 6264 37924 6316
rect 37976 6304 37982 6316
rect 38289 6307 38347 6313
rect 38289 6304 38301 6307
rect 37976 6276 38301 6304
rect 37976 6264 37982 6276
rect 38289 6273 38301 6276
rect 38335 6273 38347 6307
rect 38289 6267 38347 6273
rect 36081 6239 36139 6245
rect 36081 6236 36093 6239
rect 35452 6208 36093 6236
rect 36081 6205 36093 6208
rect 36127 6205 36139 6239
rect 36081 6199 36139 6205
rect 36998 6168 37004 6180
rect 35268 6140 37004 6168
rect 36998 6128 37004 6140
rect 37056 6128 37062 6180
rect 58158 6168 58164 6180
rect 58119 6140 58164 6168
rect 58158 6128 58164 6140
rect 58216 6128 58222 6180
rect 29362 6100 29368 6112
rect 26252 6072 29368 6100
rect 29362 6060 29368 6072
rect 29420 6060 29426 6112
rect 30190 6060 30196 6112
rect 30248 6100 30254 6112
rect 30653 6103 30711 6109
rect 30653 6100 30665 6103
rect 30248 6072 30665 6100
rect 30248 6060 30254 6072
rect 30653 6069 30665 6072
rect 30699 6069 30711 6103
rect 30653 6063 30711 6069
rect 34698 6060 34704 6112
rect 34756 6100 34762 6112
rect 34977 6103 35035 6109
rect 34977 6100 34989 6103
rect 34756 6072 34989 6100
rect 34756 6060 34762 6072
rect 34977 6069 34989 6072
rect 35023 6069 35035 6103
rect 34977 6063 35035 6069
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 5721 5899 5779 5905
rect 5721 5865 5733 5899
rect 5767 5896 5779 5899
rect 6914 5896 6920 5908
rect 5767 5868 6920 5896
rect 5767 5865 5779 5868
rect 5721 5859 5779 5865
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 12434 5896 12440 5908
rect 7300 5868 12440 5896
rect 3237 5831 3295 5837
rect 3237 5797 3249 5831
rect 3283 5828 3295 5831
rect 3283 5800 4292 5828
rect 3283 5797 3295 5800
rect 3237 5791 3295 5797
rect 4264 5769 4292 5800
rect 4798 5788 4804 5840
rect 4856 5828 4862 5840
rect 7300 5837 7328 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 12529 5899 12587 5905
rect 12529 5865 12541 5899
rect 12575 5896 12587 5899
rect 18598 5896 18604 5908
rect 12575 5868 18604 5896
rect 12575 5865 12587 5868
rect 12529 5859 12587 5865
rect 18598 5856 18604 5868
rect 18656 5856 18662 5908
rect 18693 5899 18751 5905
rect 18693 5865 18705 5899
rect 18739 5896 18751 5899
rect 19426 5896 19432 5908
rect 18739 5868 19432 5896
rect 18739 5865 18751 5868
rect 18693 5859 18751 5865
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 20622 5896 20628 5908
rect 20583 5868 20628 5896
rect 20622 5856 20628 5868
rect 20680 5896 20686 5908
rect 22649 5899 22707 5905
rect 20680 5868 22094 5896
rect 20680 5856 20686 5868
rect 7285 5831 7343 5837
rect 7285 5828 7297 5831
rect 4856 5800 7297 5828
rect 4856 5788 4862 5800
rect 7285 5797 7297 5800
rect 7331 5797 7343 5831
rect 7285 5791 7343 5797
rect 10137 5831 10195 5837
rect 10137 5797 10149 5831
rect 10183 5828 10195 5831
rect 10778 5828 10784 5840
rect 10183 5800 10784 5828
rect 10183 5797 10195 5800
rect 10137 5791 10195 5797
rect 10778 5788 10784 5800
rect 10836 5788 10842 5840
rect 11330 5828 11336 5840
rect 11291 5800 11336 5828
rect 11330 5788 11336 5800
rect 11388 5788 11394 5840
rect 16209 5831 16267 5837
rect 16209 5828 16221 5831
rect 15221 5800 16221 5828
rect 4249 5763 4307 5769
rect 4249 5729 4261 5763
rect 4295 5729 4307 5763
rect 4249 5723 4307 5729
rect 4433 5763 4491 5769
rect 4433 5729 4445 5763
rect 4479 5760 4491 5763
rect 4706 5760 4712 5772
rect 4479 5732 4712 5760
rect 4479 5729 4491 5732
rect 4433 5723 4491 5729
rect 1854 5692 1860 5704
rect 1815 5664 1860 5692
rect 1854 5652 1860 5664
rect 1912 5652 1918 5704
rect 2130 5701 2136 5704
rect 2124 5692 2136 5701
rect 2091 5664 2136 5692
rect 2124 5655 2136 5664
rect 2130 5652 2136 5655
rect 2188 5652 2194 5704
rect 3234 5652 3240 5704
rect 3292 5692 3298 5704
rect 4264 5692 4292 5723
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5760 5595 5763
rect 6546 5760 6552 5772
rect 5583 5732 6552 5760
rect 5583 5729 5595 5732
rect 5537 5723 5595 5729
rect 6546 5720 6552 5732
rect 6604 5720 6610 5772
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5760 9551 5763
rect 10226 5760 10232 5772
rect 9539 5732 10232 5760
rect 9539 5729 9551 5732
rect 9493 5723 9551 5729
rect 10226 5720 10232 5732
rect 10284 5720 10290 5772
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 3292 5664 4200 5692
rect 4264 5664 5457 5692
rect 3292 5652 3298 5664
rect 2682 5584 2688 5636
rect 2740 5624 2746 5636
rect 4172 5633 4200 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 6362 5692 6368 5704
rect 6323 5664 6368 5692
rect 5445 5655 5503 5661
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5692 8447 5695
rect 9950 5692 9956 5704
rect 8435 5664 9956 5692
rect 8435 5661 8447 5664
rect 8389 5655 8447 5661
rect 9950 5652 9956 5664
rect 10008 5652 10014 5704
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5692 10839 5695
rect 11330 5692 11336 5704
rect 10827 5664 11336 5692
rect 10827 5661 10839 5664
rect 10781 5655 10839 5661
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 11514 5692 11520 5704
rect 11475 5664 11520 5692
rect 11514 5652 11520 5664
rect 11572 5652 11578 5704
rect 12529 5695 12587 5701
rect 12529 5692 12541 5695
rect 12406 5664 12541 5692
rect 4157 5627 4215 5633
rect 2740 5596 3832 5624
rect 2740 5584 2746 5596
rect 3804 5565 3832 5596
rect 4157 5593 4169 5627
rect 4203 5624 4215 5627
rect 6549 5627 6607 5633
rect 6549 5624 6561 5627
rect 4203 5596 6561 5624
rect 4203 5593 4215 5596
rect 4157 5587 4215 5593
rect 6549 5593 6561 5596
rect 6595 5624 6607 5627
rect 6638 5624 6644 5636
rect 6595 5596 6644 5624
rect 6595 5593 6607 5596
rect 6549 5587 6607 5593
rect 6638 5584 6644 5596
rect 6696 5584 6702 5636
rect 7006 5584 7012 5636
rect 7064 5624 7070 5636
rect 7101 5627 7159 5633
rect 7101 5624 7113 5627
rect 7064 5596 7113 5624
rect 7064 5584 7070 5596
rect 7101 5593 7113 5596
rect 7147 5593 7159 5627
rect 7101 5587 7159 5593
rect 8294 5584 8300 5636
rect 8352 5624 8358 5636
rect 12406 5624 12434 5664
rect 12529 5661 12541 5664
rect 12575 5661 12587 5695
rect 12710 5692 12716 5704
rect 12671 5664 12716 5692
rect 12529 5655 12587 5661
rect 12710 5652 12716 5664
rect 12768 5652 12774 5704
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 13320 5664 13369 5692
rect 13320 5652 13326 5664
rect 13357 5661 13369 5664
rect 13403 5661 13415 5695
rect 14090 5692 14096 5704
rect 14051 5664 14096 5692
rect 13357 5655 13415 5661
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 14918 5652 14924 5704
rect 14976 5692 14982 5704
rect 15105 5695 15163 5701
rect 15105 5692 15117 5695
rect 14976 5664 15117 5692
rect 14976 5652 14982 5664
rect 15105 5661 15117 5664
rect 15151 5661 15163 5695
rect 15105 5655 15163 5661
rect 15221 5686 15249 5800
rect 16209 5797 16221 5800
rect 16255 5797 16267 5831
rect 22066 5828 22094 5868
rect 22649 5865 22661 5899
rect 22695 5896 22707 5899
rect 23290 5896 23296 5908
rect 22695 5868 23296 5896
rect 22695 5865 22707 5868
rect 22649 5859 22707 5865
rect 23290 5856 23296 5868
rect 23348 5856 23354 5908
rect 24762 5896 24768 5908
rect 24723 5868 24768 5896
rect 24762 5856 24768 5868
rect 24820 5856 24826 5908
rect 29178 5856 29184 5908
rect 29236 5896 29242 5908
rect 29549 5899 29607 5905
rect 29549 5896 29561 5899
rect 29236 5868 29561 5896
rect 29236 5856 29242 5868
rect 29549 5865 29561 5868
rect 29595 5896 29607 5899
rect 30558 5896 30564 5908
rect 29595 5868 30564 5896
rect 29595 5865 29607 5868
rect 29549 5859 29607 5865
rect 30558 5856 30564 5868
rect 30616 5856 30622 5908
rect 32677 5899 32735 5905
rect 32677 5865 32689 5899
rect 32723 5896 32735 5899
rect 33134 5896 33140 5908
rect 32723 5868 33140 5896
rect 32723 5865 32735 5868
rect 32677 5859 32735 5865
rect 33134 5856 33140 5868
rect 33192 5856 33198 5908
rect 34514 5856 34520 5908
rect 34572 5896 34578 5908
rect 35526 5896 35532 5908
rect 34572 5868 35532 5896
rect 34572 5856 34578 5868
rect 35526 5856 35532 5868
rect 35584 5856 35590 5908
rect 36173 5899 36231 5905
rect 36173 5865 36185 5899
rect 36219 5896 36231 5899
rect 36262 5896 36268 5908
rect 36219 5868 36268 5896
rect 36219 5865 36231 5868
rect 36173 5859 36231 5865
rect 36262 5856 36268 5868
rect 36320 5856 36326 5908
rect 37182 5856 37188 5908
rect 37240 5896 37246 5908
rect 38841 5899 38899 5905
rect 38841 5896 38853 5899
rect 37240 5868 38853 5896
rect 37240 5856 37246 5868
rect 38841 5865 38853 5868
rect 38887 5865 38899 5899
rect 38841 5859 38899 5865
rect 27706 5828 27712 5840
rect 22066 5800 27712 5828
rect 16209 5791 16267 5797
rect 27706 5788 27712 5800
rect 27764 5788 27770 5840
rect 15746 5720 15752 5772
rect 15804 5760 15810 5772
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 15804 5732 17601 5760
rect 15804 5720 15810 5732
rect 17589 5729 17601 5732
rect 17635 5760 17647 5763
rect 17862 5760 17868 5772
rect 17635 5732 17868 5760
rect 17635 5729 17647 5732
rect 17589 5723 17647 5729
rect 17862 5720 17868 5732
rect 17920 5760 17926 5772
rect 17920 5732 18460 5760
rect 17920 5720 17926 5732
rect 15289 5695 15347 5701
rect 15289 5686 15301 5695
rect 15221 5661 15301 5686
rect 15335 5661 15347 5695
rect 15221 5658 15347 5661
rect 15289 5655 15347 5658
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 8352 5596 12434 5624
rect 8352 5584 8358 5596
rect 14550 5584 14556 5636
rect 14608 5624 14614 5636
rect 15396 5624 15424 5655
rect 15470 5652 15476 5704
rect 15528 5692 15534 5704
rect 15528 5664 15573 5692
rect 15528 5652 15534 5664
rect 17770 5652 17776 5704
rect 17828 5692 17834 5704
rect 18049 5695 18107 5701
rect 18049 5692 18061 5695
rect 17828 5664 18061 5692
rect 17828 5652 17834 5664
rect 18049 5661 18061 5664
rect 18095 5661 18107 5695
rect 18230 5692 18236 5704
rect 18191 5664 18236 5692
rect 18049 5655 18107 5661
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 18432 5701 18460 5732
rect 19058 5720 19064 5772
rect 19116 5760 19122 5772
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 19116 5732 19257 5760
rect 19116 5720 19122 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 23201 5763 23259 5769
rect 23201 5729 23213 5763
rect 23247 5760 23259 5763
rect 23382 5760 23388 5772
rect 23247 5732 23388 5760
rect 23247 5729 23259 5732
rect 23201 5723 23259 5729
rect 23382 5720 23388 5732
rect 23440 5720 23446 5772
rect 25590 5760 25596 5772
rect 25551 5732 25596 5760
rect 25590 5720 25596 5732
rect 25648 5720 25654 5772
rect 30190 5720 30196 5772
rect 30248 5720 30254 5772
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5661 18475 5695
rect 18417 5655 18475 5661
rect 14608 5596 15424 5624
rect 16393 5627 16451 5633
rect 14608 5584 14614 5596
rect 16393 5593 16405 5627
rect 16439 5593 16451 5627
rect 16393 5587 16451 5593
rect 16577 5627 16635 5633
rect 16577 5593 16589 5627
rect 16623 5624 16635 5627
rect 17034 5624 17040 5636
rect 16623 5596 17040 5624
rect 16623 5593 16635 5596
rect 16577 5587 16635 5593
rect 3789 5559 3847 5565
rect 3789 5525 3801 5559
rect 3835 5525 3847 5559
rect 3789 5519 3847 5525
rect 4982 5516 4988 5568
rect 5040 5556 5046 5568
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 5040 5528 5089 5556
rect 5040 5516 5046 5528
rect 5077 5525 5089 5528
rect 5123 5525 5135 5559
rect 5077 5519 5135 5525
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 11977 5559 12035 5565
rect 11977 5556 11989 5559
rect 5500 5528 11989 5556
rect 5500 5516 5506 5528
rect 11977 5525 11989 5528
rect 12023 5556 12035 5559
rect 14826 5556 14832 5568
rect 12023 5528 14832 5556
rect 12023 5525 12035 5528
rect 11977 5519 12035 5525
rect 14826 5516 14832 5528
rect 14884 5516 14890 5568
rect 15749 5559 15807 5565
rect 15749 5525 15761 5559
rect 15795 5556 15807 5559
rect 16114 5556 16120 5568
rect 15795 5528 16120 5556
rect 15795 5525 15807 5528
rect 15749 5519 15807 5525
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 16408 5556 16436 5587
rect 17034 5584 17040 5596
rect 17092 5584 17098 5636
rect 17678 5584 17684 5636
rect 17736 5624 17742 5636
rect 18138 5624 18144 5636
rect 17736 5596 18144 5624
rect 17736 5584 17742 5596
rect 18138 5584 18144 5596
rect 18196 5624 18202 5636
rect 18340 5624 18368 5655
rect 18690 5652 18696 5704
rect 18748 5692 18754 5704
rect 22097 5695 22155 5701
rect 22097 5692 22109 5695
rect 18748 5664 22109 5692
rect 18748 5652 18754 5664
rect 22097 5661 22109 5664
rect 22143 5661 22155 5695
rect 22097 5655 22155 5661
rect 22186 5652 22192 5704
rect 22244 5692 22250 5704
rect 22281 5695 22339 5701
rect 22281 5692 22293 5695
rect 22244 5664 22293 5692
rect 22244 5652 22250 5664
rect 22281 5661 22293 5664
rect 22327 5661 22339 5695
rect 22281 5655 22339 5661
rect 22465 5695 22523 5701
rect 22465 5661 22477 5695
rect 22511 5692 22523 5695
rect 22830 5692 22836 5704
rect 22511 5664 22836 5692
rect 22511 5661 22523 5664
rect 22465 5655 22523 5661
rect 22830 5652 22836 5664
rect 22888 5652 22894 5704
rect 23750 5652 23756 5704
rect 23808 5692 23814 5704
rect 24581 5695 24639 5701
rect 24581 5692 24593 5695
rect 23808 5664 24593 5692
rect 23808 5652 23814 5664
rect 24581 5661 24593 5664
rect 24627 5661 24639 5695
rect 24581 5655 24639 5661
rect 25869 5695 25927 5701
rect 25869 5661 25881 5695
rect 25915 5692 25927 5695
rect 27522 5692 27528 5704
rect 25915 5664 27528 5692
rect 25915 5661 25927 5664
rect 25869 5655 25927 5661
rect 27522 5652 27528 5664
rect 27580 5652 27586 5704
rect 29546 5652 29552 5704
rect 29604 5692 29610 5704
rect 30101 5695 30159 5701
rect 30101 5692 30113 5695
rect 29604 5664 30113 5692
rect 29604 5652 29610 5664
rect 30101 5661 30113 5664
rect 30147 5661 30159 5695
rect 30208 5689 30236 5720
rect 30558 5701 30564 5704
rect 30285 5695 30343 5701
rect 30285 5689 30297 5695
rect 30208 5661 30297 5689
rect 30331 5661 30343 5695
rect 30101 5655 30159 5661
rect 30285 5655 30343 5661
rect 30377 5695 30435 5701
rect 30377 5661 30389 5695
rect 30423 5661 30435 5695
rect 30377 5655 30435 5661
rect 30515 5695 30564 5701
rect 30515 5661 30527 5695
rect 30561 5661 30564 5695
rect 30515 5655 30564 5661
rect 18196 5596 18368 5624
rect 18196 5584 18202 5596
rect 19334 5584 19340 5636
rect 19392 5624 19398 5636
rect 19490 5627 19548 5633
rect 19490 5624 19502 5627
rect 19392 5596 19502 5624
rect 19392 5584 19398 5596
rect 19490 5593 19502 5596
rect 19536 5593 19548 5627
rect 19490 5587 19548 5593
rect 22373 5627 22431 5633
rect 22373 5593 22385 5627
rect 22419 5624 22431 5627
rect 22922 5624 22928 5636
rect 22419 5596 22928 5624
rect 22419 5593 22431 5596
rect 22373 5587 22431 5593
rect 22922 5584 22928 5596
rect 22980 5584 22986 5636
rect 24394 5624 24400 5636
rect 24355 5596 24400 5624
rect 24394 5584 24400 5596
rect 24452 5584 24458 5636
rect 27062 5584 27068 5636
rect 27120 5624 27126 5636
rect 29822 5624 29828 5636
rect 27120 5596 29828 5624
rect 27120 5584 27126 5596
rect 29822 5584 29828 5596
rect 29880 5624 29886 5636
rect 30392 5624 30420 5655
rect 30558 5652 30564 5655
rect 30616 5652 30622 5704
rect 31018 5652 31024 5704
rect 31076 5692 31082 5704
rect 31297 5695 31355 5701
rect 31297 5692 31309 5695
rect 31076 5664 31309 5692
rect 31076 5652 31082 5664
rect 31297 5661 31309 5664
rect 31343 5692 31355 5695
rect 34790 5692 34796 5704
rect 31343 5664 34796 5692
rect 31343 5661 31355 5664
rect 31297 5655 31355 5661
rect 34790 5652 34796 5664
rect 34848 5692 34854 5704
rect 37461 5695 37519 5701
rect 37461 5692 37473 5695
rect 34848 5664 37473 5692
rect 34848 5652 34854 5664
rect 37461 5661 37473 5664
rect 37507 5661 37519 5695
rect 37461 5655 37519 5661
rect 37550 5652 37556 5704
rect 37608 5692 37614 5704
rect 37717 5695 37775 5701
rect 37717 5692 37729 5695
rect 37608 5664 37729 5692
rect 37608 5652 37614 5664
rect 37717 5661 37729 5664
rect 37763 5661 37775 5695
rect 37717 5655 37775 5661
rect 29880 5596 30420 5624
rect 30745 5627 30803 5633
rect 29880 5584 29886 5596
rect 30300 5568 30328 5596
rect 30745 5593 30757 5627
rect 30791 5624 30803 5627
rect 31542 5627 31600 5633
rect 31542 5624 31554 5627
rect 30791 5596 31554 5624
rect 30791 5593 30803 5596
rect 30745 5587 30803 5593
rect 31542 5593 31554 5596
rect 31588 5593 31600 5627
rect 31542 5587 31600 5593
rect 34698 5584 34704 5636
rect 34756 5624 34762 5636
rect 35038 5627 35096 5633
rect 35038 5624 35050 5627
rect 34756 5596 35050 5624
rect 34756 5584 34762 5596
rect 35038 5593 35050 5596
rect 35084 5593 35096 5627
rect 35038 5587 35096 5593
rect 18506 5556 18512 5568
rect 16408 5528 18512 5556
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 21634 5556 21640 5568
rect 21595 5528 21640 5556
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 23474 5516 23480 5568
rect 23532 5556 23538 5568
rect 23661 5559 23719 5565
rect 23661 5556 23673 5559
rect 23532 5528 23673 5556
rect 23532 5516 23538 5528
rect 23661 5525 23673 5528
rect 23707 5525 23719 5559
rect 23661 5519 23719 5525
rect 24854 5516 24860 5568
rect 24912 5556 24918 5568
rect 26973 5559 27031 5565
rect 26973 5556 26985 5559
rect 24912 5528 26985 5556
rect 24912 5516 24918 5528
rect 26973 5525 26985 5528
rect 27019 5556 27031 5559
rect 28994 5556 29000 5568
rect 27019 5528 29000 5556
rect 27019 5525 27031 5528
rect 26973 5519 27031 5525
rect 28994 5516 29000 5528
rect 29052 5516 29058 5568
rect 30282 5516 30288 5568
rect 30340 5516 30346 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 2498 5352 2504 5364
rect 2459 5324 2504 5352
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 4982 5352 4988 5364
rect 4943 5324 4988 5352
rect 4982 5312 4988 5324
rect 5040 5312 5046 5364
rect 5169 5355 5227 5361
rect 5169 5321 5181 5355
rect 5215 5352 5227 5355
rect 5626 5352 5632 5364
rect 5215 5324 5632 5352
rect 5215 5321 5227 5324
rect 5169 5315 5227 5321
rect 5626 5312 5632 5324
rect 5684 5352 5690 5364
rect 6362 5352 6368 5364
rect 5684 5324 6368 5352
rect 5684 5312 5690 5324
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 6546 5352 6552 5364
rect 6507 5324 6552 5352
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 14274 5352 14280 5364
rect 12483 5324 14280 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 14274 5312 14280 5324
rect 14332 5312 14338 5364
rect 17586 5312 17592 5364
rect 17644 5352 17650 5364
rect 17644 5324 18184 5352
rect 17644 5312 17650 5324
rect 1489 5287 1547 5293
rect 1489 5253 1501 5287
rect 1535 5284 1547 5287
rect 7834 5284 7840 5296
rect 1535 5256 4384 5284
rect 1535 5253 1547 5256
rect 1489 5247 1547 5253
rect 2682 5216 2688 5228
rect 2643 5188 2688 5216
rect 2682 5176 2688 5188
rect 2740 5176 2746 5228
rect 2869 5219 2927 5225
rect 2869 5185 2881 5219
rect 2915 5216 2927 5219
rect 3970 5216 3976 5228
rect 2915 5188 3976 5216
rect 2915 5185 2927 5188
rect 2869 5179 2927 5185
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4356 5225 4384 5256
rect 5721 5251 5779 5257
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4798 5216 4804 5228
rect 4387 5188 4804 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 4982 5176 4988 5228
rect 5040 5216 5046 5228
rect 5350 5216 5356 5228
rect 5040 5188 5356 5216
rect 5040 5176 5046 5188
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5721 5217 5733 5251
rect 5767 5217 5779 5251
rect 6748 5256 7840 5284
rect 5721 5211 5779 5217
rect 6362 5216 6368 5228
rect 3881 5151 3939 5157
rect 3881 5117 3893 5151
rect 3927 5148 3939 5151
rect 4522 5148 4528 5160
rect 3927 5120 4528 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 4706 5108 4712 5160
rect 4764 5148 4770 5160
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 4764 5120 5273 5148
rect 4764 5108 4770 5120
rect 5261 5117 5273 5120
rect 5307 5117 5319 5151
rect 5736 5148 5764 5211
rect 6323 5188 6368 5216
rect 6362 5176 6368 5188
rect 6420 5176 6426 5228
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 6748 5225 6776 5256
rect 7834 5244 7840 5256
rect 7892 5244 7898 5296
rect 18156 5284 18184 5324
rect 18230 5312 18236 5364
rect 18288 5352 18294 5364
rect 19061 5355 19119 5361
rect 19061 5352 19073 5355
rect 18288 5324 19073 5352
rect 18288 5312 18294 5324
rect 19061 5321 19073 5324
rect 19107 5321 19119 5355
rect 20990 5352 20996 5364
rect 19061 5315 19119 5321
rect 19260 5324 20996 5352
rect 18156 5256 18276 5284
rect 6733 5219 6791 5225
rect 6733 5216 6745 5219
rect 6512 5188 6745 5216
rect 6512 5176 6518 5188
rect 6733 5185 6745 5188
rect 6779 5185 6791 5219
rect 6914 5216 6920 5228
rect 6875 5188 6920 5216
rect 6733 5179 6791 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 7653 5219 7711 5225
rect 7653 5216 7665 5219
rect 7524 5188 7665 5216
rect 7524 5176 7530 5188
rect 7653 5185 7665 5188
rect 7699 5216 7711 5219
rect 7699 5188 7972 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 7837 5151 7895 5157
rect 5736 5120 6684 5148
rect 5261 5111 5319 5117
rect 5721 5083 5779 5089
rect 2746 5052 5672 5080
rect 2041 5015 2099 5021
rect 2041 4981 2053 5015
rect 2087 5012 2099 5015
rect 2746 5012 2774 5052
rect 2087 4984 2774 5012
rect 4525 5015 4583 5021
rect 2087 4981 2099 4984
rect 2041 4975 2099 4981
rect 4525 4981 4537 5015
rect 4571 5012 4583 5015
rect 5350 5012 5356 5024
rect 4571 4984 5356 5012
rect 4571 4981 4583 4984
rect 4525 4975 4583 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5644 5012 5672 5052
rect 5721 5049 5733 5083
rect 5767 5080 5779 5083
rect 6270 5080 6276 5092
rect 5767 5052 6276 5080
rect 5767 5049 5779 5052
rect 5721 5043 5779 5049
rect 6270 5040 6276 5052
rect 6328 5040 6334 5092
rect 6454 5012 6460 5024
rect 5644 4984 6460 5012
rect 6454 4972 6460 4984
rect 6512 4972 6518 5024
rect 6656 5012 6684 5120
rect 7837 5117 7849 5151
rect 7883 5117 7895 5151
rect 7944 5148 7972 5188
rect 8018 5176 8024 5228
rect 8076 5216 8082 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8076 5188 8309 5216
rect 8076 5176 8082 5188
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 9677 5219 9735 5225
rect 9677 5185 9689 5219
rect 9723 5216 9735 5219
rect 10962 5216 10968 5228
rect 9723 5188 10968 5216
rect 9723 5185 9735 5188
rect 9677 5179 9735 5185
rect 10962 5176 10968 5188
rect 11020 5176 11026 5228
rect 11514 5176 11520 5228
rect 11572 5216 11578 5228
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11572 5188 11897 5216
rect 11572 5176 11578 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 12066 5176 12072 5228
rect 12124 5216 12130 5228
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 12124 5188 12265 5216
rect 12124 5176 12130 5188
rect 12253 5185 12265 5188
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 14734 5176 14740 5228
rect 14792 5216 14798 5228
rect 15010 5216 15016 5228
rect 14792 5188 15016 5216
rect 14792 5176 14798 5188
rect 15010 5176 15016 5188
rect 15068 5176 15074 5228
rect 17770 5216 17776 5228
rect 17731 5188 17776 5216
rect 17770 5176 17776 5188
rect 17828 5176 17834 5228
rect 17862 5176 17868 5228
rect 17920 5216 17926 5228
rect 17957 5219 18015 5225
rect 17957 5216 17969 5219
rect 17920 5188 17969 5216
rect 17920 5176 17926 5188
rect 17957 5185 17969 5188
rect 18003 5185 18015 5219
rect 17957 5179 18015 5185
rect 18052 5219 18110 5225
rect 18052 5185 18064 5219
rect 18098 5185 18110 5219
rect 18052 5179 18110 5185
rect 18161 5219 18219 5225
rect 18161 5185 18173 5219
rect 18207 5216 18219 5219
rect 18248 5216 18276 5256
rect 19260 5225 19288 5324
rect 20990 5312 20996 5324
rect 21048 5312 21054 5364
rect 23750 5352 23756 5364
rect 23711 5324 23756 5352
rect 23750 5312 23756 5324
rect 23808 5312 23814 5364
rect 25590 5352 25596 5364
rect 25551 5324 25596 5352
rect 25590 5312 25596 5324
rect 25648 5312 25654 5364
rect 34790 5312 34796 5364
rect 34848 5352 34854 5364
rect 35437 5355 35495 5361
rect 35437 5352 35449 5355
rect 34848 5324 35449 5352
rect 34848 5312 34854 5324
rect 35437 5321 35449 5324
rect 35483 5321 35495 5355
rect 35437 5315 35495 5321
rect 19429 5287 19487 5293
rect 19429 5253 19441 5287
rect 19475 5284 19487 5287
rect 19518 5284 19524 5296
rect 19475 5256 19524 5284
rect 19475 5253 19487 5256
rect 19429 5247 19487 5253
rect 19518 5244 19524 5256
rect 19576 5244 19582 5296
rect 24946 5293 24952 5296
rect 24888 5287 24952 5293
rect 24888 5253 24900 5287
rect 24934 5253 24952 5287
rect 24888 5247 24952 5253
rect 24946 5244 24952 5247
rect 25004 5244 25010 5296
rect 27982 5284 27988 5296
rect 27895 5256 27988 5284
rect 27982 5244 27988 5256
rect 28040 5284 28046 5296
rect 28442 5284 28448 5296
rect 28040 5256 28448 5284
rect 28040 5244 28046 5256
rect 28442 5244 28448 5256
rect 28500 5244 28506 5296
rect 28994 5244 29000 5296
rect 29052 5284 29058 5296
rect 29914 5284 29920 5296
rect 29052 5256 29920 5284
rect 29052 5244 29058 5256
rect 29914 5244 29920 5256
rect 29972 5284 29978 5296
rect 33689 5287 33747 5293
rect 33689 5284 33701 5287
rect 29972 5256 33701 5284
rect 29972 5244 29978 5256
rect 33689 5253 33701 5256
rect 33735 5284 33747 5287
rect 34149 5287 34207 5293
rect 34149 5284 34161 5287
rect 33735 5256 34161 5284
rect 33735 5253 33747 5256
rect 33689 5247 33747 5253
rect 34149 5253 34161 5256
rect 34195 5253 34207 5287
rect 34149 5247 34207 5253
rect 18207 5188 18276 5216
rect 19245 5219 19303 5225
rect 18207 5185 18219 5188
rect 18161 5179 18219 5185
rect 19245 5185 19257 5219
rect 19291 5185 19303 5219
rect 25130 5216 25136 5228
rect 25043 5188 25136 5216
rect 19245 5179 19303 5185
rect 8754 5148 8760 5160
rect 7944 5120 8760 5148
rect 7837 5111 7895 5117
rect 7098 5040 7104 5092
rect 7156 5080 7162 5092
rect 7852 5080 7880 5111
rect 8754 5108 8760 5120
rect 8812 5108 8818 5160
rect 11238 5108 11244 5160
rect 11296 5148 11302 5160
rect 11793 5151 11851 5157
rect 11793 5148 11805 5151
rect 11296 5120 11805 5148
rect 11296 5108 11302 5120
rect 11793 5117 11805 5120
rect 11839 5117 11851 5151
rect 12434 5148 12440 5160
rect 11793 5111 11851 5117
rect 12406 5108 12440 5148
rect 12492 5108 12498 5160
rect 17678 5108 17684 5160
rect 17736 5148 17742 5160
rect 18064 5148 18092 5179
rect 25130 5176 25136 5188
rect 25188 5216 25194 5228
rect 26142 5216 26148 5228
rect 25188 5188 26148 5216
rect 25188 5176 25194 5188
rect 26142 5176 26148 5188
rect 26200 5176 26206 5228
rect 28166 5216 28172 5228
rect 28127 5188 28172 5216
rect 28166 5176 28172 5188
rect 28224 5176 28230 5228
rect 20070 5148 20076 5160
rect 17736 5120 18092 5148
rect 18340 5120 20076 5148
rect 17736 5108 17742 5120
rect 8478 5080 8484 5092
rect 7156 5052 7880 5080
rect 8439 5052 8484 5080
rect 7156 5040 7162 5052
rect 6733 5015 6791 5021
rect 6733 5012 6745 5015
rect 6656 4984 6745 5012
rect 6733 4981 6745 4984
rect 6779 5012 6791 5015
rect 7469 5015 7527 5021
rect 7469 5012 7481 5015
rect 6779 4984 7481 5012
rect 6779 4981 6791 4984
rect 6733 4975 6791 4981
rect 7469 4981 7481 4984
rect 7515 4981 7527 5015
rect 7852 5012 7880 5052
rect 8478 5040 8484 5052
rect 8536 5040 8542 5092
rect 10965 5083 11023 5089
rect 10965 5049 10977 5083
rect 11011 5080 11023 5083
rect 12406 5080 12434 5108
rect 11011 5052 12434 5080
rect 13081 5083 13139 5089
rect 11011 5049 11023 5052
rect 10965 5043 11023 5049
rect 13081 5049 13093 5083
rect 13127 5080 13139 5083
rect 15838 5080 15844 5092
rect 13127 5052 15844 5080
rect 13127 5049 13139 5052
rect 13081 5043 13139 5049
rect 15838 5040 15844 5052
rect 15896 5040 15902 5092
rect 7926 5012 7932 5024
rect 7839 4984 7932 5012
rect 7469 4975 7527 4981
rect 7926 4972 7932 4984
rect 7984 5012 7990 5024
rect 8846 5012 8852 5024
rect 7984 4984 8852 5012
rect 7984 4972 7990 4984
rect 8846 4972 8852 4984
rect 8904 4972 8910 5024
rect 10321 5015 10379 5021
rect 10321 4981 10333 5015
rect 10367 5012 10379 5015
rect 11882 5012 11888 5024
rect 10367 4984 11888 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 12250 5012 12256 5024
rect 12211 4984 12256 5012
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 13725 5015 13783 5021
rect 13725 4981 13737 5015
rect 13771 5012 13783 5015
rect 13814 5012 13820 5024
rect 13771 4984 13820 5012
rect 13771 4981 13783 4984
rect 13725 4975 13783 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 14182 5012 14188 5024
rect 14143 4984 14188 5012
rect 14182 4972 14188 4984
rect 14240 4972 14246 5024
rect 14826 5012 14832 5024
rect 14787 4984 14832 5012
rect 14826 4972 14832 4984
rect 14884 4972 14890 5024
rect 15654 4972 15660 5024
rect 15712 5012 15718 5024
rect 15749 5015 15807 5021
rect 15749 5012 15761 5015
rect 15712 4984 15761 5012
rect 15712 4972 15718 4984
rect 15749 4981 15761 4984
rect 15795 4981 15807 5015
rect 15749 4975 15807 4981
rect 17313 5015 17371 5021
rect 17313 4981 17325 5015
rect 17359 5012 17371 5015
rect 17586 5012 17592 5024
rect 17359 4984 17592 5012
rect 17359 4981 17371 4984
rect 17313 4975 17371 4981
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 17862 4972 17868 5024
rect 17920 5012 17926 5024
rect 18340 5012 18368 5120
rect 20070 5108 20076 5120
rect 20128 5108 20134 5160
rect 53742 5108 53748 5160
rect 53800 5148 53806 5160
rect 54389 5151 54447 5157
rect 54389 5148 54401 5151
rect 53800 5120 54401 5148
rect 53800 5108 53806 5120
rect 54389 5117 54401 5120
rect 54435 5117 54447 5151
rect 54389 5111 54447 5117
rect 18417 5083 18475 5089
rect 18417 5049 18429 5083
rect 18463 5080 18475 5083
rect 19334 5080 19340 5092
rect 18463 5052 19340 5080
rect 18463 5049 18475 5052
rect 18417 5043 18475 5049
rect 19334 5040 19340 5052
rect 19392 5040 19398 5092
rect 31570 5080 31576 5092
rect 25148 5052 31576 5080
rect 17920 4984 18368 5012
rect 17920 4972 17926 4984
rect 20070 4972 20076 5024
rect 20128 5012 20134 5024
rect 20165 5015 20223 5021
rect 20165 5012 20177 5015
rect 20128 4984 20177 5012
rect 20128 4972 20134 4984
rect 20165 4981 20177 4984
rect 20211 4981 20223 5015
rect 20165 4975 20223 4981
rect 20898 4972 20904 5024
rect 20956 5012 20962 5024
rect 20993 5015 21051 5021
rect 20993 5012 21005 5015
rect 20956 4984 21005 5012
rect 20956 4972 20962 4984
rect 20993 4981 21005 4984
rect 21039 4981 21051 5015
rect 20993 4975 21051 4981
rect 21726 4972 21732 5024
rect 21784 5012 21790 5024
rect 21821 5015 21879 5021
rect 21821 5012 21833 5015
rect 21784 4984 21833 5012
rect 21784 4972 21790 4984
rect 21821 4981 21833 4984
rect 21867 4981 21879 5015
rect 21821 4975 21879 4981
rect 22554 4972 22560 5024
rect 22612 5012 22618 5024
rect 22649 5015 22707 5021
rect 22649 5012 22661 5015
rect 22612 4984 22661 5012
rect 22612 4972 22618 4984
rect 22649 4981 22661 4984
rect 22695 4981 22707 5015
rect 22649 4975 22707 4981
rect 23014 4972 23020 5024
rect 23072 5012 23078 5024
rect 25148 5012 25176 5052
rect 31570 5040 31576 5052
rect 31628 5040 31634 5092
rect 54110 5040 54116 5092
rect 54168 5080 54174 5092
rect 55033 5083 55091 5089
rect 55033 5080 55045 5083
rect 54168 5052 55045 5080
rect 54168 5040 54174 5052
rect 55033 5049 55045 5052
rect 55079 5049 55091 5083
rect 55033 5043 55091 5049
rect 23072 4984 25176 5012
rect 23072 4972 23078 4984
rect 27338 4972 27344 5024
rect 27396 5012 27402 5024
rect 27801 5015 27859 5021
rect 27801 5012 27813 5015
rect 27396 4984 27813 5012
rect 27396 4972 27402 4984
rect 27801 4981 27813 4984
rect 27847 4981 27859 5015
rect 27801 4975 27859 4981
rect 53650 4972 53656 5024
rect 53708 5012 53714 5024
rect 53745 5015 53803 5021
rect 53745 5012 53757 5015
rect 53708 4984 53757 5012
rect 53708 4972 53714 4984
rect 53745 4981 53757 4984
rect 53791 4981 53803 5015
rect 58158 5012 58164 5024
rect 58119 4984 58164 5012
rect 53745 4975 53803 4981
rect 58158 4972 58164 4984
rect 58216 4972 58222 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 3237 4811 3295 4817
rect 3237 4777 3249 4811
rect 3283 4808 3295 4811
rect 4614 4808 4620 4820
rect 3283 4780 4620 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 5350 4768 5356 4820
rect 5408 4808 5414 4820
rect 5626 4808 5632 4820
rect 5408 4780 5632 4808
rect 5408 4768 5414 4780
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 6914 4808 6920 4820
rect 6875 4780 6920 4808
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7098 4768 7104 4820
rect 7156 4768 7162 4820
rect 7466 4808 7472 4820
rect 7208 4780 7472 4808
rect 2041 4743 2099 4749
rect 2041 4709 2053 4743
rect 2087 4740 2099 4743
rect 6270 4740 6276 4752
rect 2087 4712 6276 4740
rect 2087 4709 2099 4712
rect 2041 4703 2099 4709
rect 6270 4700 6276 4712
rect 6328 4700 6334 4752
rect 6825 4743 6883 4749
rect 6825 4709 6837 4743
rect 6871 4740 6883 4743
rect 7116 4740 7144 4768
rect 6871 4712 7144 4740
rect 6871 4709 6883 4712
rect 6825 4703 6883 4709
rect 5810 4672 5816 4684
rect 2746 4644 5816 4672
rect 1489 4539 1547 4545
rect 1489 4505 1501 4539
rect 1535 4536 1547 4539
rect 2746 4536 2774 4644
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 6641 4675 6699 4681
rect 6641 4641 6653 4675
rect 6687 4672 6699 4675
rect 7098 4672 7104 4684
rect 6687 4644 7104 4672
rect 6687 4641 6699 4644
rect 6641 4635 6699 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 3050 4604 3056 4616
rect 2963 4576 3056 4604
rect 3050 4564 3056 4576
rect 3108 4564 3114 4616
rect 3326 4564 3332 4616
rect 3384 4604 3390 4616
rect 3881 4607 3939 4613
rect 3881 4604 3893 4607
rect 3384 4576 3893 4604
rect 3384 4564 3390 4576
rect 3881 4573 3893 4576
rect 3927 4573 3939 4607
rect 4706 4604 4712 4616
rect 4667 4576 4712 4604
rect 3881 4567 3939 4573
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 5166 4604 5172 4616
rect 4939 4576 5172 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 6181 4607 6239 4613
rect 6181 4573 6193 4607
rect 6227 4604 6239 4607
rect 6730 4604 6736 4616
rect 6227 4576 6736 4604
rect 6227 4573 6239 4576
rect 6181 4567 6239 4573
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7208 4604 7236 4780
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7926 4808 7932 4820
rect 7887 4780 7932 4808
rect 7926 4768 7932 4780
rect 7984 4768 7990 4820
rect 8297 4811 8355 4817
rect 8297 4777 8309 4811
rect 8343 4808 8355 4811
rect 8386 4808 8392 4820
rect 8343 4780 8392 4808
rect 8343 4777 8355 4780
rect 8297 4771 8355 4777
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 8938 4808 8944 4820
rect 8899 4780 8944 4808
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 9401 4811 9459 4817
rect 9401 4808 9413 4811
rect 9364 4780 9413 4808
rect 9364 4768 9370 4780
rect 9401 4777 9413 4780
rect 9447 4777 9459 4811
rect 9401 4771 9459 4777
rect 10321 4811 10379 4817
rect 10321 4777 10333 4811
rect 10367 4808 10379 4811
rect 10870 4808 10876 4820
rect 10367 4780 10876 4808
rect 10367 4777 10379 4780
rect 10321 4771 10379 4777
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 11422 4808 11428 4820
rect 10980 4780 11428 4808
rect 7282 4700 7288 4752
rect 7340 4740 7346 4752
rect 10505 4743 10563 4749
rect 10505 4740 10517 4743
rect 7340 4712 10517 4740
rect 7340 4700 7346 4712
rect 10505 4709 10517 4712
rect 10551 4740 10563 4743
rect 10980 4740 11008 4780
rect 11422 4768 11428 4780
rect 11480 4808 11486 4820
rect 11701 4811 11759 4817
rect 11701 4808 11713 4811
rect 11480 4780 11713 4808
rect 11480 4768 11486 4780
rect 11701 4777 11713 4780
rect 11747 4777 11759 4811
rect 11701 4771 11759 4777
rect 10551 4712 11008 4740
rect 10551 4709 10563 4712
rect 10505 4703 10563 4709
rect 11514 4700 11520 4752
rect 11572 4740 11578 4752
rect 11609 4743 11667 4749
rect 11609 4740 11621 4743
rect 11572 4712 11621 4740
rect 11572 4700 11578 4712
rect 11609 4709 11621 4712
rect 11655 4709 11667 4743
rect 11716 4740 11744 4771
rect 11790 4768 11796 4820
rect 11848 4808 11854 4820
rect 11885 4811 11943 4817
rect 11885 4808 11897 4811
rect 11848 4780 11897 4808
rect 11848 4768 11854 4780
rect 11885 4777 11897 4780
rect 11931 4808 11943 4811
rect 21082 4808 21088 4820
rect 11931 4780 21088 4808
rect 11931 4777 11943 4780
rect 11885 4771 11943 4777
rect 21082 4768 21088 4780
rect 21140 4768 21146 4820
rect 22465 4811 22523 4817
rect 22465 4777 22477 4811
rect 22511 4808 22523 4811
rect 22922 4808 22928 4820
rect 22511 4780 22928 4808
rect 22511 4777 22523 4780
rect 22465 4771 22523 4777
rect 22922 4768 22928 4780
rect 22980 4768 22986 4820
rect 23198 4768 23204 4820
rect 23256 4808 23262 4820
rect 42058 4808 42064 4820
rect 23256 4780 42064 4808
rect 23256 4768 23262 4780
rect 42058 4768 42064 4780
rect 42116 4768 42122 4820
rect 12250 4740 12256 4752
rect 11716 4712 12256 4740
rect 11609 4703 11667 4709
rect 12250 4700 12256 4712
rect 12308 4700 12314 4752
rect 17405 4743 17463 4749
rect 17405 4709 17417 4743
rect 17451 4740 17463 4743
rect 18690 4740 18696 4752
rect 17451 4712 18696 4740
rect 17451 4709 17463 4712
rect 17405 4703 17463 4709
rect 18690 4700 18696 4712
rect 18748 4700 18754 4752
rect 26418 4740 26424 4752
rect 26379 4712 26424 4740
rect 26418 4700 26424 4712
rect 26476 4700 26482 4752
rect 52178 4700 52184 4752
rect 52236 4740 52242 4752
rect 52825 4743 52883 4749
rect 52825 4740 52837 4743
rect 52236 4712 52837 4740
rect 52236 4700 52242 4712
rect 52825 4709 52837 4712
rect 52871 4709 52883 4743
rect 52825 4703 52883 4709
rect 53926 4700 53932 4752
rect 53984 4740 53990 4752
rect 55309 4743 55367 4749
rect 55309 4740 55321 4743
rect 53984 4712 55321 4740
rect 53984 4700 53990 4712
rect 55309 4709 55321 4712
rect 55355 4709 55367 4743
rect 55309 4703 55367 4709
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8128 4644 9045 4672
rect 7466 4604 7472 4616
rect 6963 4576 7236 4604
rect 7427 4576 7472 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7466 4564 7472 4576
rect 7524 4564 7530 4616
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 7616 4576 7661 4604
rect 7616 4564 7622 4576
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 7995 4607 8053 4613
rect 7995 4604 8007 4607
rect 7892 4576 8007 4604
rect 7892 4564 7898 4576
rect 7995 4573 8007 4576
rect 8041 4604 8053 4607
rect 8128 4604 8156 4644
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9033 4635 9091 4641
rect 9140 4644 9352 4672
rect 8041 4576 8156 4604
rect 8041 4573 8053 4576
rect 7995 4567 8053 4573
rect 8846 4564 8852 4616
rect 8904 4604 8910 4616
rect 8941 4607 8999 4613
rect 8941 4604 8953 4607
rect 8904 4576 8953 4604
rect 8904 4564 8910 4576
rect 8941 4573 8953 4576
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 1535 4508 2774 4536
rect 3068 4536 3096 4564
rect 3970 4536 3976 4548
rect 3068 4508 3976 4536
rect 1535 4505 1547 4508
rect 1489 4499 1547 4505
rect 3970 4496 3976 4508
rect 4028 4496 4034 4548
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 9140 4536 9168 4644
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 7156 4508 9168 4536
rect 7156 4496 7162 4508
rect 2593 4471 2651 4477
rect 2593 4437 2605 4471
rect 2639 4468 2651 4471
rect 3234 4468 3240 4480
rect 2639 4440 3240 4468
rect 2639 4437 2651 4440
rect 2593 4431 2651 4437
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 4065 4471 4123 4477
rect 4065 4437 4077 4471
rect 4111 4468 4123 4471
rect 4338 4468 4344 4480
rect 4111 4440 4344 4468
rect 4111 4437 4123 4440
rect 4065 4431 4123 4437
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 4522 4468 4528 4480
rect 4483 4440 4528 4468
rect 4522 4428 4528 4440
rect 4580 4428 4586 4480
rect 5445 4471 5503 4477
rect 5445 4437 5457 4471
rect 5491 4468 5503 4471
rect 5902 4468 5908 4480
rect 5491 4440 5908 4468
rect 5491 4437 5503 4440
rect 5445 4431 5503 4437
rect 5902 4428 5908 4440
rect 5960 4428 5966 4480
rect 5997 4471 6055 4477
rect 5997 4437 6009 4471
rect 6043 4468 6055 4471
rect 6546 4468 6552 4480
rect 6043 4440 6552 4468
rect 6043 4437 6055 4440
rect 5997 4431 6055 4437
rect 6546 4428 6552 4440
rect 6604 4428 6610 4480
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 9232 4468 9260 4567
rect 9324 4536 9352 4644
rect 9398 4632 9404 4684
rect 9456 4672 9462 4684
rect 10413 4675 10471 4681
rect 10413 4672 10425 4675
rect 9456 4644 10425 4672
rect 9456 4632 9462 4644
rect 10413 4641 10425 4644
rect 10459 4672 10471 4675
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 10459 4644 11805 4672
rect 10459 4641 10471 4644
rect 10413 4635 10471 4641
rect 11793 4641 11805 4644
rect 11839 4672 11851 4675
rect 12066 4672 12072 4684
rect 11839 4644 12072 4672
rect 11839 4641 11851 4644
rect 11793 4635 11851 4641
rect 12066 4632 12072 4644
rect 12124 4632 12130 4684
rect 12897 4675 12955 4681
rect 12897 4641 12909 4675
rect 12943 4672 12955 4675
rect 13538 4672 13544 4684
rect 12943 4644 13544 4672
rect 12943 4641 12955 4644
rect 12897 4635 12955 4641
rect 13538 4632 13544 4644
rect 13596 4632 13602 4684
rect 16117 4675 16175 4681
rect 16117 4641 16129 4675
rect 16163 4672 16175 4675
rect 17034 4672 17040 4684
rect 16163 4644 17040 4672
rect 16163 4641 16175 4644
rect 16117 4635 16175 4641
rect 17034 4632 17040 4644
rect 17092 4632 17098 4684
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4672 18107 4675
rect 18966 4672 18972 4684
rect 18095 4644 18972 4672
rect 18095 4641 18107 4644
rect 18049 4635 18107 4641
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 23845 4675 23903 4681
rect 23845 4641 23857 4675
rect 23891 4672 23903 4675
rect 25130 4672 25136 4684
rect 23891 4644 25136 4672
rect 23891 4641 23903 4644
rect 23845 4635 23903 4641
rect 25130 4632 25136 4644
rect 25188 4632 25194 4684
rect 10634 4607 10692 4613
rect 10634 4573 10646 4607
rect 10680 4604 10692 4607
rect 11238 4604 11244 4616
rect 10680 4576 11244 4604
rect 10680 4573 10692 4576
rect 10634 4567 10692 4573
rect 11238 4564 11244 4576
rect 11296 4564 11302 4616
rect 13354 4604 13360 4616
rect 13267 4576 13360 4604
rect 13354 4564 13360 4576
rect 13412 4604 13418 4616
rect 14274 4604 14280 4616
rect 13412 4576 14280 4604
rect 13412 4564 13418 4576
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14829 4607 14887 4613
rect 14829 4573 14841 4607
rect 14875 4604 14887 4607
rect 15378 4604 15384 4616
rect 14875 4576 15384 4604
rect 14875 4573 14887 4576
rect 14829 4567 14887 4573
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 15473 4607 15531 4613
rect 15473 4573 15485 4607
rect 15519 4604 15531 4607
rect 15930 4604 15936 4616
rect 15519 4576 15936 4604
rect 15519 4573 15531 4576
rect 15473 4567 15531 4573
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 16761 4607 16819 4613
rect 16761 4573 16773 4607
rect 16807 4573 16819 4607
rect 16761 4567 16819 4573
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4604 18751 4607
rect 19242 4604 19248 4616
rect 18739 4576 19248 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 10781 4539 10839 4545
rect 10781 4536 10793 4539
rect 9324 4508 10793 4536
rect 10781 4505 10793 4508
rect 10827 4536 10839 4539
rect 11514 4536 11520 4548
rect 10827 4508 11520 4536
rect 10827 4505 10839 4508
rect 10781 4499 10839 4505
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 16776 4536 16804 4567
rect 19242 4564 19248 4576
rect 19300 4564 19306 4616
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19392 4576 19441 4604
rect 19392 4564 19398 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 20073 4607 20131 4613
rect 20073 4573 20085 4607
rect 20119 4604 20131 4607
rect 20622 4604 20628 4616
rect 20119 4576 20628 4604
rect 20119 4573 20131 4576
rect 20073 4567 20131 4573
rect 20622 4564 20628 4576
rect 20680 4564 20686 4616
rect 20717 4607 20775 4613
rect 20717 4573 20729 4607
rect 20763 4604 20775 4607
rect 21082 4604 21088 4616
rect 20763 4576 21088 4604
rect 20763 4573 20775 4576
rect 20717 4567 20775 4573
rect 21082 4564 21088 4576
rect 21140 4564 21146 4616
rect 21361 4607 21419 4613
rect 21361 4573 21373 4607
rect 21407 4604 21419 4607
rect 21910 4604 21916 4616
rect 21407 4576 21916 4604
rect 21407 4573 21419 4576
rect 21361 4567 21419 4573
rect 21910 4564 21916 4576
rect 21968 4564 21974 4616
rect 22005 4607 22063 4613
rect 22005 4573 22017 4607
rect 22051 4604 22063 4607
rect 22186 4604 22192 4616
rect 22051 4576 22192 4604
rect 22051 4573 22063 4576
rect 22005 4567 22063 4573
rect 22186 4564 22192 4576
rect 22244 4564 22250 4616
rect 23566 4564 23572 4616
rect 23624 4613 23630 4616
rect 23624 4604 23636 4613
rect 24949 4607 25007 4613
rect 24949 4604 24961 4607
rect 23624 4576 23669 4604
rect 23860 4576 24961 4604
rect 23624 4567 23636 4576
rect 23624 4564 23630 4567
rect 18046 4536 18052 4548
rect 16776 4508 18052 4536
rect 18046 4496 18052 4508
rect 18104 4496 18110 4548
rect 23290 4496 23296 4548
rect 23348 4536 23354 4548
rect 23750 4536 23756 4548
rect 23348 4508 23756 4536
rect 23348 4496 23354 4508
rect 23750 4496 23756 4508
rect 23808 4496 23814 4548
rect 8260 4440 9260 4468
rect 13541 4471 13599 4477
rect 8260 4428 8266 4440
rect 13541 4437 13553 4471
rect 13587 4468 13599 4471
rect 13906 4468 13912 4480
rect 13587 4440 13912 4468
rect 13587 4437 13599 4440
rect 13541 4431 13599 4437
rect 13906 4428 13912 4440
rect 13964 4428 13970 4480
rect 14185 4471 14243 4477
rect 14185 4437 14197 4471
rect 14231 4468 14243 4471
rect 17862 4468 17868 4480
rect 14231 4440 17868 4468
rect 14231 4437 14243 4440
rect 14185 4431 14243 4437
rect 17862 4428 17868 4440
rect 17920 4428 17926 4480
rect 22370 4428 22376 4480
rect 22428 4468 22434 4480
rect 23860 4468 23888 4576
rect 24949 4573 24961 4576
rect 24995 4573 25007 4607
rect 26436 4604 26464 4700
rect 27062 4632 27068 4684
rect 27120 4672 27126 4684
rect 31481 4675 31539 4681
rect 31481 4672 31493 4675
rect 27120 4644 27292 4672
rect 27120 4632 27126 4644
rect 27264 4613 27292 4644
rect 30208 4644 31493 4672
rect 27157 4607 27215 4613
rect 27157 4604 27169 4607
rect 26436 4576 27169 4604
rect 24949 4567 25007 4573
rect 27157 4573 27169 4576
rect 27203 4573 27215 4607
rect 27157 4567 27215 4573
rect 27249 4607 27307 4613
rect 27249 4573 27261 4607
rect 27295 4573 27307 4607
rect 27249 4567 27307 4573
rect 27338 4564 27344 4616
rect 27396 4604 27402 4616
rect 27396 4576 27441 4604
rect 27396 4564 27402 4576
rect 27522 4564 27528 4616
rect 27580 4604 27586 4616
rect 30208 4613 30236 4644
rect 31481 4641 31493 4644
rect 31527 4641 31539 4675
rect 31481 4635 31539 4641
rect 53190 4632 53196 4684
rect 53248 4672 53254 4684
rect 54113 4675 54171 4681
rect 54113 4672 54125 4675
rect 53248 4644 54125 4672
rect 53248 4632 53254 4644
rect 54113 4641 54125 4644
rect 54159 4641 54171 4675
rect 54113 4635 54171 4641
rect 54294 4632 54300 4684
rect 54352 4672 54358 4684
rect 55953 4675 56011 4681
rect 55953 4672 55965 4675
rect 54352 4644 55965 4672
rect 54352 4632 54358 4644
rect 55953 4641 55965 4644
rect 55999 4641 56011 4675
rect 55953 4635 56011 4641
rect 30009 4607 30067 4613
rect 30009 4604 30021 4607
rect 27580 4576 30021 4604
rect 27580 4564 27586 4576
rect 30009 4573 30021 4576
rect 30055 4573 30067 4607
rect 30009 4567 30067 4573
rect 30193 4607 30251 4613
rect 30193 4573 30205 4607
rect 30239 4573 30251 4607
rect 30193 4567 30251 4573
rect 30282 4564 30288 4616
rect 30340 4604 30346 4616
rect 30423 4607 30481 4613
rect 30340 4576 30385 4604
rect 30340 4564 30346 4576
rect 30423 4573 30435 4607
rect 30469 4604 30481 4607
rect 30834 4604 30840 4616
rect 30469 4576 30840 4604
rect 30469 4573 30481 4576
rect 30423 4567 30481 4573
rect 30834 4564 30840 4576
rect 30892 4564 30898 4616
rect 31110 4604 31116 4616
rect 31071 4576 31116 4604
rect 31110 4564 31116 4576
rect 31168 4564 31174 4616
rect 31297 4607 31355 4613
rect 31297 4573 31309 4607
rect 31343 4604 31355 4607
rect 32398 4604 32404 4616
rect 31343 4576 32404 4604
rect 31343 4573 31355 4576
rect 31297 4567 31355 4573
rect 32398 4564 32404 4576
rect 32456 4564 32462 4616
rect 52086 4564 52092 4616
rect 52144 4604 52150 4616
rect 52181 4607 52239 4613
rect 52181 4604 52193 4607
rect 52144 4576 52193 4604
rect 52144 4564 52150 4576
rect 52181 4573 52193 4576
rect 52227 4573 52239 4607
rect 52181 4567 52239 4573
rect 52638 4564 52644 4616
rect 52696 4604 52702 4616
rect 53469 4607 53527 4613
rect 53469 4604 53481 4607
rect 52696 4576 53481 4604
rect 52696 4564 52702 4576
rect 53469 4573 53481 4576
rect 53515 4573 53527 4607
rect 53469 4567 53527 4573
rect 23934 4496 23940 4548
rect 23992 4536 23998 4548
rect 25501 4539 25559 4545
rect 25501 4536 25513 4539
rect 23992 4508 25513 4536
rect 23992 4496 23998 4508
rect 25501 4505 25513 4508
rect 25547 4505 25559 4539
rect 25501 4499 25559 4505
rect 24394 4468 24400 4480
rect 22428 4440 23888 4468
rect 24355 4440 24400 4468
rect 22428 4428 22434 4440
rect 24394 4428 24400 4440
rect 24452 4428 24458 4480
rect 26878 4468 26884 4480
rect 26839 4440 26884 4468
rect 26878 4428 26884 4440
rect 26936 4428 26942 4480
rect 30650 4468 30656 4480
rect 30611 4440 30656 4468
rect 30650 4428 30656 4440
rect 30708 4428 30714 4480
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 4706 4224 4712 4276
rect 4764 4264 4770 4276
rect 6086 4264 6092 4276
rect 4764 4236 6092 4264
rect 4764 4224 4770 4236
rect 6086 4224 6092 4236
rect 6144 4264 6150 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6144 4236 6561 4264
rect 6144 4224 6150 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 7926 4224 7932 4276
rect 7984 4224 7990 4276
rect 8754 4264 8760 4276
rect 8715 4236 8760 4264
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 8938 4224 8944 4276
rect 8996 4264 9002 4276
rect 9766 4264 9772 4276
rect 8996 4236 9168 4264
rect 9727 4236 9772 4264
rect 8996 4224 9002 4236
rect 4890 4196 4896 4208
rect 4851 4168 4896 4196
rect 4890 4156 4896 4168
rect 4948 4196 4954 4208
rect 5350 4196 5356 4208
rect 4948 4168 5356 4196
rect 4948 4156 4954 4168
rect 5350 4156 5356 4168
rect 5408 4156 5414 4208
rect 6362 4196 6368 4208
rect 6323 4168 6368 4196
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 7653 4199 7711 4205
rect 7653 4165 7665 4199
rect 7699 4196 7711 4199
rect 7944 4196 7972 4224
rect 7699 4168 7972 4196
rect 7699 4165 7711 4168
rect 7653 4159 7711 4165
rect 2317 4131 2375 4137
rect 2317 4097 2329 4131
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 2332 4060 2360 4091
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 2832 4100 2877 4128
rect 2832 4088 2838 4100
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3421 4131 3479 4137
rect 3421 4128 3433 4131
rect 3200 4100 3433 4128
rect 3200 4088 3206 4100
rect 3421 4097 3433 4100
rect 3467 4097 3479 4131
rect 4062 4128 4068 4140
rect 4023 4100 4068 4128
rect 3421 4091 3479 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 5810 4128 5816 4140
rect 4396 4100 4936 4128
rect 5723 4100 5816 4128
rect 4396 4088 4402 4100
rect 4522 4060 4528 4072
rect 2332 4032 4528 4060
rect 4522 4020 4528 4032
rect 4580 4020 4586 4072
rect 4908 4060 4936 4100
rect 5810 4088 5816 4100
rect 5868 4128 5874 4140
rect 7282 4128 7288 4140
rect 5868 4100 7288 4128
rect 5868 4088 5874 4100
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 7524 4100 8125 4128
rect 7524 4088 7530 4100
rect 8113 4097 8125 4100
rect 8159 4128 8171 4131
rect 8202 4128 8208 4140
rect 8159 4100 8208 4128
rect 8159 4097 8171 4100
rect 8113 4091 8171 4097
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8846 4088 8852 4140
rect 8904 4128 8910 4140
rect 9140 4137 9168 4236
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 16390 4224 16396 4276
rect 16448 4264 16454 4276
rect 16448 4236 22094 4264
rect 16448 4224 16454 4236
rect 22066 4196 22094 4236
rect 22462 4224 22468 4276
rect 22520 4264 22526 4276
rect 25866 4264 25872 4276
rect 22520 4236 25872 4264
rect 22520 4224 22526 4236
rect 25866 4224 25872 4236
rect 25924 4224 25930 4276
rect 29914 4264 29920 4276
rect 29827 4236 29920 4264
rect 29914 4224 29920 4236
rect 29972 4264 29978 4276
rect 30834 4264 30840 4276
rect 29972 4236 30840 4264
rect 29972 4224 29978 4236
rect 30834 4224 30840 4236
rect 30892 4224 30898 4276
rect 26418 4196 26424 4208
rect 16684 4168 17080 4196
rect 22066 4168 26424 4196
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8904 4100 8953 4128
rect 8904 4088 8910 4100
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 9125 4131 9183 4137
rect 9125 4097 9137 4131
rect 9171 4097 9183 4131
rect 9125 4091 9183 4097
rect 4908 4032 6583 4060
rect 2961 3995 3019 4001
rect 2961 3961 2973 3995
rect 3007 3992 3019 3995
rect 5902 3992 5908 4004
rect 3007 3964 5908 3992
rect 3007 3961 3019 3964
rect 2961 3955 3019 3961
rect 5902 3952 5908 3964
rect 5960 3952 5966 4004
rect 1670 3924 1676 3936
rect 1631 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 2130 3924 2136 3936
rect 2091 3896 2136 3924
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 3605 3927 3663 3933
rect 3605 3893 3617 3927
rect 3651 3924 3663 3927
rect 3786 3924 3792 3936
rect 3651 3896 3792 3924
rect 3651 3893 3663 3896
rect 3605 3887 3663 3893
rect 3786 3884 3792 3896
rect 3844 3884 3850 3936
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 4890 3924 4896 3936
rect 4295 3896 4896 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 4985 3927 5043 3933
rect 4985 3893 4997 3927
rect 5031 3924 5043 3927
rect 5442 3924 5448 3936
rect 5031 3896 5448 3924
rect 5031 3893 5043 3896
rect 4985 3887 5043 3893
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 5629 3927 5687 3933
rect 5629 3893 5641 3927
rect 5675 3924 5687 3927
rect 5994 3924 6000 3936
rect 5675 3896 6000 3924
rect 5675 3893 5687 3896
rect 5629 3887 5687 3893
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 6555 3933 6583 4032
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7892 4032 7941 4060
rect 7892 4020 7898 4032
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 8018 3952 8024 4004
rect 8076 3992 8082 4004
rect 8220 3992 8248 4088
rect 8754 4020 8760 4072
rect 8812 4060 8818 4072
rect 9140 4060 9168 4091
rect 9214 4088 9220 4140
rect 9272 4128 9278 4140
rect 9585 4131 9643 4137
rect 9585 4128 9597 4131
rect 9272 4100 9597 4128
rect 9272 4088 9278 4100
rect 9585 4097 9597 4100
rect 9631 4097 9643 4131
rect 10594 4128 10600 4140
rect 10555 4100 10600 4128
rect 9585 4091 9643 4097
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 11514 4128 11520 4140
rect 11475 4100 11520 4128
rect 11514 4088 11520 4100
rect 11572 4088 11578 4140
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 14090 4128 14096 4140
rect 12768 4100 14096 4128
rect 12768 4088 12774 4100
rect 14090 4088 14096 4100
rect 14148 4088 14154 4140
rect 16684 4137 16712 4168
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4097 16727 4131
rect 16936 4131 16994 4137
rect 16936 4128 16948 4131
rect 16669 4091 16727 4097
rect 16776 4100 16948 4128
rect 12066 4060 12072 4072
rect 8812 4032 9168 4060
rect 12027 4032 12072 4060
rect 8812 4020 8818 4032
rect 12066 4020 12072 4032
rect 12124 4020 12130 4072
rect 12345 4063 12403 4069
rect 12345 4029 12357 4063
rect 12391 4060 12403 4063
rect 13078 4060 13084 4072
rect 12391 4032 13084 4060
rect 12391 4029 12403 4032
rect 12345 4023 12403 4029
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 14829 4063 14887 4069
rect 14829 4029 14841 4063
rect 14875 4060 14887 4063
rect 16022 4060 16028 4072
rect 14875 4032 16028 4060
rect 14875 4029 14887 4032
rect 14829 4023 14887 4029
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 16114 4020 16120 4072
rect 16172 4060 16178 4072
rect 16776 4060 16804 4100
rect 16936 4097 16948 4100
rect 16982 4097 16994 4131
rect 17052 4128 17080 4168
rect 26418 4156 26424 4168
rect 26476 4156 26482 4208
rect 19058 4128 19064 4140
rect 17052 4100 19064 4128
rect 16936 4091 16994 4097
rect 19058 4088 19064 4100
rect 19116 4128 19122 4140
rect 19429 4131 19487 4137
rect 19429 4128 19441 4131
rect 19116 4100 19441 4128
rect 19116 4088 19122 4100
rect 19429 4097 19441 4100
rect 19475 4097 19487 4131
rect 19429 4091 19487 4097
rect 19518 4088 19524 4140
rect 19576 4128 19582 4140
rect 19685 4131 19743 4137
rect 19685 4128 19697 4131
rect 19576 4100 19697 4128
rect 19576 4088 19582 4100
rect 19685 4097 19697 4100
rect 19731 4097 19743 4131
rect 19685 4091 19743 4097
rect 20990 4088 20996 4140
rect 21048 4088 21054 4140
rect 34790 4088 34796 4140
rect 34848 4128 34854 4140
rect 34885 4131 34943 4137
rect 34885 4128 34897 4131
rect 34848 4100 34897 4128
rect 34848 4088 34854 4100
rect 34885 4097 34897 4100
rect 34931 4097 34943 4131
rect 34885 4091 34943 4097
rect 35152 4131 35210 4137
rect 35152 4097 35164 4131
rect 35198 4128 35210 4131
rect 35434 4128 35440 4140
rect 35198 4100 35440 4128
rect 35198 4097 35210 4100
rect 35152 4091 35210 4097
rect 35434 4088 35440 4100
rect 35492 4088 35498 4140
rect 53006 4088 53012 4140
rect 53064 4128 53070 4140
rect 54665 4131 54723 4137
rect 54665 4128 54677 4131
rect 53064 4100 54677 4128
rect 53064 4088 53070 4100
rect 54665 4097 54677 4100
rect 54711 4097 54723 4131
rect 54665 4091 54723 4097
rect 16172 4032 16804 4060
rect 21008 4060 21036 4088
rect 26326 4060 26332 4072
rect 21008 4032 26332 4060
rect 16172 4020 16178 4032
rect 8076 3964 8984 3992
rect 8076 3952 8082 3964
rect 6549 3927 6607 3933
rect 6549 3893 6561 3927
rect 6595 3893 6607 3927
rect 6730 3924 6736 3936
rect 6691 3896 6736 3924
rect 6549 3887 6607 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 7558 3884 7564 3936
rect 7616 3924 7622 3936
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 7616 3896 7757 3924
rect 7616 3884 7622 3896
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 8294 3924 8300 3936
rect 8255 3896 8300 3924
rect 7745 3887 7803 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8956 3933 8984 3964
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 10413 3995 10471 4001
rect 10413 3992 10425 3995
rect 9272 3964 10425 3992
rect 9272 3952 9278 3964
rect 10413 3961 10425 3964
rect 10459 3961 10471 3995
rect 10413 3955 10471 3961
rect 11422 3952 11428 4004
rect 11480 3992 11486 4004
rect 11977 3995 12035 4001
rect 11977 3992 11989 3995
rect 11480 3964 11989 3992
rect 11480 3952 11486 3964
rect 11977 3961 11989 3964
rect 12023 3961 12035 3995
rect 11977 3955 12035 3961
rect 12618 3952 12624 4004
rect 12676 3992 12682 4004
rect 13630 3992 13636 4004
rect 12676 3964 13636 3992
rect 12676 3952 12682 3964
rect 13630 3952 13636 3964
rect 13688 3952 13694 4004
rect 14185 3995 14243 4001
rect 14185 3961 14197 3995
rect 14231 3992 14243 3995
rect 15194 3992 15200 4004
rect 14231 3964 15200 3992
rect 14231 3961 14243 3964
rect 14185 3955 14243 3961
rect 15194 3952 15200 3964
rect 15252 3952 15258 4004
rect 15473 3995 15531 4001
rect 15473 3961 15485 3995
rect 15519 3992 15531 3995
rect 16666 3992 16672 4004
rect 15519 3964 16672 3992
rect 15519 3961 15531 3964
rect 15473 3955 15531 3961
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 18414 3992 18420 4004
rect 17972 3964 18420 3992
rect 8941 3927 8999 3933
rect 8941 3893 8953 3927
rect 8987 3893 8999 3927
rect 8941 3887 8999 3893
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 11885 3927 11943 3933
rect 11885 3924 11897 3927
rect 11296 3896 11897 3924
rect 11296 3884 11302 3896
rect 11885 3893 11897 3896
rect 11931 3893 11943 3927
rect 11885 3887 11943 3893
rect 13541 3927 13599 3933
rect 13541 3893 13553 3927
rect 13587 3924 13599 3927
rect 14642 3924 14648 3936
rect 13587 3896 14648 3924
rect 13587 3893 13599 3896
rect 13541 3887 13599 3893
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 16117 3927 16175 3933
rect 16117 3893 16129 3927
rect 16163 3924 16175 3927
rect 17972 3924 18000 3964
rect 18414 3952 18420 3964
rect 18472 3952 18478 4004
rect 20809 3995 20867 4001
rect 20809 3961 20821 3995
rect 20855 3992 20867 3995
rect 21008 3992 21036 4032
rect 26326 4020 26332 4032
rect 26384 4020 26390 4072
rect 51810 4020 51816 4072
rect 51868 4060 51874 4072
rect 52733 4063 52791 4069
rect 52733 4060 52745 4063
rect 51868 4032 52745 4060
rect 51868 4020 51874 4032
rect 52733 4029 52745 4032
rect 52779 4029 52791 4063
rect 52733 4023 52791 4029
rect 54018 4020 54024 4072
rect 54076 4060 54082 4072
rect 55953 4063 56011 4069
rect 55953 4060 55965 4063
rect 54076 4032 55965 4060
rect 54076 4020 54082 4032
rect 55953 4029 55965 4032
rect 55999 4029 56011 4063
rect 55953 4023 56011 4029
rect 20855 3964 21036 3992
rect 20855 3961 20867 3964
rect 20809 3955 20867 3961
rect 21542 3952 21548 4004
rect 21600 3992 21606 4004
rect 26053 3995 26111 4001
rect 26053 3992 26065 3995
rect 21600 3964 26065 3992
rect 21600 3952 21606 3964
rect 26053 3961 26065 3964
rect 26099 3961 26111 3995
rect 26053 3955 26111 3961
rect 52822 3952 52828 4004
rect 52880 3992 52886 4004
rect 52880 3964 54064 3992
rect 52880 3952 52886 3964
rect 16163 3896 18000 3924
rect 18049 3927 18107 3933
rect 16163 3893 16175 3896
rect 16117 3887 16175 3893
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 18506 3924 18512 3936
rect 18095 3896 18512 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 18506 3884 18512 3896
rect 18564 3884 18570 3936
rect 18874 3884 18880 3936
rect 18932 3924 18938 3936
rect 18969 3927 19027 3933
rect 18969 3924 18981 3927
rect 18932 3896 18981 3924
rect 18932 3884 18938 3896
rect 18969 3893 18981 3896
rect 19015 3893 19027 3927
rect 18969 3887 19027 3893
rect 19426 3884 19432 3936
rect 19484 3924 19490 3936
rect 20346 3924 20352 3936
rect 19484 3896 20352 3924
rect 19484 3884 19490 3896
rect 20346 3884 20352 3896
rect 20404 3884 20410 3936
rect 22373 3927 22431 3933
rect 22373 3893 22385 3927
rect 22419 3924 22431 3927
rect 22922 3924 22928 3936
rect 22419 3896 22928 3924
rect 22419 3893 22431 3896
rect 22373 3887 22431 3893
rect 22922 3884 22928 3896
rect 22980 3884 22986 3936
rect 23017 3927 23075 3933
rect 23017 3893 23029 3927
rect 23063 3924 23075 3927
rect 23106 3924 23112 3936
rect 23063 3896 23112 3924
rect 23063 3893 23075 3896
rect 23017 3887 23075 3893
rect 23106 3884 23112 3896
rect 23164 3884 23170 3936
rect 23382 3884 23388 3936
rect 23440 3924 23446 3936
rect 23477 3927 23535 3933
rect 23477 3924 23489 3927
rect 23440 3896 23489 3924
rect 23440 3884 23446 3896
rect 23477 3893 23489 3896
rect 23523 3893 23535 3927
rect 23477 3887 23535 3893
rect 24210 3884 24216 3936
rect 24268 3924 24274 3936
rect 24305 3927 24363 3933
rect 24305 3924 24317 3927
rect 24268 3896 24317 3924
rect 24268 3884 24274 3896
rect 24305 3893 24317 3896
rect 24351 3893 24363 3927
rect 24305 3887 24363 3893
rect 25314 3884 25320 3936
rect 25372 3924 25378 3936
rect 25409 3927 25467 3933
rect 25409 3924 25421 3927
rect 25372 3896 25421 3924
rect 25372 3884 25378 3896
rect 25409 3893 25421 3896
rect 25455 3893 25467 3927
rect 25409 3887 25467 3893
rect 35618 3884 35624 3936
rect 35676 3924 35682 3936
rect 36265 3927 36323 3933
rect 36265 3924 36277 3927
rect 35676 3896 36277 3924
rect 35676 3884 35682 3896
rect 36265 3893 36277 3896
rect 36311 3893 36323 3927
rect 36265 3887 36323 3893
rect 51074 3884 51080 3936
rect 51132 3924 51138 3936
rect 51169 3927 51227 3933
rect 51169 3924 51181 3927
rect 51132 3896 51181 3924
rect 51132 3884 51138 3896
rect 51169 3893 51181 3896
rect 51215 3893 51227 3927
rect 51169 3887 51227 3893
rect 51350 3884 51356 3936
rect 51408 3924 51414 3936
rect 51813 3927 51871 3933
rect 51813 3924 51825 3927
rect 51408 3896 51825 3924
rect 51408 3884 51414 3896
rect 51813 3893 51825 3896
rect 51859 3893 51871 3927
rect 51813 3887 51871 3893
rect 52454 3884 52460 3936
rect 52512 3924 52518 3936
rect 54036 3933 54064 3964
rect 53377 3927 53435 3933
rect 53377 3924 53389 3927
rect 52512 3896 53389 3924
rect 52512 3884 52518 3896
rect 53377 3893 53389 3896
rect 53423 3893 53435 3927
rect 53377 3887 53435 3893
rect 54021 3927 54079 3933
rect 54021 3893 54033 3927
rect 54067 3893 54079 3927
rect 55306 3924 55312 3936
rect 55267 3896 55312 3924
rect 54021 3887 54079 3893
rect 55306 3884 55312 3896
rect 55364 3884 55370 3936
rect 58161 3927 58219 3933
rect 58161 3893 58173 3927
rect 58207 3924 58219 3927
rect 58434 3924 58440 3936
rect 58207 3896 58440 3924
rect 58207 3893 58219 3896
rect 58161 3887 58219 3893
rect 58434 3884 58440 3896
rect 58492 3884 58498 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 3237 3723 3295 3729
rect 3237 3689 3249 3723
rect 3283 3720 3295 3723
rect 4062 3720 4068 3732
rect 3283 3692 4068 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 4062 3680 4068 3692
rect 4120 3680 4126 3732
rect 4890 3680 4896 3732
rect 4948 3720 4954 3732
rect 5718 3720 5724 3732
rect 4948 3692 5724 3720
rect 4948 3680 4954 3692
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 5902 3720 5908 3732
rect 5863 3692 5908 3720
rect 5902 3680 5908 3692
rect 5960 3680 5966 3732
rect 6086 3720 6092 3732
rect 6047 3692 6092 3720
rect 6086 3680 6092 3692
rect 6144 3680 6150 3732
rect 8294 3720 8300 3732
rect 8255 3692 8300 3720
rect 8294 3680 8300 3692
rect 8352 3680 8358 3732
rect 9122 3680 9128 3732
rect 9180 3720 9186 3732
rect 9401 3723 9459 3729
rect 9401 3720 9413 3723
rect 9180 3692 9413 3720
rect 9180 3680 9186 3692
rect 9401 3689 9413 3692
rect 9447 3689 9459 3723
rect 9401 3683 9459 3689
rect 9490 3680 9496 3732
rect 9548 3680 9554 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 10505 3723 10563 3729
rect 10505 3720 10517 3723
rect 9640 3692 10517 3720
rect 9640 3680 9646 3692
rect 10505 3689 10517 3692
rect 10551 3689 10563 3723
rect 10505 3683 10563 3689
rect 12253 3723 12311 3729
rect 12253 3689 12265 3723
rect 12299 3720 12311 3723
rect 14366 3720 14372 3732
rect 12299 3692 14372 3720
rect 12299 3689 12311 3692
rect 12253 3683 12311 3689
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 16114 3720 16120 3732
rect 16075 3692 16120 3720
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 17037 3723 17095 3729
rect 17037 3689 17049 3723
rect 17083 3720 17095 3723
rect 17126 3720 17132 3732
rect 17083 3692 17132 3720
rect 17083 3689 17095 3692
rect 17037 3683 17095 3689
rect 17126 3680 17132 3692
rect 17184 3680 17190 3732
rect 17770 3720 17776 3732
rect 17731 3692 17776 3720
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 18598 3720 18604 3732
rect 18559 3692 18604 3720
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 18782 3680 18788 3732
rect 18840 3720 18846 3732
rect 20993 3723 21051 3729
rect 20993 3720 21005 3723
rect 18840 3692 21005 3720
rect 18840 3680 18846 3692
rect 20993 3689 21005 3692
rect 21039 3689 21051 3723
rect 27982 3720 27988 3732
rect 27943 3692 27988 3720
rect 20993 3683 21051 3689
rect 27982 3680 27988 3692
rect 28040 3680 28046 3732
rect 32398 3720 32404 3732
rect 32359 3692 32404 3720
rect 32398 3680 32404 3692
rect 32456 3680 32462 3732
rect 52730 3680 52736 3732
rect 52788 3720 52794 3732
rect 52788 3692 55214 3720
rect 52788 3680 52794 3692
rect 3418 3612 3424 3664
rect 3476 3652 3482 3664
rect 3786 3652 3792 3664
rect 3476 3624 3792 3652
rect 3476 3612 3482 3624
rect 3786 3612 3792 3624
rect 3844 3652 3850 3664
rect 3881 3655 3939 3661
rect 3881 3652 3893 3655
rect 3844 3624 3893 3652
rect 3844 3612 3850 3624
rect 3881 3621 3893 3624
rect 3927 3621 3939 3655
rect 3881 3615 3939 3621
rect 7558 3612 7564 3664
rect 7616 3652 7622 3664
rect 8754 3652 8760 3664
rect 7616 3624 8760 3652
rect 7616 3612 7622 3624
rect 8754 3612 8760 3624
rect 8812 3652 8818 3664
rect 8941 3655 8999 3661
rect 8941 3652 8953 3655
rect 8812 3624 8953 3652
rect 8812 3612 8818 3624
rect 8941 3621 8953 3624
rect 8987 3621 8999 3655
rect 8941 3615 8999 3621
rect 9030 3612 9036 3664
rect 9088 3652 9094 3664
rect 9309 3655 9367 3661
rect 9309 3652 9321 3655
rect 9088 3624 9321 3652
rect 9088 3612 9094 3624
rect 9309 3621 9321 3624
rect 9355 3652 9367 3655
rect 9508 3652 9536 3680
rect 9355 3624 9536 3652
rect 13541 3655 13599 3661
rect 9355 3621 9367 3624
rect 9309 3615 9367 3621
rect 13541 3621 13553 3655
rect 13587 3652 13599 3655
rect 14829 3655 14887 3661
rect 14829 3652 14841 3655
rect 13587 3624 14841 3652
rect 13587 3621 13599 3624
rect 13541 3615 13599 3621
rect 14829 3621 14841 3624
rect 14875 3621 14887 3655
rect 14829 3615 14887 3621
rect 16850 3612 16856 3664
rect 16908 3652 16914 3664
rect 17954 3652 17960 3664
rect 16908 3624 17960 3652
rect 16908 3612 16914 3624
rect 17954 3612 17960 3624
rect 18012 3612 18018 3664
rect 20346 3652 20352 3664
rect 20307 3624 20352 3652
rect 20346 3612 20352 3624
rect 20404 3612 20410 3664
rect 21358 3612 21364 3664
rect 21416 3652 21422 3664
rect 21729 3655 21787 3661
rect 21729 3652 21741 3655
rect 21416 3624 21741 3652
rect 21416 3612 21422 3624
rect 21729 3621 21741 3624
rect 21775 3621 21787 3655
rect 21729 3615 21787 3621
rect 26142 3612 26148 3664
rect 26200 3652 26206 3664
rect 26200 3624 26648 3652
rect 26200 3612 26206 3624
rect 5261 3587 5319 3593
rect 5261 3553 5273 3587
rect 5307 3584 5319 3587
rect 5442 3584 5448 3596
rect 5307 3556 5448 3584
rect 5307 3553 5319 3556
rect 5261 3547 5319 3553
rect 1854 3516 1860 3528
rect 1767 3488 1860 3516
rect 1854 3476 1860 3488
rect 1912 3516 1918 3528
rect 2406 3516 2412 3528
rect 1912 3488 2412 3516
rect 1912 3476 1918 3488
rect 2406 3476 2412 3488
rect 2464 3516 2470 3528
rect 5276 3516 5304 3547
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 6549 3587 6607 3593
rect 6549 3584 6561 3587
rect 6512 3556 6561 3584
rect 6512 3544 6518 3556
rect 6549 3553 6561 3556
rect 6595 3553 6607 3587
rect 6822 3584 6828 3596
rect 6783 3556 6828 3584
rect 6549 3547 6607 3553
rect 6822 3544 6828 3556
rect 6880 3584 6886 3596
rect 6880 3556 8616 3584
rect 6880 3544 6886 3556
rect 2464 3488 5304 3516
rect 2464 3476 2470 3488
rect 5350 3476 5356 3528
rect 5408 3516 5414 3528
rect 5408 3488 6592 3516
rect 5408 3476 5414 3488
rect 6564 3460 6592 3488
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 7800 3488 8033 3516
rect 7800 3476 7806 3488
rect 8021 3485 8033 3488
rect 8067 3516 8079 3519
rect 8202 3516 8208 3528
rect 8067 3488 8208 3516
rect 8067 3485 8079 3488
rect 8021 3479 8079 3485
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8588 3516 8616 3556
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 9493 3587 9551 3593
rect 9493 3584 9505 3587
rect 8720 3556 9505 3584
rect 8720 3544 8726 3556
rect 9493 3553 9505 3556
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 9861 3587 9919 3593
rect 9861 3553 9873 3587
rect 9907 3584 9919 3587
rect 12618 3584 12624 3596
rect 9907 3556 12624 3584
rect 9907 3553 9919 3556
rect 9861 3547 9919 3553
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 12728 3556 13860 3584
rect 9398 3516 9404 3528
rect 8588 3488 9404 3516
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 9582 3476 9588 3528
rect 9640 3516 9646 3528
rect 10318 3516 10324 3528
rect 9640 3488 10324 3516
rect 9640 3476 9646 3488
rect 10318 3476 10324 3488
rect 10376 3476 10382 3528
rect 10686 3476 10692 3528
rect 10744 3516 10750 3528
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 10744 3488 11069 3516
rect 10744 3476 10750 3488
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 11057 3479 11115 3485
rect 12526 3476 12532 3528
rect 12584 3516 12590 3528
rect 12728 3525 12756 3556
rect 12713 3519 12771 3525
rect 12713 3516 12725 3519
rect 12584 3488 12725 3516
rect 12584 3476 12590 3488
rect 12713 3485 12725 3488
rect 12759 3485 12771 3519
rect 12713 3479 12771 3485
rect 13170 3476 13176 3528
rect 13228 3516 13234 3528
rect 13357 3519 13415 3525
rect 13357 3516 13369 3519
rect 13228 3488 13369 3516
rect 13228 3476 13234 3488
rect 13357 3485 13369 3488
rect 13403 3485 13415 3519
rect 13832 3516 13860 3556
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 14369 3587 14427 3593
rect 14369 3584 14381 3587
rect 13964 3556 14381 3584
rect 13964 3544 13970 3556
rect 14369 3553 14381 3556
rect 14415 3553 14427 3587
rect 14369 3547 14427 3553
rect 15838 3544 15844 3596
rect 15896 3584 15902 3596
rect 17494 3584 17500 3596
rect 15896 3556 17500 3584
rect 15896 3544 15902 3556
rect 17494 3544 17500 3556
rect 17552 3584 17558 3596
rect 19613 3587 19671 3593
rect 17552 3556 17632 3584
rect 17552 3544 17558 3556
rect 14458 3516 14464 3528
rect 13832 3488 14464 3516
rect 13357 3479 13415 3485
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 15746 3476 15752 3528
rect 15804 3516 15810 3528
rect 15933 3519 15991 3525
rect 15933 3516 15945 3519
rect 15804 3488 15945 3516
rect 15804 3476 15810 3488
rect 15933 3485 15945 3488
rect 15979 3516 15991 3519
rect 16574 3516 16580 3528
rect 15979 3488 16580 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 16850 3516 16856 3528
rect 16811 3488 16856 3516
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 17604 3525 17632 3556
rect 19613 3553 19625 3587
rect 19659 3584 19671 3587
rect 21450 3584 21456 3596
rect 19659 3556 21456 3584
rect 19659 3553 19671 3556
rect 19613 3547 19671 3553
rect 21450 3544 21456 3556
rect 21508 3544 21514 3596
rect 26620 3593 26648 3624
rect 46290 3612 46296 3664
rect 46348 3652 46354 3664
rect 46937 3655 46995 3661
rect 46937 3652 46949 3655
rect 46348 3624 46949 3652
rect 46348 3612 46354 3624
rect 46937 3621 46949 3624
rect 46983 3621 46995 3655
rect 46937 3615 46995 3621
rect 51442 3612 51448 3664
rect 51500 3652 51506 3664
rect 52825 3655 52883 3661
rect 52825 3652 52837 3655
rect 51500 3624 52837 3652
rect 51500 3612 51506 3624
rect 52825 3621 52837 3624
rect 52871 3621 52883 3655
rect 55186 3652 55214 3692
rect 55309 3655 55367 3661
rect 55309 3652 55321 3655
rect 55186 3624 55321 3652
rect 52825 3615 52883 3621
rect 55309 3621 55321 3624
rect 55355 3621 55367 3655
rect 55309 3615 55367 3621
rect 26605 3587 26663 3593
rect 26605 3553 26617 3587
rect 26651 3553 26663 3587
rect 31018 3584 31024 3596
rect 30979 3556 31024 3584
rect 26605 3547 26663 3553
rect 31018 3544 31024 3556
rect 31076 3544 31082 3596
rect 50798 3544 50804 3596
rect 50856 3584 50862 3596
rect 51537 3587 51595 3593
rect 51537 3584 51549 3587
rect 50856 3556 51549 3584
rect 50856 3544 50862 3556
rect 51537 3553 51549 3556
rect 51583 3553 51595 3587
rect 51537 3547 51595 3553
rect 51626 3544 51632 3596
rect 51684 3584 51690 3596
rect 53469 3587 53527 3593
rect 53469 3584 53481 3587
rect 51684 3556 53481 3584
rect 51684 3544 51690 3556
rect 53469 3553 53481 3556
rect 53515 3553 53527 3587
rect 53469 3547 53527 3553
rect 53834 3544 53840 3596
rect 53892 3584 53898 3596
rect 56597 3587 56655 3593
rect 56597 3584 56609 3587
rect 53892 3556 56609 3584
rect 53892 3544 53898 3556
rect 56597 3553 56609 3556
rect 56643 3553 56655 3587
rect 56597 3547 56655 3553
rect 17589 3519 17647 3525
rect 17589 3485 17601 3519
rect 17635 3485 17647 3519
rect 17589 3479 17647 3485
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 18509 3519 18567 3525
rect 18509 3516 18521 3519
rect 18380 3488 18521 3516
rect 18380 3476 18386 3488
rect 18509 3485 18521 3488
rect 18555 3485 18567 3519
rect 18509 3479 18567 3485
rect 20806 3476 20812 3528
rect 20864 3516 20870 3528
rect 21085 3519 21143 3525
rect 21085 3516 21097 3519
rect 20864 3488 21097 3516
rect 20864 3476 20870 3488
rect 21085 3485 21097 3488
rect 21131 3485 21143 3519
rect 21085 3479 21143 3485
rect 21634 3476 21640 3528
rect 21692 3516 21698 3528
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21692 3488 21925 3516
rect 21692 3476 21698 3488
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3516 23259 3519
rect 23658 3516 23664 3528
rect 23247 3488 23664 3516
rect 23247 3485 23259 3488
rect 23201 3479 23259 3485
rect 23658 3476 23664 3488
rect 23716 3476 23722 3528
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3516 23903 3519
rect 23934 3516 23940 3528
rect 23891 3488 23940 3516
rect 23891 3485 23903 3488
rect 23845 3479 23903 3485
rect 23934 3476 23940 3488
rect 23992 3476 23998 3528
rect 24673 3519 24731 3525
rect 24673 3485 24685 3519
rect 24719 3516 24731 3519
rect 24762 3516 24768 3528
rect 24719 3488 24768 3516
rect 24719 3485 24731 3488
rect 24673 3479 24731 3485
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 25501 3519 25559 3525
rect 25501 3485 25513 3519
rect 25547 3516 25559 3519
rect 25590 3516 25596 3528
rect 25547 3488 25596 3516
rect 25547 3485 25559 3488
rect 25501 3479 25559 3485
rect 25590 3476 25596 3488
rect 25648 3476 25654 3528
rect 26142 3516 26148 3528
rect 26103 3488 26148 3516
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26878 3525 26884 3528
rect 26872 3516 26884 3525
rect 26839 3488 26884 3516
rect 26872 3479 26884 3488
rect 26878 3476 26884 3479
rect 26936 3476 26942 3528
rect 28626 3476 28632 3528
rect 28684 3516 28690 3528
rect 28721 3519 28779 3525
rect 28721 3516 28733 3519
rect 28684 3488 28733 3516
rect 28684 3476 28690 3488
rect 28721 3485 28733 3488
rect 28767 3485 28779 3519
rect 28721 3479 28779 3485
rect 30650 3476 30656 3528
rect 30708 3516 30714 3528
rect 31277 3519 31335 3525
rect 31277 3516 31289 3519
rect 30708 3488 31289 3516
rect 30708 3476 30714 3488
rect 31277 3485 31289 3488
rect 31323 3485 31335 3519
rect 31277 3479 31335 3485
rect 34698 3476 34704 3528
rect 34756 3516 34762 3528
rect 34793 3519 34851 3525
rect 34793 3516 34805 3519
rect 34756 3488 34805 3516
rect 34756 3476 34762 3488
rect 34793 3485 34805 3488
rect 34839 3485 34851 3519
rect 34793 3479 34851 3485
rect 35342 3476 35348 3528
rect 35400 3516 35406 3528
rect 35437 3519 35495 3525
rect 35437 3516 35449 3519
rect 35400 3488 35449 3516
rect 35400 3476 35406 3488
rect 35437 3485 35449 3488
rect 35483 3485 35495 3519
rect 35437 3479 35495 3485
rect 35802 3476 35808 3528
rect 35860 3516 35866 3528
rect 36081 3519 36139 3525
rect 36081 3516 36093 3519
rect 35860 3488 36093 3516
rect 35860 3476 35866 3488
rect 36081 3485 36093 3488
rect 36127 3485 36139 3519
rect 36081 3479 36139 3485
rect 36630 3476 36636 3528
rect 36688 3516 36694 3528
rect 36725 3519 36783 3525
rect 36725 3516 36737 3519
rect 36688 3488 36737 3516
rect 36688 3476 36694 3488
rect 36725 3485 36737 3488
rect 36771 3485 36783 3519
rect 36725 3479 36783 3485
rect 37458 3476 37464 3528
rect 37516 3516 37522 3528
rect 37553 3519 37611 3525
rect 37553 3516 37565 3519
rect 37516 3488 37565 3516
rect 37516 3476 37522 3488
rect 37553 3485 37565 3488
rect 37599 3485 37611 3519
rect 37553 3479 37611 3485
rect 38562 3476 38568 3528
rect 38620 3516 38626 3528
rect 38657 3519 38715 3525
rect 38657 3516 38669 3519
rect 38620 3488 38669 3516
rect 38620 3476 38626 3488
rect 38657 3485 38669 3488
rect 38703 3485 38715 3519
rect 38657 3479 38715 3485
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 40000 3488 40049 3516
rect 40000 3476 40006 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 40494 3476 40500 3528
rect 40552 3516 40558 3528
rect 40681 3519 40739 3525
rect 40681 3516 40693 3519
rect 40552 3488 40693 3516
rect 40552 3476 40558 3488
rect 40681 3485 40693 3488
rect 40727 3485 40739 3519
rect 40681 3479 40739 3485
rect 41046 3476 41052 3528
rect 41104 3516 41110 3528
rect 41325 3519 41383 3525
rect 41325 3516 41337 3519
rect 41104 3488 41337 3516
rect 41104 3476 41110 3488
rect 41325 3485 41337 3488
rect 41371 3485 41383 3519
rect 41325 3479 41383 3485
rect 42426 3476 42432 3528
rect 42484 3516 42490 3528
rect 42521 3519 42579 3525
rect 42521 3516 42533 3519
rect 42484 3488 42533 3516
rect 42484 3476 42490 3488
rect 42521 3485 42533 3488
rect 42567 3485 42579 3519
rect 42521 3479 42579 3485
rect 42702 3476 42708 3528
rect 42760 3516 42766 3528
rect 43165 3519 43223 3525
rect 43165 3516 43177 3519
rect 42760 3488 43177 3516
rect 42760 3476 42766 3488
rect 43165 3485 43177 3488
rect 43211 3485 43223 3519
rect 43165 3479 43223 3485
rect 44358 3476 44364 3528
rect 44416 3516 44422 3528
rect 45005 3519 45063 3525
rect 45005 3516 45017 3519
rect 44416 3488 45017 3516
rect 44416 3476 44422 3488
rect 45005 3485 45017 3488
rect 45051 3485 45063 3519
rect 45005 3479 45063 3485
rect 45186 3476 45192 3528
rect 45244 3516 45250 3528
rect 45649 3519 45707 3525
rect 45649 3516 45661 3519
rect 45244 3488 45661 3516
rect 45244 3476 45250 3488
rect 45649 3485 45661 3488
rect 45695 3485 45707 3519
rect 45649 3479 45707 3485
rect 46014 3476 46020 3528
rect 46072 3516 46078 3528
rect 46293 3519 46351 3525
rect 46293 3516 46305 3519
rect 46072 3488 46305 3516
rect 46072 3476 46078 3488
rect 46293 3485 46305 3488
rect 46339 3485 46351 3519
rect 46293 3479 46351 3485
rect 47670 3476 47676 3528
rect 47728 3516 47734 3528
rect 47765 3519 47823 3525
rect 47765 3516 47777 3519
rect 47728 3488 47777 3516
rect 47728 3476 47734 3488
rect 47765 3485 47777 3488
rect 47811 3485 47823 3519
rect 47765 3479 47823 3485
rect 48222 3476 48228 3528
rect 48280 3516 48286 3528
rect 48409 3519 48467 3525
rect 48409 3516 48421 3519
rect 48280 3488 48421 3516
rect 48280 3476 48286 3488
rect 48409 3485 48421 3488
rect 48455 3485 48467 3519
rect 48409 3479 48467 3485
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50249 3519 50307 3525
rect 50249 3516 50261 3519
rect 50212 3488 50261 3516
rect 50212 3476 50218 3488
rect 50249 3485 50261 3488
rect 50295 3485 50307 3519
rect 50249 3479 50307 3485
rect 50614 3476 50620 3528
rect 50672 3516 50678 3528
rect 50893 3519 50951 3525
rect 50893 3516 50905 3519
rect 50672 3488 50905 3516
rect 50672 3476 50678 3488
rect 50893 3485 50905 3488
rect 50939 3485 50951 3519
rect 50893 3479 50951 3485
rect 51166 3476 51172 3528
rect 51224 3516 51230 3528
rect 52181 3519 52239 3525
rect 52181 3516 52193 3519
rect 51224 3488 52193 3516
rect 51224 3476 51230 3488
rect 52181 3485 52193 3488
rect 52227 3485 52239 3519
rect 52181 3479 52239 3485
rect 52270 3476 52276 3528
rect 52328 3516 52334 3528
rect 54113 3519 54171 3525
rect 54113 3516 54125 3519
rect 52328 3488 54125 3516
rect 52328 3476 52334 3488
rect 54113 3485 54125 3488
rect 54159 3485 54171 3519
rect 55953 3519 56011 3525
rect 55953 3516 55965 3519
rect 54113 3479 54171 3485
rect 55186 3488 55965 3516
rect 2130 3457 2136 3460
rect 2124 3448 2136 3457
rect 2091 3420 2136 3448
rect 2124 3411 2136 3420
rect 2130 3408 2136 3411
rect 2188 3408 2194 3460
rect 5016 3451 5074 3457
rect 5016 3417 5028 3451
rect 5062 3448 5074 3451
rect 5258 3448 5264 3460
rect 5062 3420 5264 3448
rect 5062 3417 5074 3420
rect 5016 3411 5074 3417
rect 5258 3408 5264 3420
rect 5316 3408 5322 3460
rect 5626 3408 5632 3460
rect 5684 3448 5690 3460
rect 5721 3451 5779 3457
rect 5721 3448 5733 3451
rect 5684 3420 5733 3448
rect 5684 3408 5690 3420
rect 5721 3417 5733 3420
rect 5767 3417 5779 3451
rect 5721 3411 5779 3417
rect 6546 3408 6552 3460
rect 6604 3408 6610 3460
rect 8294 3408 8300 3460
rect 8352 3448 8358 3460
rect 14277 3451 14335 3457
rect 14277 3448 14289 3451
rect 8352 3420 11284 3448
rect 8352 3408 8358 3420
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 4890 3380 4896 3392
rect 2832 3352 4896 3380
rect 2832 3340 2838 3352
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 5902 3340 5908 3392
rect 5960 3389 5966 3392
rect 5960 3383 5979 3389
rect 5967 3349 5979 3383
rect 5960 3343 5979 3349
rect 5960 3340 5966 3343
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 9214 3380 9220 3392
rect 8628 3352 9220 3380
rect 8628 3340 8634 3352
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 11256 3389 11284 3420
rect 12912 3420 14289 3448
rect 12912 3389 12940 3420
rect 14277 3417 14289 3420
rect 14323 3417 14335 3451
rect 14826 3448 14832 3460
rect 14787 3420 14832 3448
rect 14277 3411 14335 3417
rect 14826 3408 14832 3420
rect 14884 3408 14890 3460
rect 15473 3451 15531 3457
rect 15473 3417 15485 3451
rect 15519 3448 15531 3451
rect 20165 3451 20223 3457
rect 20165 3448 20177 3451
rect 15519 3420 20177 3448
rect 15519 3417 15531 3420
rect 15473 3411 15531 3417
rect 20165 3417 20177 3420
rect 20211 3417 20223 3451
rect 20165 3411 20223 3417
rect 11241 3383 11299 3389
rect 11241 3349 11253 3383
rect 11287 3349 11299 3383
rect 11241 3343 11299 3349
rect 12897 3383 12955 3389
rect 12897 3349 12909 3383
rect 12943 3349 12955 3383
rect 14090 3380 14096 3392
rect 14051 3352 14096 3380
rect 12897 3343 12955 3349
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 16666 3340 16672 3392
rect 16724 3380 16730 3392
rect 16942 3380 16948 3392
rect 16724 3352 16948 3380
rect 16724 3340 16730 3352
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 17770 3340 17776 3392
rect 17828 3380 17834 3392
rect 19426 3380 19432 3392
rect 17828 3352 19432 3380
rect 17828 3340 17834 3352
rect 19426 3340 19432 3352
rect 19484 3340 19490 3392
rect 20180 3380 20208 3411
rect 53282 3408 53288 3460
rect 53340 3448 53346 3460
rect 55186 3448 55214 3488
rect 55953 3485 55965 3488
rect 55999 3485 56011 3519
rect 57514 3516 57520 3528
rect 57475 3488 57520 3516
rect 55953 3479 56011 3485
rect 57514 3476 57520 3488
rect 57572 3476 57578 3528
rect 58158 3516 58164 3528
rect 58119 3488 58164 3516
rect 58158 3476 58164 3488
rect 58216 3476 58222 3528
rect 53340 3420 55214 3448
rect 53340 3408 53346 3420
rect 20254 3380 20260 3392
rect 20180 3352 20260 3380
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 22557 3383 22615 3389
rect 22557 3349 22569 3383
rect 22603 3380 22615 3383
rect 22830 3380 22836 3392
rect 22603 3352 22836 3380
rect 22603 3349 22615 3352
rect 22557 3343 22615 3349
rect 22830 3340 22836 3352
rect 22888 3340 22894 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 1728 3148 3648 3176
rect 1728 3136 1734 3148
rect 2676 3111 2734 3117
rect 2676 3077 2688 3111
rect 2722 3108 2734 3111
rect 3510 3108 3516 3120
rect 2722 3080 3516 3108
rect 2722 3077 2734 3080
rect 2676 3071 2734 3077
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 3620 3108 3648 3148
rect 3694 3136 3700 3188
rect 3752 3176 3758 3188
rect 3789 3179 3847 3185
rect 3789 3176 3801 3179
rect 3752 3148 3801 3176
rect 3752 3136 3758 3148
rect 3789 3145 3801 3148
rect 3835 3176 3847 3179
rect 4062 3176 4068 3188
rect 3835 3148 4068 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 4062 3136 4068 3148
rect 4120 3136 4126 3188
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 5902 3176 5908 3188
rect 4856 3148 5908 3176
rect 4856 3136 4862 3148
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 8938 3176 8944 3188
rect 8899 3148 8944 3176
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 11609 3179 11667 3185
rect 11609 3176 11621 3179
rect 9180 3148 11621 3176
rect 9180 3136 9186 3148
rect 11609 3145 11621 3148
rect 11655 3145 11667 3179
rect 14550 3176 14556 3188
rect 14511 3148 14556 3176
rect 11609 3139 11667 3145
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 15286 3176 15292 3188
rect 15247 3148 15292 3176
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 15933 3179 15991 3185
rect 15933 3145 15945 3179
rect 15979 3176 15991 3179
rect 16114 3176 16120 3188
rect 15979 3148 16120 3176
rect 15979 3145 15991 3148
rect 15933 3139 15991 3145
rect 16114 3136 16120 3148
rect 16172 3136 16178 3188
rect 17405 3179 17463 3185
rect 17405 3145 17417 3179
rect 17451 3176 17463 3179
rect 17678 3176 17684 3188
rect 17451 3148 17684 3176
rect 17451 3145 17463 3148
rect 17405 3139 17463 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 18138 3176 18144 3188
rect 18099 3148 18144 3176
rect 18138 3136 18144 3148
rect 18196 3136 18202 3188
rect 19426 3136 19432 3188
rect 19484 3176 19490 3188
rect 19613 3179 19671 3185
rect 19613 3176 19625 3179
rect 19484 3148 19625 3176
rect 19484 3136 19490 3148
rect 19613 3145 19625 3148
rect 19659 3145 19671 3179
rect 20346 3176 20352 3188
rect 20307 3148 20352 3176
rect 19613 3139 19671 3145
rect 20346 3136 20352 3148
rect 20404 3136 20410 3188
rect 22278 3176 22284 3188
rect 22239 3148 22284 3176
rect 22278 3136 22284 3148
rect 22336 3136 22342 3188
rect 23017 3179 23075 3185
rect 23017 3145 23029 3179
rect 23063 3176 23075 3179
rect 23198 3176 23204 3188
rect 23063 3148 23204 3176
rect 23063 3145 23075 3148
rect 23017 3139 23075 3145
rect 23198 3136 23204 3148
rect 23256 3136 23262 3188
rect 8754 3108 8760 3120
rect 3620 3080 8760 3108
rect 8754 3068 8760 3080
rect 8812 3068 8818 3120
rect 8846 3068 8852 3120
rect 8904 3108 8910 3120
rect 9214 3108 9220 3120
rect 8904 3080 9220 3108
rect 8904 3068 8910 3080
rect 9214 3068 9220 3080
rect 9272 3108 9278 3120
rect 11238 3108 11244 3120
rect 9272 3080 11244 3108
rect 9272 3068 9278 3080
rect 11238 3068 11244 3080
rect 11296 3068 11302 3120
rect 13446 3108 13452 3120
rect 11808 3080 13452 3108
rect 1762 3040 1768 3052
rect 1723 3012 1768 3040
rect 1762 3000 1768 3012
rect 1820 3000 1826 3052
rect 2406 3040 2412 3052
rect 2367 3012 2412 3040
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 5074 3040 5080 3052
rect 5035 3012 5080 3040
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 5810 3040 5816 3052
rect 5771 3012 5816 3040
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 6730 3000 6736 3052
rect 6788 3040 6794 3052
rect 7926 3040 7932 3052
rect 6788 3012 7932 3040
rect 6788 3000 6794 3012
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 8076 3012 8125 3040
rect 8076 3000 8082 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8772 3040 8800 3068
rect 9585 3043 9643 3049
rect 9585 3040 9597 3043
rect 8772 3012 9597 3040
rect 8113 3003 8171 3009
rect 9585 3009 9597 3012
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 9953 3043 10011 3049
rect 9953 3009 9965 3043
rect 9999 3040 10011 3043
rect 10042 3040 10048 3052
rect 9999 3012 10048 3040
rect 9999 3009 10011 3012
rect 9953 3003 10011 3009
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10410 3000 10416 3052
rect 10468 3040 10474 3052
rect 10505 3043 10563 3049
rect 10505 3040 10517 3043
rect 10468 3012 10517 3040
rect 10468 3000 10474 3012
rect 10505 3009 10517 3012
rect 10551 3009 10563 3043
rect 10870 3040 10876 3052
rect 10831 3012 10876 3040
rect 10505 3003 10563 3009
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11808 3049 11836 3080
rect 13446 3068 13452 3080
rect 13504 3068 13510 3120
rect 14384 3080 15332 3108
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 11793 3003 11851 3009
rect 11974 3000 11980 3052
rect 12032 3040 12038 3052
rect 12253 3043 12311 3049
rect 12253 3040 12265 3043
rect 12032 3012 12265 3040
rect 12032 3000 12038 3012
rect 12253 3009 12265 3012
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14384 3049 14412 3080
rect 15304 3052 15332 3080
rect 17862 3068 17868 3120
rect 17920 3108 17926 3120
rect 18233 3111 18291 3117
rect 18233 3108 18245 3111
rect 17920 3080 18245 3108
rect 17920 3068 17926 3080
rect 18233 3077 18245 3080
rect 18279 3108 18291 3111
rect 18598 3108 18604 3120
rect 18279 3080 18604 3108
rect 18279 3077 18291 3080
rect 18233 3071 18291 3077
rect 18598 3068 18604 3080
rect 18656 3068 18662 3120
rect 18782 3108 18788 3120
rect 18743 3080 18788 3108
rect 18782 3068 18788 3080
rect 18840 3068 18846 3120
rect 18969 3111 19027 3117
rect 18969 3077 18981 3111
rect 19015 3108 19027 3111
rect 19058 3108 19064 3120
rect 19015 3080 19064 3108
rect 19015 3077 19027 3080
rect 18969 3071 19027 3077
rect 19058 3068 19064 3080
rect 19116 3108 19122 3120
rect 20162 3108 20168 3120
rect 19116 3080 20168 3108
rect 19116 3068 19122 3080
rect 20162 3068 20168 3080
rect 20220 3068 20226 3120
rect 20441 3111 20499 3117
rect 20441 3077 20453 3111
rect 20487 3108 20499 3111
rect 20530 3108 20536 3120
rect 20487 3080 20536 3108
rect 20487 3077 20499 3080
rect 20441 3071 20499 3077
rect 20530 3068 20536 3080
rect 20588 3108 20594 3120
rect 20714 3108 20720 3120
rect 20588 3080 20720 3108
rect 20588 3068 20594 3080
rect 20714 3068 20720 3080
rect 20772 3068 20778 3120
rect 20990 3108 20996 3120
rect 20951 3080 20996 3108
rect 20990 3068 20996 3080
rect 21048 3068 21054 3120
rect 21174 3108 21180 3120
rect 21135 3080 21180 3108
rect 21174 3068 21180 3080
rect 21232 3068 21238 3120
rect 22094 3068 22100 3120
rect 22152 3108 22158 3120
rect 22189 3111 22247 3117
rect 22189 3108 22201 3111
rect 22152 3080 22201 3108
rect 22152 3068 22158 3080
rect 22189 3077 22201 3080
rect 22235 3108 22247 3111
rect 24394 3108 24400 3120
rect 22235 3080 24400 3108
rect 22235 3077 22247 3080
rect 22189 3071 22247 3077
rect 24394 3068 24400 3080
rect 24452 3068 24458 3120
rect 51902 3068 51908 3120
rect 51960 3108 51966 3120
rect 51960 3080 54708 3108
rect 51960 3068 51966 3080
rect 14369 3043 14427 3049
rect 14369 3040 14381 3043
rect 14056 3012 14381 3040
rect 14056 3000 14062 3012
rect 14369 3009 14381 3012
rect 14415 3009 14427 3043
rect 15102 3040 15108 3052
rect 15063 3012 15108 3040
rect 14369 3003 14427 3009
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 15286 3000 15292 3052
rect 15344 3000 15350 3052
rect 16117 3043 16175 3049
rect 16117 3009 16129 3043
rect 16163 3040 16175 3043
rect 16666 3040 16672 3052
rect 16163 3012 16672 3040
rect 16163 3009 16175 3012
rect 16117 3003 16175 3009
rect 16666 3000 16672 3012
rect 16724 3040 16730 3052
rect 17218 3040 17224 3052
rect 16724 3012 17224 3040
rect 16724 3000 16730 3012
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3040 17647 3043
rect 17770 3040 17776 3052
rect 17635 3012 17776 3040
rect 17635 3009 17647 3012
rect 17589 3003 17647 3009
rect 17770 3000 17776 3012
rect 17828 3000 17834 3052
rect 18506 3000 18512 3052
rect 18564 3040 18570 3052
rect 19797 3043 19855 3049
rect 18564 3012 19564 3040
rect 18564 3000 18570 3012
rect 3418 2932 3424 2984
rect 3476 2972 3482 2984
rect 5994 2972 6000 2984
rect 3476 2944 6000 2972
rect 3476 2932 3482 2944
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 6270 2932 6276 2984
rect 6328 2972 6334 2984
rect 6822 2972 6828 2984
rect 6328 2944 6828 2972
rect 6328 2932 6334 2944
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 7098 2972 7104 2984
rect 7059 2944 7104 2972
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 7650 2932 7656 2984
rect 7708 2972 7714 2984
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 7708 2944 8677 2972
rect 7708 2932 7714 2944
rect 8665 2941 8677 2944
rect 8711 2941 8723 2975
rect 8665 2935 8723 2941
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 10428 2972 10456 3000
rect 8996 2944 10456 2972
rect 13909 2975 13967 2981
rect 8996 2932 9002 2944
rect 13909 2941 13921 2975
rect 13955 2972 13967 2975
rect 17310 2972 17316 2984
rect 13955 2944 17316 2972
rect 13955 2941 13967 2944
rect 13909 2935 13967 2941
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 4341 2907 4399 2913
rect 4341 2873 4353 2907
rect 4387 2904 4399 2907
rect 5442 2904 5448 2916
rect 4387 2876 5448 2904
rect 4387 2873 4399 2876
rect 4341 2867 4399 2873
rect 5442 2864 5448 2876
rect 5500 2864 5506 2916
rect 7374 2904 7380 2916
rect 5552 2876 7380 2904
rect 1949 2839 2007 2845
rect 1949 2805 1961 2839
rect 1995 2836 2007 2839
rect 3602 2836 3608 2848
rect 1995 2808 3608 2836
rect 1995 2805 2007 2808
rect 1949 2799 2007 2805
rect 3602 2796 3608 2808
rect 3660 2796 3666 2848
rect 4893 2839 4951 2845
rect 4893 2805 4905 2839
rect 4939 2836 4951 2839
rect 5552 2836 5580 2876
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 8573 2907 8631 2913
rect 8573 2873 8585 2907
rect 8619 2904 8631 2907
rect 9030 2904 9036 2916
rect 8619 2876 9036 2904
rect 8619 2873 8631 2876
rect 8573 2867 8631 2873
rect 9030 2864 9036 2876
rect 9088 2864 9094 2916
rect 13265 2907 13323 2913
rect 13265 2873 13277 2907
rect 13311 2904 13323 2907
rect 16482 2904 16488 2916
rect 13311 2876 16488 2904
rect 13311 2873 13323 2876
rect 13265 2867 13323 2873
rect 16482 2864 16488 2876
rect 16540 2864 16546 2916
rect 16853 2907 16911 2913
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 19426 2904 19432 2916
rect 16899 2876 19432 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 19536 2904 19564 3012
rect 19797 3009 19809 3043
rect 19843 3040 19855 3043
rect 19978 3040 19984 3052
rect 19843 3012 19984 3040
rect 19843 3009 19855 3012
rect 19797 3003 19855 3009
rect 19978 3000 19984 3012
rect 20036 3000 20042 3052
rect 22830 3040 22836 3052
rect 22791 3012 22836 3040
rect 22830 3000 22836 3012
rect 22888 3000 22894 3052
rect 51718 3000 51724 3052
rect 51776 3040 51782 3052
rect 54680 3049 54708 3080
rect 54021 3043 54079 3049
rect 54021 3040 54033 3043
rect 51776 3012 54033 3040
rect 51776 3000 51782 3012
rect 54021 3009 54033 3012
rect 54067 3009 54079 3043
rect 54021 3003 54079 3009
rect 54665 3043 54723 3049
rect 54665 3009 54677 3043
rect 54711 3009 54723 3043
rect 54665 3003 54723 3009
rect 54754 3000 54760 3052
rect 54812 3040 54818 3052
rect 55309 3043 55367 3049
rect 55309 3040 55321 3043
rect 54812 3012 55321 3040
rect 54812 3000 54818 3012
rect 55309 3009 55321 3012
rect 55355 3009 55367 3043
rect 55309 3003 55367 3009
rect 20254 2932 20260 2984
rect 20312 2972 20318 2984
rect 20438 2972 20444 2984
rect 20312 2944 20444 2972
rect 20312 2932 20318 2944
rect 20438 2932 20444 2944
rect 20496 2932 20502 2984
rect 23845 2975 23903 2981
rect 23845 2941 23857 2975
rect 23891 2972 23903 2975
rect 24486 2972 24492 2984
rect 23891 2944 24492 2972
rect 23891 2941 23903 2944
rect 23845 2935 23903 2941
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 25777 2975 25835 2981
rect 25777 2941 25789 2975
rect 25823 2972 25835 2975
rect 26418 2972 26424 2984
rect 25823 2944 26424 2972
rect 25823 2941 25835 2944
rect 25777 2935 25835 2941
rect 26418 2932 26424 2944
rect 26476 2932 26482 2984
rect 32766 2932 32772 2984
rect 32824 2972 32830 2984
rect 33413 2975 33471 2981
rect 33413 2972 33425 2975
rect 32824 2944 33425 2972
rect 32824 2932 32830 2944
rect 33413 2941 33425 2944
rect 33459 2941 33471 2975
rect 33413 2935 33471 2941
rect 38286 2932 38292 2984
rect 38344 2972 38350 2984
rect 39209 2975 39267 2981
rect 39209 2972 39221 2975
rect 38344 2944 39221 2972
rect 38344 2932 38350 2944
rect 39209 2941 39221 2944
rect 39255 2941 39267 2975
rect 39209 2935 39267 2941
rect 42150 2932 42156 2984
rect 42208 2972 42214 2984
rect 43073 2975 43131 2981
rect 43073 2972 43085 2975
rect 42208 2944 43085 2972
rect 42208 2932 42214 2944
rect 43073 2941 43085 2944
rect 43119 2941 43131 2975
rect 43073 2935 43131 2941
rect 53098 2932 53104 2984
rect 53156 2972 53162 2984
rect 55953 2975 56011 2981
rect 55953 2972 55965 2975
rect 53156 2944 55965 2972
rect 53156 2932 53162 2944
rect 55953 2941 55965 2944
rect 55999 2941 56011 2975
rect 56594 2972 56600 2984
rect 56555 2944 56600 2972
rect 55953 2935 56011 2941
rect 56594 2932 56600 2944
rect 56652 2932 56658 2984
rect 23290 2904 23296 2916
rect 19536 2876 23296 2904
rect 23290 2864 23296 2876
rect 23348 2864 23354 2916
rect 33318 2864 33324 2916
rect 33376 2904 33382 2916
rect 34057 2907 34115 2913
rect 34057 2904 34069 2907
rect 33376 2876 34069 2904
rect 33376 2864 33382 2876
rect 34057 2873 34069 2876
rect 34103 2873 34115 2907
rect 34057 2867 34115 2873
rect 34422 2864 34428 2916
rect 34480 2904 34486 2916
rect 35345 2907 35403 2913
rect 35345 2904 35357 2907
rect 34480 2876 35357 2904
rect 34480 2864 34486 2876
rect 35345 2873 35357 2876
rect 35391 2873 35403 2907
rect 35345 2867 35403 2873
rect 37182 2864 37188 2916
rect 37240 2904 37246 2916
rect 37921 2907 37979 2913
rect 37921 2904 37933 2907
rect 37240 2876 37933 2904
rect 37240 2864 37246 2876
rect 37921 2873 37933 2876
rect 37967 2873 37979 2907
rect 37921 2867 37979 2873
rect 39114 2864 39120 2916
rect 39172 2904 39178 2916
rect 39853 2907 39911 2913
rect 39853 2904 39865 2907
rect 39172 2876 39865 2904
rect 39172 2864 39178 2876
rect 39853 2873 39865 2876
rect 39899 2873 39911 2907
rect 39853 2867 39911 2873
rect 40218 2864 40224 2916
rect 40276 2904 40282 2916
rect 41141 2907 41199 2913
rect 41141 2904 41153 2907
rect 40276 2876 41153 2904
rect 40276 2864 40282 2876
rect 41141 2873 41153 2876
rect 41187 2873 41199 2907
rect 41141 2867 41199 2873
rect 42978 2864 42984 2916
rect 43036 2904 43042 2916
rect 43717 2907 43775 2913
rect 43717 2904 43729 2907
rect 43036 2876 43729 2904
rect 43036 2864 43042 2876
rect 43717 2873 43729 2876
rect 43763 2873 43775 2907
rect 43717 2867 43775 2873
rect 44082 2864 44088 2916
rect 44140 2904 44146 2916
rect 45005 2907 45063 2913
rect 45005 2904 45017 2907
rect 44140 2876 45017 2904
rect 44140 2864 44146 2876
rect 45005 2873 45017 2876
rect 45051 2873 45063 2907
rect 45649 2907 45707 2913
rect 45649 2904 45661 2907
rect 45005 2867 45063 2873
rect 45112 2876 45661 2904
rect 4939 2808 5580 2836
rect 5629 2839 5687 2845
rect 4939 2805 4951 2808
rect 4893 2799 4951 2805
rect 5629 2805 5641 2839
rect 5675 2836 5687 2839
rect 8018 2836 8024 2848
rect 5675 2808 8024 2836
rect 5675 2805 5687 2808
rect 5629 2799 5687 2805
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 8481 2839 8539 2845
rect 8481 2805 8493 2839
rect 8527 2836 8539 2839
rect 9490 2836 9496 2848
rect 8527 2808 9496 2836
rect 8527 2805 8539 2808
rect 8481 2799 8539 2805
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 9766 2796 9772 2848
rect 9824 2836 9830 2848
rect 12437 2839 12495 2845
rect 12437 2836 12449 2839
rect 9824 2808 12449 2836
rect 9824 2796 9830 2808
rect 12437 2805 12449 2808
rect 12483 2805 12495 2839
rect 12437 2799 12495 2805
rect 13170 2796 13176 2848
rect 13228 2836 13234 2848
rect 15010 2836 15016 2848
rect 13228 2808 15016 2836
rect 13228 2796 13234 2808
rect 15010 2796 15016 2808
rect 15068 2796 15074 2848
rect 15102 2796 15108 2848
rect 15160 2836 15166 2848
rect 15562 2836 15568 2848
rect 15160 2808 15568 2836
rect 15160 2796 15166 2808
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 18874 2796 18880 2848
rect 18932 2836 18938 2848
rect 20438 2836 20444 2848
rect 18932 2808 20444 2836
rect 18932 2796 18938 2808
rect 20438 2796 20444 2808
rect 20496 2796 20502 2848
rect 21266 2796 21272 2848
rect 21324 2836 21330 2848
rect 21818 2836 21824 2848
rect 21324 2808 21824 2836
rect 21324 2796 21330 2808
rect 21818 2796 21824 2808
rect 21876 2836 21882 2848
rect 23474 2836 23480 2848
rect 21876 2808 23480 2836
rect 21876 2796 21882 2808
rect 23474 2796 23480 2808
rect 23532 2796 23538 2848
rect 24489 2839 24547 2845
rect 24489 2805 24501 2839
rect 24535 2836 24547 2839
rect 25038 2836 25044 2848
rect 24535 2808 25044 2836
rect 24535 2805 24547 2808
rect 24489 2799 24547 2805
rect 25038 2796 25044 2808
rect 25096 2796 25102 2848
rect 25133 2839 25191 2845
rect 25133 2805 25145 2839
rect 25179 2836 25191 2839
rect 25866 2836 25872 2848
rect 25179 2808 25872 2836
rect 25179 2805 25191 2808
rect 25133 2799 25191 2805
rect 25866 2796 25872 2808
rect 25924 2796 25930 2848
rect 26421 2839 26479 2845
rect 26421 2805 26433 2839
rect 26467 2836 26479 2839
rect 26970 2836 26976 2848
rect 26467 2808 26976 2836
rect 26467 2805 26479 2808
rect 26421 2799 26479 2805
rect 26970 2796 26976 2808
rect 27028 2796 27034 2848
rect 27617 2839 27675 2845
rect 27617 2805 27629 2839
rect 27663 2836 27675 2839
rect 27798 2836 27804 2848
rect 27663 2808 27804 2836
rect 27663 2805 27675 2808
rect 27617 2799 27675 2805
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 28074 2836 28080 2848
rect 28035 2808 28080 2836
rect 28074 2796 28080 2808
rect 28132 2796 28138 2848
rect 28905 2839 28963 2845
rect 28905 2805 28917 2839
rect 28951 2836 28963 2839
rect 29178 2836 29184 2848
rect 28951 2808 29184 2836
rect 28951 2805 28963 2808
rect 28905 2799 28963 2805
rect 29178 2796 29184 2808
rect 29236 2796 29242 2848
rect 29549 2839 29607 2845
rect 29549 2805 29561 2839
rect 29595 2836 29607 2839
rect 29730 2836 29736 2848
rect 29595 2808 29736 2836
rect 29595 2805 29607 2808
rect 29549 2799 29607 2805
rect 29730 2796 29736 2808
rect 29788 2796 29794 2848
rect 30006 2836 30012 2848
rect 29967 2808 30012 2836
rect 30006 2796 30012 2808
rect 30064 2796 30070 2848
rect 30558 2796 30564 2848
rect 30616 2836 30622 2848
rect 30653 2839 30711 2845
rect 30653 2836 30665 2839
rect 30616 2808 30665 2836
rect 30616 2796 30622 2808
rect 30653 2805 30665 2808
rect 30699 2805 30711 2839
rect 30653 2799 30711 2805
rect 31662 2796 31668 2848
rect 31720 2836 31726 2848
rect 32125 2839 32183 2845
rect 32125 2836 32137 2839
rect 31720 2808 32137 2836
rect 31720 2796 31726 2808
rect 32125 2805 32137 2808
rect 32171 2805 32183 2839
rect 32125 2799 32183 2805
rect 32214 2796 32220 2848
rect 32272 2836 32278 2848
rect 32769 2839 32827 2845
rect 32769 2836 32781 2839
rect 32272 2808 32781 2836
rect 32272 2796 32278 2808
rect 32769 2805 32781 2808
rect 32815 2805 32827 2839
rect 32769 2799 32827 2805
rect 33870 2796 33876 2848
rect 33928 2836 33934 2848
rect 34701 2839 34759 2845
rect 34701 2836 34713 2839
rect 33928 2808 34713 2836
rect 33928 2796 33934 2808
rect 34701 2805 34713 2808
rect 34747 2805 34759 2839
rect 34701 2799 34759 2805
rect 35434 2796 35440 2848
rect 35492 2836 35498 2848
rect 35989 2839 36047 2845
rect 35989 2836 36001 2839
rect 35492 2808 36001 2836
rect 35492 2796 35498 2808
rect 35989 2805 36001 2808
rect 36035 2805 36047 2839
rect 35989 2799 36047 2805
rect 36354 2796 36360 2848
rect 36412 2836 36418 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36412 2808 37289 2836
rect 36412 2796 36418 2808
rect 37277 2805 37289 2808
rect 37323 2805 37335 2839
rect 37277 2799 37335 2805
rect 37734 2796 37740 2848
rect 37792 2836 37798 2848
rect 38565 2839 38623 2845
rect 38565 2836 38577 2839
rect 37792 2808 38577 2836
rect 37792 2796 37798 2808
rect 38565 2805 38577 2808
rect 38611 2805 38623 2839
rect 38565 2799 38623 2805
rect 39666 2796 39672 2848
rect 39724 2836 39730 2848
rect 40497 2839 40555 2845
rect 40497 2836 40509 2839
rect 39724 2808 40509 2836
rect 39724 2796 39730 2808
rect 40497 2805 40509 2808
rect 40543 2805 40555 2839
rect 40497 2799 40555 2805
rect 41598 2796 41604 2848
rect 41656 2836 41662 2848
rect 42429 2839 42487 2845
rect 42429 2836 42441 2839
rect 41656 2808 42441 2836
rect 41656 2796 41662 2808
rect 42429 2805 42441 2808
rect 42475 2805 42487 2839
rect 42429 2799 42487 2805
rect 43530 2796 43536 2848
rect 43588 2836 43594 2848
rect 44361 2839 44419 2845
rect 44361 2836 44373 2839
rect 43588 2808 44373 2836
rect 43588 2796 43594 2808
rect 44361 2805 44373 2808
rect 44407 2805 44419 2839
rect 44361 2799 44419 2805
rect 44910 2796 44916 2848
rect 44968 2836 44974 2848
rect 45112 2836 45140 2876
rect 45649 2873 45661 2876
rect 45695 2873 45707 2907
rect 45649 2867 45707 2873
rect 47394 2864 47400 2916
rect 47452 2904 47458 2916
rect 48225 2907 48283 2913
rect 48225 2904 48237 2907
rect 47452 2876 48237 2904
rect 47452 2864 47458 2876
rect 48225 2873 48237 2876
rect 48271 2873 48283 2907
rect 48225 2867 48283 2873
rect 48774 2864 48780 2916
rect 48832 2904 48838 2916
rect 49513 2907 49571 2913
rect 49513 2904 49525 2907
rect 48832 2876 49525 2904
rect 48832 2864 48838 2876
rect 49513 2873 49525 2876
rect 49559 2873 49571 2907
rect 49513 2867 49571 2873
rect 49878 2864 49884 2916
rect 49936 2904 49942 2916
rect 50801 2907 50859 2913
rect 50801 2904 50813 2907
rect 49936 2876 50813 2904
rect 49936 2864 49942 2876
rect 50801 2873 50813 2876
rect 50847 2873 50859 2907
rect 50801 2867 50859 2873
rect 50982 2864 50988 2916
rect 51040 2904 51046 2916
rect 52733 2907 52791 2913
rect 52733 2904 52745 2907
rect 51040 2876 52745 2904
rect 51040 2864 51046 2876
rect 52733 2873 52745 2876
rect 52779 2873 52791 2907
rect 52733 2867 52791 2873
rect 54202 2864 54208 2916
rect 54260 2904 54266 2916
rect 57885 2907 57943 2913
rect 57885 2904 57897 2907
rect 54260 2876 57897 2904
rect 54260 2864 54266 2876
rect 57885 2873 57897 2876
rect 57931 2873 57943 2907
rect 57885 2867 57943 2873
rect 44968 2808 45140 2836
rect 44968 2796 44974 2808
rect 45462 2796 45468 2848
rect 45520 2836 45526 2848
rect 46293 2839 46351 2845
rect 46293 2836 46305 2839
rect 45520 2808 46305 2836
rect 45520 2796 45526 2808
rect 46293 2805 46305 2808
rect 46339 2805 46351 2839
rect 46293 2799 46351 2805
rect 46842 2796 46848 2848
rect 46900 2836 46906 2848
rect 47581 2839 47639 2845
rect 47581 2836 47593 2839
rect 46900 2808 47593 2836
rect 46900 2796 46906 2808
rect 47581 2805 47593 2808
rect 47627 2805 47639 2839
rect 47581 2799 47639 2805
rect 47946 2796 47952 2848
rect 48004 2836 48010 2848
rect 48869 2839 48927 2845
rect 48869 2836 48881 2839
rect 48004 2808 48881 2836
rect 48004 2796 48010 2808
rect 48869 2805 48881 2808
rect 48915 2805 48927 2839
rect 48869 2799 48927 2805
rect 49326 2796 49332 2848
rect 49384 2836 49390 2848
rect 50157 2839 50215 2845
rect 50157 2836 50169 2839
rect 49384 2808 50169 2836
rect 49384 2796 49390 2808
rect 50157 2805 50169 2808
rect 50203 2805 50215 2839
rect 50157 2799 50215 2805
rect 50706 2796 50712 2848
rect 50764 2836 50770 2848
rect 51445 2839 51503 2845
rect 51445 2836 51457 2839
rect 50764 2808 51457 2836
rect 50764 2796 50770 2808
rect 51445 2805 51457 2808
rect 51491 2805 51503 2839
rect 51445 2799 51503 2805
rect 51534 2796 51540 2848
rect 51592 2836 51598 2848
rect 53377 2839 53435 2845
rect 53377 2836 53389 2839
rect 51592 2808 53389 2836
rect 51592 2796 51598 2808
rect 53377 2805 53389 2808
rect 53423 2805 53435 2839
rect 53377 2799 53435 2805
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 3970 2592 3976 2644
rect 4028 2632 4034 2644
rect 5626 2632 5632 2644
rect 4028 2604 5632 2632
rect 4028 2592 4034 2604
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 10410 2632 10416 2644
rect 10371 2604 10416 2632
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 10594 2592 10600 2644
rect 10652 2632 10658 2644
rect 12437 2635 12495 2641
rect 12437 2632 12449 2635
rect 10652 2604 12449 2632
rect 10652 2592 10658 2604
rect 12437 2601 12449 2604
rect 12483 2601 12495 2635
rect 13446 2632 13452 2644
rect 13407 2604 13452 2632
rect 12437 2595 12495 2601
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 14550 2632 14556 2644
rect 14511 2604 14556 2632
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 15838 2632 15844 2644
rect 15120 2604 15844 2632
rect 2317 2567 2375 2573
rect 2317 2533 2329 2567
rect 2363 2564 2375 2567
rect 2958 2564 2964 2576
rect 2363 2536 2964 2564
rect 2363 2533 2375 2536
rect 2317 2527 2375 2533
rect 2958 2524 2964 2536
rect 3016 2524 3022 2576
rect 3053 2567 3111 2573
rect 3053 2533 3065 2567
rect 3099 2564 3111 2567
rect 7006 2564 7012 2576
rect 3099 2536 7012 2564
rect 3099 2533 3111 2536
rect 3053 2527 3111 2533
rect 7006 2524 7012 2536
rect 7064 2524 7070 2576
rect 7116 2536 9352 2564
rect 3786 2496 3792 2508
rect 2516 2468 3792 2496
rect 1578 2428 1584 2440
rect 1539 2400 1584 2428
rect 1578 2388 1584 2400
rect 1636 2388 1642 2440
rect 2516 2437 2544 2468
rect 3786 2456 3792 2468
rect 3844 2456 3850 2508
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4120 2468 4384 2496
rect 4120 2456 4126 2468
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 3234 2428 3240 2440
rect 3195 2400 3240 2428
rect 2501 2391 2559 2397
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 4249 2431 4307 2437
rect 4249 2428 4261 2431
rect 3936 2400 4261 2428
rect 3936 2388 3942 2400
rect 4249 2397 4261 2400
rect 4295 2397 4307 2431
rect 4356 2428 4384 2468
rect 4982 2456 4988 2508
rect 5040 2496 5046 2508
rect 5537 2499 5595 2505
rect 5537 2496 5549 2499
rect 5040 2468 5549 2496
rect 5040 2456 5046 2468
rect 5537 2465 5549 2468
rect 5583 2465 5595 2499
rect 7116 2496 7144 2536
rect 5537 2459 5595 2465
rect 5644 2468 7144 2496
rect 7837 2499 7895 2505
rect 5644 2428 5672 2468
rect 7837 2465 7849 2499
rect 7883 2496 7895 2499
rect 9214 2496 9220 2508
rect 7883 2468 9220 2496
rect 7883 2465 7895 2468
rect 7837 2459 7895 2465
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 4356 2400 5672 2428
rect 5813 2431 5871 2437
rect 4249 2391 4307 2397
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6270 2428 6276 2440
rect 5859 2400 6276 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 5828 2360 5856 2391
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 6730 2428 6736 2440
rect 6691 2400 6736 2428
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 8110 2428 8116 2440
rect 8071 2400 8116 2428
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 9324 2428 9352 2536
rect 9398 2524 9404 2576
rect 9456 2564 9462 2576
rect 11701 2567 11759 2573
rect 11701 2564 11713 2567
rect 9456 2536 11713 2564
rect 9456 2524 9462 2536
rect 11701 2533 11713 2536
rect 11747 2533 11759 2567
rect 11701 2527 11759 2533
rect 13722 2524 13728 2576
rect 13780 2564 13786 2576
rect 15120 2564 15148 2604
rect 15838 2592 15844 2604
rect 15896 2592 15902 2644
rect 17402 2632 17408 2644
rect 17363 2604 17408 2632
rect 17402 2592 17408 2604
rect 17460 2592 17466 2644
rect 25406 2592 25412 2644
rect 25464 2632 25470 2644
rect 29270 2632 29276 2644
rect 25464 2604 29276 2632
rect 25464 2592 25470 2604
rect 29270 2592 29276 2604
rect 29328 2592 29334 2644
rect 51994 2592 52000 2644
rect 52052 2632 52058 2644
rect 55309 2635 55367 2641
rect 55309 2632 55321 2635
rect 52052 2604 55321 2632
rect 52052 2592 52058 2604
rect 55309 2601 55321 2604
rect 55355 2601 55367 2635
rect 55309 2595 55367 2601
rect 13780 2536 15148 2564
rect 15197 2567 15255 2573
rect 13780 2524 13786 2536
rect 15197 2533 15209 2567
rect 15243 2533 15255 2567
rect 15197 2527 15255 2533
rect 16117 2567 16175 2573
rect 16117 2533 16129 2567
rect 16163 2564 16175 2567
rect 16206 2564 16212 2576
rect 16163 2536 16212 2564
rect 16163 2533 16175 2536
rect 16117 2527 16175 2533
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 14918 2496 14924 2508
rect 9631 2468 14924 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 14918 2456 14924 2468
rect 14976 2456 14982 2508
rect 15212 2496 15240 2527
rect 16206 2524 16212 2536
rect 16264 2524 16270 2576
rect 18046 2564 18052 2576
rect 18007 2536 18052 2564
rect 18046 2524 18052 2536
rect 18104 2524 18110 2576
rect 19150 2524 19156 2576
rect 19208 2564 19214 2576
rect 19245 2567 19303 2573
rect 19245 2564 19257 2567
rect 19208 2536 19257 2564
rect 19208 2524 19214 2536
rect 19245 2533 19257 2536
rect 19291 2533 19303 2567
rect 19245 2527 19303 2533
rect 20162 2524 20168 2576
rect 20220 2564 20226 2576
rect 20257 2567 20315 2573
rect 20257 2564 20269 2567
rect 20220 2536 20269 2564
rect 20220 2524 20226 2536
rect 20257 2533 20269 2536
rect 20303 2533 20315 2567
rect 20257 2527 20315 2533
rect 21085 2567 21143 2573
rect 21085 2533 21097 2567
rect 21131 2564 21143 2567
rect 22462 2564 22468 2576
rect 21131 2536 22468 2564
rect 21131 2533 21143 2536
rect 21085 2527 21143 2533
rect 22462 2524 22468 2536
rect 22520 2524 22526 2576
rect 22741 2567 22799 2573
rect 22741 2533 22753 2567
rect 22787 2564 22799 2567
rect 22922 2564 22928 2576
rect 22787 2536 22928 2564
rect 22787 2533 22799 2536
rect 22741 2527 22799 2533
rect 22922 2524 22928 2536
rect 22980 2524 22986 2576
rect 23569 2567 23627 2573
rect 23569 2533 23581 2567
rect 23615 2564 23627 2567
rect 25777 2567 25835 2573
rect 23615 2536 25452 2564
rect 23615 2533 23627 2536
rect 23569 2527 23627 2533
rect 25424 2496 25452 2536
rect 25777 2533 25789 2567
rect 25823 2564 25835 2567
rect 27246 2564 27252 2576
rect 25823 2536 27252 2564
rect 25823 2533 25835 2536
rect 25777 2527 25835 2533
rect 27246 2524 27252 2536
rect 27304 2524 27310 2576
rect 27709 2567 27767 2573
rect 27709 2533 27721 2567
rect 27755 2564 27767 2567
rect 28350 2564 28356 2576
rect 27755 2536 28356 2564
rect 27755 2533 27767 2536
rect 27709 2527 27767 2533
rect 28350 2524 28356 2536
rect 28408 2524 28414 2576
rect 34146 2524 34152 2576
rect 34204 2564 34210 2576
rect 35989 2567 36047 2573
rect 35989 2564 36001 2567
rect 34204 2536 36001 2564
rect 34204 2524 34210 2536
rect 35989 2533 36001 2536
rect 36035 2533 36047 2567
rect 35989 2527 36047 2533
rect 38010 2524 38016 2576
rect 38068 2564 38074 2576
rect 39853 2567 39911 2573
rect 39853 2564 39865 2567
rect 38068 2536 39865 2564
rect 38068 2524 38074 2536
rect 39853 2533 39865 2536
rect 39899 2533 39911 2567
rect 39853 2527 39911 2533
rect 41874 2524 41880 2576
rect 41932 2564 41938 2576
rect 43717 2567 43775 2573
rect 43717 2564 43729 2567
rect 41932 2536 43729 2564
rect 41932 2524 41938 2536
rect 43717 2533 43729 2536
rect 43763 2533 43775 2567
rect 43717 2527 43775 2533
rect 45738 2524 45744 2576
rect 45796 2564 45802 2576
rect 47581 2567 47639 2573
rect 47581 2564 47593 2567
rect 45796 2536 47593 2564
rect 45796 2524 45802 2536
rect 47581 2533 47593 2536
rect 47627 2533 47639 2567
rect 47581 2527 47639 2533
rect 49602 2524 49608 2576
rect 49660 2564 49666 2576
rect 51445 2567 51503 2573
rect 51445 2564 51457 2567
rect 49660 2536 51457 2564
rect 49660 2524 49666 2536
rect 51445 2533 51457 2536
rect 51491 2533 51503 2567
rect 51445 2527 51503 2533
rect 54021 2567 54079 2573
rect 54021 2533 54033 2567
rect 54067 2533 54079 2567
rect 54021 2527 54079 2533
rect 26234 2496 26240 2508
rect 15212 2468 25268 2496
rect 25424 2468 26240 2496
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 9324 2400 11529 2428
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 11698 2388 11704 2440
rect 11756 2428 11762 2440
rect 12253 2431 12311 2437
rect 12253 2428 12265 2431
rect 11756 2400 12265 2428
rect 11756 2388 11762 2400
rect 12253 2397 12265 2400
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2397 13323 2431
rect 13265 2391 13323 2397
rect 7742 2360 7748 2372
rect 2648 2332 5856 2360
rect 6380 2332 7748 2360
rect 2648 2320 2654 2332
rect 1762 2292 1768 2304
rect 1723 2264 1768 2292
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 4433 2295 4491 2301
rect 4433 2261 4445 2295
rect 4479 2292 4491 2295
rect 6380 2292 6408 2332
rect 7742 2320 7748 2332
rect 7800 2320 7806 2372
rect 8478 2320 8484 2372
rect 8536 2360 8542 2372
rect 10137 2363 10195 2369
rect 10137 2360 10149 2363
rect 8536 2332 10149 2360
rect 8536 2320 8542 2332
rect 10137 2329 10149 2332
rect 10183 2329 10195 2363
rect 10137 2323 10195 2329
rect 10318 2320 10324 2372
rect 10376 2360 10382 2372
rect 13280 2360 13308 2391
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 14369 2431 14427 2437
rect 14369 2428 14381 2431
rect 14056 2400 14381 2428
rect 14056 2388 14062 2400
rect 14369 2397 14381 2400
rect 14415 2428 14427 2431
rect 14550 2428 14556 2440
rect 14415 2400 14556 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 15381 2431 15439 2437
rect 15381 2397 15393 2431
rect 15427 2428 15439 2431
rect 15470 2428 15476 2440
rect 15427 2400 15476 2428
rect 15427 2397 15439 2400
rect 15381 2391 15439 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 15838 2388 15844 2440
rect 15896 2428 15902 2440
rect 15933 2431 15991 2437
rect 15933 2428 15945 2431
rect 15896 2400 15945 2428
rect 15896 2388 15902 2400
rect 15933 2397 15945 2400
rect 15979 2397 15991 2431
rect 15933 2391 15991 2397
rect 16853 2431 16911 2437
rect 16853 2397 16865 2431
rect 16899 2428 16911 2431
rect 17862 2428 17868 2440
rect 16899 2400 17868 2428
rect 16899 2397 16911 2400
rect 16853 2391 16911 2397
rect 17862 2388 17868 2400
rect 17920 2388 17926 2440
rect 18233 2431 18291 2437
rect 18233 2397 18245 2431
rect 18279 2428 18291 2431
rect 19518 2428 19524 2440
rect 18279 2400 19524 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 19518 2388 19524 2400
rect 19576 2388 19582 2440
rect 21266 2428 21272 2440
rect 21227 2400 21272 2428
rect 21266 2388 21272 2400
rect 21324 2388 21330 2440
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2428 22247 2431
rect 22370 2428 22376 2440
rect 22235 2400 22376 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 22370 2388 22376 2400
rect 22428 2388 22434 2440
rect 22925 2431 22983 2437
rect 22925 2397 22937 2431
rect 22971 2428 22983 2431
rect 23014 2428 23020 2440
rect 22971 2400 23020 2428
rect 22971 2397 22983 2400
rect 22925 2391 22983 2397
rect 23014 2388 23020 2400
rect 23072 2388 23078 2440
rect 23290 2388 23296 2440
rect 23348 2428 23354 2440
rect 23385 2431 23443 2437
rect 23385 2428 23397 2431
rect 23348 2400 23397 2428
rect 23348 2388 23354 2400
rect 23385 2397 23397 2400
rect 23431 2428 23443 2431
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 23431 2400 24409 2428
rect 23431 2397 23443 2400
rect 23385 2391 23443 2397
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 24397 2391 24455 2397
rect 25133 2431 25191 2437
rect 25133 2397 25145 2431
rect 25179 2397 25191 2431
rect 25240 2428 25268 2468
rect 26234 2456 26240 2468
rect 26292 2456 26298 2508
rect 26510 2496 26516 2508
rect 26344 2468 26516 2496
rect 26344 2428 26372 2468
rect 26510 2456 26516 2468
rect 26568 2456 26574 2508
rect 31938 2456 31944 2508
rect 31996 2496 32002 2508
rect 32769 2499 32827 2505
rect 32769 2496 32781 2499
rect 31996 2468 32781 2496
rect 31996 2456 32002 2468
rect 32769 2465 32781 2468
rect 32815 2465 32827 2499
rect 32769 2459 32827 2465
rect 33042 2456 33048 2508
rect 33100 2496 33106 2508
rect 34701 2499 34759 2505
rect 34701 2496 34713 2499
rect 33100 2468 34713 2496
rect 33100 2456 33106 2468
rect 34701 2465 34713 2468
rect 34747 2465 34759 2499
rect 34701 2459 34759 2465
rect 35526 2456 35532 2508
rect 35584 2496 35590 2508
rect 37277 2499 37335 2505
rect 37277 2496 37289 2499
rect 35584 2468 37289 2496
rect 35584 2456 35590 2468
rect 37277 2465 37289 2468
rect 37323 2465 37335 2499
rect 37277 2459 37335 2465
rect 38838 2456 38844 2508
rect 38896 2496 38902 2508
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 38896 2468 40509 2496
rect 38896 2456 38902 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 40497 2459 40555 2465
rect 40770 2456 40776 2508
rect 40828 2496 40834 2508
rect 42429 2499 42487 2505
rect 42429 2496 42441 2499
rect 40828 2468 42441 2496
rect 40828 2456 40834 2468
rect 42429 2465 42441 2468
rect 42475 2465 42487 2499
rect 42429 2459 42487 2465
rect 43254 2456 43260 2508
rect 43312 2496 43318 2508
rect 45005 2499 45063 2505
rect 45005 2496 45017 2499
rect 43312 2468 45017 2496
rect 43312 2456 43318 2468
rect 45005 2465 45017 2468
rect 45051 2465 45063 2499
rect 45005 2459 45063 2465
rect 46566 2456 46572 2508
rect 46624 2496 46630 2508
rect 48225 2499 48283 2505
rect 48225 2496 48237 2499
rect 46624 2468 48237 2496
rect 46624 2456 46630 2468
rect 48225 2465 48237 2468
rect 48271 2465 48283 2499
rect 48225 2459 48283 2465
rect 48498 2456 48504 2508
rect 48556 2496 48562 2508
rect 50157 2499 50215 2505
rect 50157 2496 50169 2499
rect 48556 2468 50169 2496
rect 48556 2456 48562 2468
rect 50157 2465 50169 2468
rect 50203 2465 50215 2499
rect 52733 2499 52791 2505
rect 52733 2496 52745 2499
rect 50157 2459 50215 2465
rect 51046 2468 52745 2496
rect 25240 2400 26372 2428
rect 26421 2431 26479 2437
rect 25133 2391 25191 2397
rect 26421 2397 26433 2431
rect 26467 2428 26479 2431
rect 27522 2428 27528 2440
rect 26467 2400 27528 2428
rect 26467 2397 26479 2400
rect 26421 2391 26479 2397
rect 10376 2332 13308 2360
rect 15488 2360 15516 2388
rect 17218 2360 17224 2372
rect 15488 2332 17224 2360
rect 10376 2320 10382 2332
rect 4479 2264 6408 2292
rect 6641 2295 6699 2301
rect 4479 2261 4491 2264
rect 4433 2255 4491 2261
rect 6641 2261 6653 2295
rect 6687 2292 6699 2295
rect 6730 2292 6736 2304
rect 6687 2264 6736 2292
rect 6687 2261 6699 2264
rect 6641 2255 6699 2261
rect 6730 2252 6736 2264
rect 6788 2252 6794 2304
rect 13280 2292 13308 2332
rect 17218 2320 17224 2332
rect 17276 2320 17282 2372
rect 17497 2363 17555 2369
rect 17497 2329 17509 2363
rect 17543 2329 17555 2363
rect 17497 2323 17555 2329
rect 19429 2363 19487 2369
rect 19429 2329 19441 2363
rect 19475 2360 19487 2363
rect 20254 2360 20260 2372
rect 19475 2332 20260 2360
rect 19475 2329 19487 2332
rect 19429 2323 19487 2329
rect 16022 2292 16028 2304
rect 13280 2264 16028 2292
rect 16022 2252 16028 2264
rect 16080 2252 16086 2304
rect 17512 2292 17540 2323
rect 20254 2320 20260 2332
rect 20312 2320 20318 2372
rect 20441 2363 20499 2369
rect 20441 2329 20453 2363
rect 20487 2360 20499 2363
rect 21542 2360 21548 2372
rect 20487 2332 21548 2360
rect 20487 2329 20499 2332
rect 20441 2323 20499 2329
rect 21542 2320 21548 2332
rect 21600 2320 21606 2372
rect 25148 2360 25176 2391
rect 27522 2388 27528 2400
rect 27580 2388 27586 2440
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 28902 2428 28908 2440
rect 28399 2400 28908 2428
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 28902 2388 28908 2400
rect 28960 2388 28966 2440
rect 28997 2431 29055 2437
rect 28997 2397 29009 2431
rect 29043 2428 29055 2431
rect 29454 2428 29460 2440
rect 29043 2400 29460 2428
rect 29043 2397 29055 2400
rect 28997 2391 29055 2397
rect 29454 2388 29460 2400
rect 29512 2388 29518 2440
rect 30101 2431 30159 2437
rect 30101 2397 30113 2431
rect 30147 2428 30159 2431
rect 30282 2428 30288 2440
rect 30147 2400 30288 2428
rect 30147 2397 30159 2400
rect 30101 2391 30159 2397
rect 30282 2388 30288 2400
rect 30340 2388 30346 2440
rect 30745 2431 30803 2437
rect 30745 2397 30757 2431
rect 30791 2428 30803 2431
rect 30834 2428 30840 2440
rect 30791 2400 30840 2428
rect 30791 2397 30803 2400
rect 30745 2391 30803 2397
rect 30834 2388 30840 2400
rect 30892 2388 30898 2440
rect 31110 2388 31116 2440
rect 31168 2428 31174 2440
rect 31205 2431 31263 2437
rect 31205 2428 31217 2431
rect 31168 2400 31217 2428
rect 31168 2388 31174 2400
rect 31205 2397 31217 2400
rect 31251 2397 31263 2431
rect 31205 2391 31263 2397
rect 31386 2388 31392 2440
rect 31444 2428 31450 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31444 2400 32137 2428
rect 31444 2388 31450 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 32490 2388 32496 2440
rect 32548 2428 32554 2440
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 32548 2400 33425 2428
rect 32548 2388 32554 2400
rect 33413 2397 33425 2400
rect 33459 2397 33471 2431
rect 33413 2391 33471 2397
rect 33594 2388 33600 2440
rect 33652 2428 33658 2440
rect 35345 2431 35403 2437
rect 35345 2428 35357 2431
rect 33652 2400 35357 2428
rect 33652 2388 33658 2400
rect 35345 2397 35357 2400
rect 35391 2397 35403 2431
rect 35345 2391 35403 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 37921 2431 37979 2437
rect 37921 2428 37933 2431
rect 36136 2400 37933 2428
rect 36136 2388 36142 2400
rect 37921 2397 37933 2400
rect 37967 2397 37979 2431
rect 37921 2391 37979 2397
rect 38565 2431 38623 2437
rect 38565 2397 38577 2431
rect 38611 2397 38623 2431
rect 38565 2391 38623 2397
rect 26694 2360 26700 2372
rect 25148 2332 26700 2360
rect 26694 2320 26700 2332
rect 26752 2320 26758 2372
rect 36906 2320 36912 2372
rect 36964 2360 36970 2372
rect 38580 2360 38608 2391
rect 39390 2388 39396 2440
rect 39448 2428 39454 2440
rect 41141 2431 41199 2437
rect 41141 2428 41153 2431
rect 39448 2400 41153 2428
rect 39448 2388 39454 2400
rect 41141 2397 41153 2400
rect 41187 2397 41199 2431
rect 41141 2391 41199 2397
rect 41322 2388 41328 2440
rect 41380 2428 41386 2440
rect 43073 2431 43131 2437
rect 43073 2428 43085 2431
rect 41380 2400 43085 2428
rect 41380 2388 41386 2400
rect 43073 2397 43085 2400
rect 43119 2397 43131 2431
rect 43073 2391 43131 2397
rect 43806 2388 43812 2440
rect 43864 2428 43870 2440
rect 45649 2431 45707 2437
rect 45649 2428 45661 2431
rect 43864 2400 45661 2428
rect 43864 2388 43870 2400
rect 45649 2397 45661 2400
rect 45695 2397 45707 2431
rect 45649 2391 45707 2397
rect 46293 2431 46351 2437
rect 46293 2397 46305 2431
rect 46339 2397 46351 2431
rect 46293 2391 46351 2397
rect 36964 2332 38608 2360
rect 36964 2320 36970 2332
rect 44634 2320 44640 2372
rect 44692 2360 44698 2372
rect 46308 2360 46336 2391
rect 47118 2388 47124 2440
rect 47176 2428 47182 2440
rect 48869 2431 48927 2437
rect 48869 2428 48881 2431
rect 47176 2400 48881 2428
rect 47176 2388 47182 2400
rect 48869 2397 48881 2400
rect 48915 2397 48927 2431
rect 48869 2391 48927 2397
rect 49050 2388 49056 2440
rect 49108 2428 49114 2440
rect 50801 2431 50859 2437
rect 50801 2428 50813 2431
rect 49108 2400 50813 2428
rect 49108 2388 49114 2400
rect 50801 2397 50813 2400
rect 50847 2397 50859 2431
rect 50801 2391 50859 2397
rect 50890 2388 50896 2440
rect 50948 2428 50954 2440
rect 51046 2428 51074 2468
rect 52733 2465 52745 2468
rect 52779 2465 52791 2499
rect 54036 2496 54064 2527
rect 57882 2496 57888 2508
rect 54036 2468 54156 2496
rect 57843 2468 57888 2496
rect 52733 2459 52791 2465
rect 50948 2400 51074 2428
rect 50948 2388 50954 2400
rect 52546 2388 52552 2440
rect 52604 2428 52610 2440
rect 53377 2431 53435 2437
rect 53377 2428 53389 2431
rect 52604 2400 53389 2428
rect 52604 2388 52610 2400
rect 53377 2397 53389 2400
rect 53423 2397 53435 2431
rect 53377 2391 53435 2397
rect 44692 2332 46336 2360
rect 44692 2320 44698 2332
rect 18506 2292 18512 2304
rect 17512 2264 18512 2292
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 22002 2292 22008 2304
rect 21963 2264 22008 2292
rect 22002 2252 22008 2264
rect 22060 2252 22066 2304
rect 23014 2252 23020 2304
rect 23072 2292 23078 2304
rect 26973 2295 27031 2301
rect 26973 2292 26985 2295
rect 23072 2264 26985 2292
rect 23072 2252 23078 2264
rect 26973 2261 26985 2264
rect 27019 2261 27031 2295
rect 26973 2255 27031 2261
rect 51258 2252 51264 2304
rect 51316 2292 51322 2304
rect 54128 2292 54156 2468
rect 57882 2456 57888 2468
rect 57940 2456 57946 2508
rect 55950 2428 55956 2440
rect 55911 2400 55956 2428
rect 55950 2388 55956 2400
rect 56008 2388 56014 2440
rect 56594 2428 56600 2440
rect 56555 2400 56600 2428
rect 56594 2388 56600 2400
rect 56652 2388 56658 2440
rect 51316 2264 54156 2292
rect 51316 2252 51322 2264
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 7190 2048 7196 2100
rect 7248 2088 7254 2100
rect 10318 2088 10324 2100
rect 7248 2060 10324 2088
rect 7248 2048 7254 2060
rect 10318 2048 10324 2060
rect 10376 2048 10382 2100
rect 10686 2048 10692 2100
rect 10744 2088 10750 2100
rect 13998 2088 14004 2100
rect 10744 2060 14004 2088
rect 10744 2048 10750 2060
rect 13998 2048 14004 2060
rect 14056 2048 14062 2100
rect 25406 2088 25412 2100
rect 14200 2060 25412 2088
rect 9490 2020 9496 2032
rect 2746 1992 9496 2020
rect 1762 1912 1768 1964
rect 1820 1952 1826 1964
rect 2746 1952 2774 1992
rect 9490 1980 9496 1992
rect 9548 1980 9554 2032
rect 10410 1980 10416 2032
rect 10468 2020 10474 2032
rect 14200 2020 14228 2060
rect 25406 2048 25412 2060
rect 25464 2048 25470 2100
rect 26234 2048 26240 2100
rect 26292 2088 26298 2100
rect 34606 2088 34612 2100
rect 26292 2060 34612 2088
rect 26292 2048 26298 2060
rect 34606 2048 34612 2060
rect 34664 2048 34670 2100
rect 52362 2048 52368 2100
rect 52420 2088 52426 2100
rect 55950 2088 55956 2100
rect 52420 2060 55956 2088
rect 52420 2048 52426 2060
rect 55950 2048 55956 2060
rect 56008 2048 56014 2100
rect 10468 1992 14228 2020
rect 10468 1980 10474 1992
rect 14550 1980 14556 2032
rect 14608 2020 14614 2032
rect 16390 2020 16396 2032
rect 14608 1992 16396 2020
rect 14608 1980 14614 1992
rect 16390 1980 16396 1992
rect 16448 1980 16454 2032
rect 22002 1980 22008 2032
rect 22060 2020 22066 2032
rect 45554 2020 45560 2032
rect 22060 1992 45560 2020
rect 22060 1980 22066 1992
rect 45554 1980 45560 1992
rect 45612 1980 45618 2032
rect 53558 1980 53564 2032
rect 53616 2020 53622 2032
rect 57882 2020 57888 2032
rect 53616 1992 57888 2020
rect 53616 1980 53622 1992
rect 57882 1980 57888 1992
rect 57940 1980 57946 2032
rect 1820 1924 2774 1952
rect 1820 1912 1826 1924
rect 6730 1912 6736 1964
rect 6788 1952 6794 1964
rect 28810 1952 28816 1964
rect 6788 1924 28816 1952
rect 6788 1912 6794 1924
rect 28810 1912 28816 1924
rect 28868 1912 28874 1964
rect 5442 1844 5448 1896
rect 5500 1884 5506 1896
rect 10686 1884 10692 1896
rect 5500 1856 10692 1884
rect 5500 1844 5506 1856
rect 10686 1844 10692 1856
rect 10744 1844 10750 1896
rect 15838 1844 15844 1896
rect 15896 1884 15902 1896
rect 18046 1884 18052 1896
rect 15896 1856 18052 1884
rect 15896 1844 15902 1856
rect 18046 1844 18052 1856
rect 18104 1844 18110 1896
rect 1578 1708 1584 1760
rect 1636 1748 1642 1760
rect 1636 1720 2774 1748
rect 1636 1708 1642 1720
rect 2746 1612 2774 1720
rect 7190 1708 7196 1760
rect 7248 1748 7254 1760
rect 8110 1748 8116 1760
rect 7248 1720 8116 1748
rect 7248 1708 7254 1720
rect 8110 1708 8116 1720
rect 8168 1708 8174 1760
rect 18506 1708 18512 1760
rect 18564 1748 18570 1760
rect 18874 1748 18880 1760
rect 18564 1720 18880 1748
rect 18564 1708 18570 1720
rect 18874 1708 18880 1720
rect 18932 1708 18938 1760
rect 21082 1640 21088 1692
rect 21140 1680 21146 1692
rect 21542 1680 21548 1692
rect 21140 1652 21548 1680
rect 21140 1640 21146 1652
rect 21542 1640 21548 1652
rect 21600 1640 21606 1692
rect 8110 1612 8116 1624
rect 2746 1584 8116 1612
rect 8110 1572 8116 1584
rect 8168 1572 8174 1624
rect 20254 1572 20260 1624
rect 20312 1572 20318 1624
rect 5994 1504 6000 1556
rect 6052 1544 6058 1556
rect 6362 1544 6368 1556
rect 6052 1516 6368 1544
rect 6052 1504 6058 1516
rect 6362 1504 6368 1516
rect 6420 1504 6426 1556
rect 20272 1488 20300 1572
rect 20346 1504 20352 1556
rect 20404 1504 20410 1556
rect 20254 1436 20260 1488
rect 20312 1436 20318 1488
rect 2958 1368 2964 1420
rect 3016 1408 3022 1420
rect 3016 1380 6316 1408
rect 3016 1368 3022 1380
rect 6288 1216 6316 1380
rect 8846 1368 8852 1420
rect 8904 1408 8910 1420
rect 10594 1408 10600 1420
rect 8904 1380 10600 1408
rect 8904 1368 8910 1380
rect 10594 1368 10600 1380
rect 10652 1368 10658 1420
rect 19334 1300 19340 1352
rect 19392 1340 19398 1352
rect 19794 1340 19800 1352
rect 19392 1312 19800 1340
rect 19392 1300 19398 1312
rect 19794 1300 19800 1312
rect 19852 1300 19858 1352
rect 19978 1300 19984 1352
rect 20036 1340 20042 1352
rect 20364 1340 20392 1504
rect 52730 1368 52736 1420
rect 52788 1408 52794 1420
rect 53006 1408 53012 1420
rect 52788 1380 53012 1408
rect 52788 1368 52794 1380
rect 53006 1368 53012 1380
rect 53064 1368 53070 1420
rect 56594 1408 56600 1420
rect 53116 1380 56600 1408
rect 20036 1312 20392 1340
rect 20036 1300 20042 1312
rect 19426 1232 19432 1284
rect 19484 1232 19490 1284
rect 6270 1164 6276 1216
rect 6328 1164 6334 1216
rect 19444 932 19472 1232
rect 52546 1136 52552 1148
rect 51000 1108 52552 1136
rect 51000 944 51028 1108
rect 52546 1096 52552 1108
rect 52604 1096 52610 1148
rect 19518 932 19524 944
rect 19444 904 19524 932
rect 19518 892 19524 904
rect 19576 892 19582 944
rect 50982 892 50988 944
rect 51040 892 51046 944
rect 52546 892 52552 944
rect 52604 892 52610 944
rect 52914 892 52920 944
rect 52972 932 52978 944
rect 53116 932 53144 1380
rect 56594 1368 56600 1380
rect 56652 1368 56658 1420
rect 52972 904 53144 932
rect 52972 892 52978 904
rect 52564 864 52592 892
rect 54754 864 54760 876
rect 52564 836 54760 864
rect 54754 824 54760 836
rect 54812 824 54818 876
<< via1 >>
rect 5264 57740 5316 57792
rect 18328 57740 18380 57792
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 1768 57536 1820 57588
rect 3332 57536 3384 57588
rect 4896 57536 4948 57588
rect 6460 57536 6512 57588
rect 8024 57536 8076 57588
rect 9680 57536 9732 57588
rect 11152 57536 11204 57588
rect 12716 57536 12768 57588
rect 14280 57536 14332 57588
rect 15844 57536 15896 57588
rect 17408 57536 17460 57588
rect 19340 57536 19392 57588
rect 20720 57536 20772 57588
rect 22100 57536 22152 57588
rect 23664 57536 23716 57588
rect 25228 57536 25280 57588
rect 26792 57536 26844 57588
rect 28356 57536 28408 57588
rect 29920 57536 29972 57588
rect 31484 57536 31536 57588
rect 33140 57536 33192 57588
rect 34612 57536 34664 57588
rect 36176 57536 36228 57588
rect 37740 57536 37792 57588
rect 39304 57536 39356 57588
rect 40868 57536 40920 57588
rect 42432 57536 42484 57588
rect 44180 57536 44232 57588
rect 45560 57536 45612 57588
rect 47124 57536 47176 57588
rect 2688 57400 2740 57452
rect 4068 57443 4120 57452
rect 4068 57409 4077 57443
rect 4077 57409 4111 57443
rect 4111 57409 4120 57443
rect 4068 57400 4120 57409
rect 5264 57443 5316 57452
rect 5264 57409 5273 57443
rect 5273 57409 5307 57443
rect 5307 57409 5316 57443
rect 5264 57400 5316 57409
rect 19156 57468 19208 57520
rect 11796 57443 11848 57452
rect 2688 57239 2740 57248
rect 2688 57205 2697 57239
rect 2697 57205 2731 57239
rect 2731 57205 2740 57239
rect 2688 57196 2740 57205
rect 11796 57409 11805 57443
rect 11805 57409 11839 57443
rect 11839 57409 11848 57443
rect 11796 57400 11848 57409
rect 13084 57443 13136 57452
rect 13084 57409 13093 57443
rect 13093 57409 13127 57443
rect 13127 57409 13136 57443
rect 13084 57400 13136 57409
rect 15936 57400 15988 57452
rect 16948 57443 17000 57452
rect 16948 57409 16957 57443
rect 16957 57409 16991 57443
rect 16991 57409 17000 57443
rect 16948 57400 17000 57409
rect 17500 57443 17552 57452
rect 17500 57409 17509 57443
rect 17509 57409 17543 57443
rect 17543 57409 17552 57443
rect 17500 57400 17552 57409
rect 19248 57443 19300 57452
rect 19248 57409 19257 57443
rect 19257 57409 19291 57443
rect 19291 57409 19300 57443
rect 19248 57400 19300 57409
rect 19340 57400 19392 57452
rect 22192 57443 22244 57452
rect 22192 57409 22201 57443
rect 22201 57409 22235 57443
rect 22235 57409 22244 57443
rect 22192 57400 22244 57409
rect 24400 57443 24452 57452
rect 24400 57409 24409 57443
rect 24409 57409 24443 57443
rect 24443 57409 24452 57443
rect 24400 57400 24452 57409
rect 25320 57443 25372 57452
rect 25320 57409 25329 57443
rect 25329 57409 25363 57443
rect 25363 57409 25372 57443
rect 25320 57400 25372 57409
rect 26976 57443 27028 57452
rect 26976 57409 26985 57443
rect 26985 57409 27019 57443
rect 27019 57409 27028 57443
rect 26976 57400 27028 57409
rect 28448 57443 28500 57452
rect 28448 57409 28457 57443
rect 28457 57409 28491 57443
rect 28491 57409 28500 57443
rect 28448 57400 28500 57409
rect 30012 57443 30064 57452
rect 30012 57409 30021 57443
rect 30021 57409 30055 57443
rect 30055 57409 30064 57443
rect 30012 57400 30064 57409
rect 27620 57332 27672 57384
rect 30380 57332 30432 57384
rect 33232 57400 33284 57452
rect 34796 57400 34848 57452
rect 37832 57443 37884 57452
rect 37832 57409 37841 57443
rect 37841 57409 37875 57443
rect 37875 57409 37884 57443
rect 37832 57400 37884 57409
rect 37924 57400 37976 57452
rect 40960 57443 41012 57452
rect 40960 57409 40969 57443
rect 40969 57409 41003 57443
rect 41003 57409 41012 57443
rect 40960 57400 41012 57409
rect 42340 57400 42392 57452
rect 44088 57443 44140 57452
rect 44088 57409 44097 57443
rect 44097 57409 44131 57443
rect 44131 57409 44140 57443
rect 44088 57400 44140 57409
rect 45652 57443 45704 57452
rect 45652 57409 45661 57443
rect 45661 57409 45695 57443
rect 45695 57409 45704 57443
rect 45652 57400 45704 57409
rect 47584 57443 47636 57452
rect 47584 57409 47593 57443
rect 47593 57409 47627 57443
rect 47627 57409 47636 57443
rect 47584 57400 47636 57409
rect 48688 57400 48740 57452
rect 50160 57400 50212 57452
rect 51816 57400 51868 57452
rect 53380 57400 53432 57452
rect 56600 57443 56652 57452
rect 56600 57409 56609 57443
rect 56609 57409 56643 57443
rect 56643 57409 56652 57443
rect 56600 57400 56652 57409
rect 58072 57400 58124 57452
rect 54944 57332 54996 57384
rect 18420 57264 18472 57316
rect 17868 57196 17920 57248
rect 18512 57196 18564 57248
rect 20076 57239 20128 57248
rect 20076 57205 20085 57239
rect 20085 57205 20119 57239
rect 20119 57205 20128 57239
rect 20076 57196 20128 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 18328 57035 18380 57044
rect 18328 57001 18337 57035
rect 18337 57001 18371 57035
rect 18371 57001 18380 57035
rect 18328 56992 18380 57001
rect 19156 56992 19208 57044
rect 57520 57035 57572 57044
rect 57520 57001 57529 57035
rect 57529 57001 57563 57035
rect 57563 57001 57572 57035
rect 57520 56992 57572 57001
rect 11796 56924 11848 56976
rect 19432 56924 19484 56976
rect 18512 56831 18564 56840
rect 18512 56797 18521 56831
rect 18521 56797 18555 56831
rect 18555 56797 18564 56831
rect 18512 56788 18564 56797
rect 20076 56788 20128 56840
rect 18052 56652 18104 56704
rect 19984 56652 20036 56704
rect 20720 56695 20772 56704
rect 20720 56661 20729 56695
rect 20729 56661 20763 56695
rect 20763 56661 20772 56695
rect 20720 56652 20772 56661
rect 22284 56695 22336 56704
rect 22284 56661 22293 56695
rect 22293 56661 22327 56695
rect 22327 56661 22336 56695
rect 22284 56652 22336 56661
rect 25136 56652 25188 56704
rect 57888 56788 57940 56840
rect 30012 56720 30064 56772
rect 26608 56695 26660 56704
rect 26608 56661 26617 56695
rect 26617 56661 26651 56695
rect 26651 56661 26660 56695
rect 26608 56652 26660 56661
rect 42340 56695 42392 56704
rect 42340 56661 42349 56695
rect 42349 56661 42383 56695
rect 42383 56661 42392 56695
rect 42340 56652 42392 56661
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 13084 56448 13136 56500
rect 15936 56491 15988 56500
rect 15936 56457 15945 56491
rect 15945 56457 15979 56491
rect 15979 56457 15988 56491
rect 15936 56448 15988 56457
rect 17500 56448 17552 56500
rect 17868 56491 17920 56500
rect 17868 56457 17877 56491
rect 17877 56457 17911 56491
rect 17911 56457 17920 56491
rect 17868 56448 17920 56457
rect 18420 56448 18472 56500
rect 19340 56491 19392 56500
rect 19340 56457 19349 56491
rect 19349 56457 19383 56491
rect 19383 56457 19392 56491
rect 19340 56448 19392 56457
rect 13728 56355 13780 56364
rect 13728 56321 13737 56355
rect 13737 56321 13771 56355
rect 13771 56321 13780 56355
rect 13728 56312 13780 56321
rect 16212 56312 16264 56364
rect 17408 56312 17460 56364
rect 18052 56355 18104 56364
rect 18052 56321 18061 56355
rect 18061 56321 18095 56355
rect 18095 56321 18104 56355
rect 18880 56380 18932 56432
rect 18696 56355 18748 56364
rect 18052 56312 18104 56321
rect 18696 56321 18705 56355
rect 18705 56321 18739 56355
rect 18739 56321 18748 56355
rect 18696 56312 18748 56321
rect 18972 56312 19024 56364
rect 2688 56244 2740 56296
rect 22192 56448 22244 56500
rect 24400 56448 24452 56500
rect 26976 56448 27028 56500
rect 27620 56448 27672 56500
rect 30380 56448 30432 56500
rect 33232 56448 33284 56500
rect 34796 56448 34848 56500
rect 37924 56448 37976 56500
rect 45652 56448 45704 56500
rect 47584 56448 47636 56500
rect 19984 56355 20036 56364
rect 19984 56321 19993 56355
rect 19993 56321 20027 56355
rect 20027 56321 20036 56355
rect 19984 56312 20036 56321
rect 20536 56312 20588 56364
rect 20720 56312 20772 56364
rect 21088 56355 21140 56364
rect 21088 56321 21097 56355
rect 21097 56321 21131 56355
rect 21131 56321 21140 56355
rect 21088 56312 21140 56321
rect 21640 56312 21692 56364
rect 22284 56312 22336 56364
rect 22560 56312 22612 56364
rect 23940 56355 23992 56364
rect 23940 56321 23949 56355
rect 23949 56321 23983 56355
rect 23983 56321 23992 56355
rect 23940 56312 23992 56321
rect 24952 56355 25004 56364
rect 24952 56321 24961 56355
rect 24961 56321 24995 56355
rect 24995 56321 25004 56355
rect 24952 56312 25004 56321
rect 25596 56355 25648 56364
rect 25596 56321 25605 56355
rect 25605 56321 25639 56355
rect 25639 56321 25648 56355
rect 25596 56312 25648 56321
rect 26608 56312 26660 56364
rect 27160 56355 27212 56364
rect 27160 56321 27169 56355
rect 27169 56321 27203 56355
rect 27203 56321 27212 56355
rect 27160 56312 27212 56321
rect 29644 56355 29696 56364
rect 29644 56321 29653 56355
rect 29653 56321 29687 56355
rect 29687 56321 29696 56355
rect 29644 56312 29696 56321
rect 42340 56380 42392 56432
rect 31668 56312 31720 56364
rect 32128 56355 32180 56364
rect 32128 56321 32137 56355
rect 32137 56321 32171 56355
rect 32171 56321 32180 56355
rect 32128 56312 32180 56321
rect 33968 56355 34020 56364
rect 33968 56321 33977 56355
rect 33977 56321 34011 56355
rect 34011 56321 34020 56355
rect 33968 56312 34020 56321
rect 35808 56355 35860 56364
rect 35808 56321 35817 56355
rect 35817 56321 35851 56355
rect 35851 56321 35860 56355
rect 35808 56312 35860 56321
rect 4068 56176 4120 56228
rect 25320 56176 25372 56228
rect 40960 56176 41012 56228
rect 13728 56108 13780 56160
rect 18788 56108 18840 56160
rect 25136 56151 25188 56160
rect 25136 56117 25145 56151
rect 25145 56117 25179 56151
rect 25179 56117 25188 56151
rect 25136 56108 25188 56117
rect 44088 56176 44140 56228
rect 42064 56108 42116 56160
rect 45560 56355 45612 56364
rect 45560 56321 45569 56355
rect 45569 56321 45603 56355
rect 45603 56321 45612 56355
rect 45560 56312 45612 56321
rect 58440 56312 58492 56364
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 16948 55904 17000 55956
rect 19248 55904 19300 55956
rect 19432 55904 19484 55956
rect 25136 55904 25188 55956
rect 37832 55904 37884 55956
rect 28448 55836 28500 55888
rect 17316 55768 17368 55820
rect 21088 55768 21140 55820
rect 17132 55700 17184 55752
rect 26332 55700 26384 55752
rect 16212 55607 16264 55616
rect 16212 55573 16221 55607
rect 16221 55573 16255 55607
rect 16255 55573 16264 55607
rect 16212 55564 16264 55573
rect 18052 55607 18104 55616
rect 18052 55573 18061 55607
rect 18061 55573 18095 55607
rect 18095 55573 18104 55607
rect 18052 55564 18104 55573
rect 20352 55607 20404 55616
rect 20352 55573 20361 55607
rect 20361 55573 20395 55607
rect 20395 55573 20404 55607
rect 20352 55564 20404 55573
rect 22560 55607 22612 55616
rect 22560 55573 22569 55607
rect 22569 55573 22603 55607
rect 22603 55573 22612 55607
rect 22560 55564 22612 55573
rect 24952 55564 25004 55616
rect 25596 55564 25648 55616
rect 26148 55564 26200 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 18696 55360 18748 55412
rect 19156 55360 19208 55412
rect 17132 55335 17184 55344
rect 17132 55301 17141 55335
rect 17141 55301 17175 55335
rect 17175 55301 17184 55335
rect 17132 55292 17184 55301
rect 18972 55335 19024 55344
rect 18972 55301 18981 55335
rect 18981 55301 19015 55335
rect 19015 55301 19024 55335
rect 18972 55292 19024 55301
rect 58164 55131 58216 55140
rect 58164 55097 58173 55131
rect 58173 55097 58207 55131
rect 58207 55097 58216 55131
rect 58164 55088 58216 55097
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 57888 53932 57940 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 57888 52436 57940 52488
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 58164 51391 58216 51400
rect 58164 51357 58173 51391
rect 58173 51357 58207 51391
rect 58207 51357 58216 51391
rect 58164 51348 58216 51357
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 58164 49759 58216 49768
rect 58164 49725 58173 49759
rect 58173 49725 58207 49759
rect 58207 49725 58216 49759
rect 58164 49716 58216 49725
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 58164 48535 58216 48544
rect 58164 48501 58173 48535
rect 58173 48501 58207 48535
rect 58207 48501 58216 48535
rect 58164 48492 58216 48501
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 15292 47540 15344 47592
rect 33968 47540 34020 47592
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 58164 47039 58216 47048
rect 58164 47005 58173 47039
rect 58173 47005 58207 47039
rect 58207 47005 58216 47039
rect 58164 46996 58216 47005
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 58164 45951 58216 45960
rect 58164 45917 58173 45951
rect 58173 45917 58207 45951
rect 58207 45917 58216 45951
rect 58164 45908 58216 45917
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 58164 44251 58216 44260
rect 58164 44217 58173 44251
rect 58173 44217 58207 44251
rect 58207 44217 58216 44251
rect 58164 44208 58216 44217
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 58164 43095 58216 43104
rect 58164 43061 58173 43095
rect 58173 43061 58207 43095
rect 58207 43061 58216 43095
rect 58164 43052 58216 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 12808 42236 12860 42288
rect 13820 42168 13872 42220
rect 14924 42211 14976 42220
rect 14924 42177 14933 42211
rect 14933 42177 14967 42211
rect 14967 42177 14976 42211
rect 14924 42168 14976 42177
rect 16672 42168 16724 42220
rect 13360 41964 13412 42016
rect 15568 41964 15620 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 12164 41488 12216 41540
rect 13360 41599 13412 41608
rect 13360 41565 13369 41599
rect 13369 41565 13403 41599
rect 13403 41565 13412 41599
rect 13360 41556 13412 41565
rect 13544 41599 13596 41608
rect 13544 41565 13553 41599
rect 13553 41565 13587 41599
rect 13587 41565 13596 41599
rect 13544 41556 13596 41565
rect 12532 41420 12584 41472
rect 12624 41420 12676 41472
rect 13636 41488 13688 41540
rect 13820 41556 13872 41608
rect 14924 41556 14976 41608
rect 15384 41556 15436 41608
rect 15752 41599 15804 41608
rect 15752 41565 15761 41599
rect 15761 41565 15795 41599
rect 15795 41565 15804 41599
rect 15752 41556 15804 41565
rect 20168 41556 20220 41608
rect 58164 41599 58216 41608
rect 58164 41565 58173 41599
rect 58173 41565 58207 41599
rect 58207 41565 58216 41599
rect 58164 41556 58216 41565
rect 13820 41420 13872 41472
rect 15200 41488 15252 41540
rect 16764 41488 16816 41540
rect 18420 41488 18472 41540
rect 19432 41531 19484 41540
rect 19432 41497 19441 41531
rect 19441 41497 19475 41531
rect 19475 41497 19484 41531
rect 19432 41488 19484 41497
rect 17684 41420 17736 41472
rect 19340 41420 19392 41472
rect 20260 41420 20312 41472
rect 20720 41420 20772 41472
rect 23480 41420 23532 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 10416 41216 10468 41268
rect 11796 41216 11848 41268
rect 12532 41148 12584 41200
rect 9864 41123 9916 41132
rect 9864 41089 9873 41123
rect 9873 41089 9907 41123
rect 9907 41089 9916 41123
rect 9864 41080 9916 41089
rect 9680 40944 9732 40996
rect 10968 41080 11020 41132
rect 13452 41123 13504 41132
rect 13452 41089 13461 41123
rect 13461 41089 13495 41123
rect 13495 41089 13504 41123
rect 15384 41123 15436 41132
rect 13452 41080 13504 41089
rect 15384 41089 15393 41123
rect 15393 41089 15427 41123
rect 15427 41089 15436 41123
rect 15384 41080 15436 41089
rect 15568 41216 15620 41268
rect 13636 41012 13688 41064
rect 13912 40987 13964 40996
rect 8300 40876 8352 40928
rect 9864 40876 9916 40928
rect 11428 40876 11480 40928
rect 13912 40953 13921 40987
rect 13921 40953 13955 40987
rect 13955 40953 13964 40987
rect 13912 40944 13964 40953
rect 19524 41080 19576 41132
rect 25320 41216 25372 41268
rect 23388 41148 23440 41200
rect 24400 41148 24452 41200
rect 20720 41123 20772 41132
rect 20720 41089 20729 41123
rect 20729 41089 20763 41123
rect 20763 41089 20772 41123
rect 20720 41080 20772 41089
rect 22192 41080 22244 41132
rect 23020 41123 23072 41132
rect 23020 41089 23029 41123
rect 23029 41089 23063 41123
rect 23063 41089 23072 41123
rect 23020 41080 23072 41089
rect 23112 41123 23164 41132
rect 23112 41089 23121 41123
rect 23121 41089 23155 41123
rect 23155 41089 23164 41123
rect 23112 41080 23164 41089
rect 23664 41080 23716 41132
rect 22928 41012 22980 41064
rect 15752 40944 15804 40996
rect 17776 40944 17828 40996
rect 20444 40944 20496 40996
rect 20628 40944 20680 40996
rect 15016 40876 15068 40928
rect 17500 40876 17552 40928
rect 18604 40876 18656 40928
rect 23296 40944 23348 40996
rect 22284 40876 22336 40928
rect 23480 40919 23532 40928
rect 23480 40885 23489 40919
rect 23489 40885 23523 40919
rect 23523 40885 23532 40919
rect 23480 40876 23532 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 12164 40672 12216 40724
rect 20628 40672 20680 40724
rect 23020 40672 23072 40724
rect 22100 40604 22152 40656
rect 23112 40604 23164 40656
rect 5264 40468 5316 40520
rect 9864 40468 9916 40520
rect 11428 40468 11480 40520
rect 5632 40400 5684 40452
rect 6460 40400 6512 40452
rect 6552 40375 6604 40384
rect 6552 40341 6561 40375
rect 6561 40341 6595 40375
rect 6595 40341 6604 40375
rect 6552 40332 6604 40341
rect 7564 40332 7616 40384
rect 12624 40468 12676 40520
rect 13728 40468 13780 40520
rect 16580 40468 16632 40520
rect 17500 40468 17552 40520
rect 20260 40536 20312 40588
rect 19340 40468 19392 40520
rect 13820 40400 13872 40452
rect 14280 40443 14332 40452
rect 14280 40409 14289 40443
rect 14289 40409 14323 40443
rect 14323 40409 14332 40443
rect 14280 40400 14332 40409
rect 16764 40400 16816 40452
rect 18420 40400 18472 40452
rect 20076 40468 20128 40520
rect 20628 40468 20680 40520
rect 22928 40511 22980 40520
rect 22928 40477 22937 40511
rect 22937 40477 22971 40511
rect 22971 40477 22980 40511
rect 22928 40468 22980 40477
rect 20444 40400 20496 40452
rect 21824 40400 21876 40452
rect 23020 40400 23072 40452
rect 23296 40511 23348 40520
rect 23296 40477 23325 40511
rect 23325 40477 23348 40511
rect 23296 40468 23348 40477
rect 32220 40468 32272 40520
rect 58164 40511 58216 40520
rect 58164 40477 58173 40511
rect 58173 40477 58207 40511
rect 58207 40477 58216 40511
rect 58164 40468 58216 40477
rect 24400 40443 24452 40452
rect 24400 40409 24409 40443
rect 24409 40409 24443 40443
rect 24443 40409 24452 40443
rect 24400 40400 24452 40409
rect 24860 40400 24912 40452
rect 30840 40400 30892 40452
rect 12348 40332 12400 40384
rect 12808 40332 12860 40384
rect 14924 40332 14976 40384
rect 15200 40332 15252 40384
rect 16028 40375 16080 40384
rect 16028 40341 16037 40375
rect 16037 40341 16071 40375
rect 16071 40341 16080 40375
rect 16028 40332 16080 40341
rect 20352 40332 20404 40384
rect 22192 40375 22244 40384
rect 22192 40341 22201 40375
rect 22201 40341 22235 40375
rect 22235 40341 22244 40375
rect 22192 40332 22244 40341
rect 22652 40332 22704 40384
rect 23572 40375 23624 40384
rect 23572 40341 23581 40375
rect 23581 40341 23615 40375
rect 23615 40341 23624 40375
rect 23572 40332 23624 40341
rect 32036 40332 32088 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4988 40128 5040 40180
rect 5540 40060 5592 40112
rect 3792 39992 3844 40044
rect 4804 39992 4856 40044
rect 6460 39992 6512 40044
rect 2504 39967 2556 39976
rect 2504 39933 2513 39967
rect 2513 39933 2547 39967
rect 2547 39933 2556 39967
rect 2504 39924 2556 39933
rect 6828 40035 6880 40044
rect 11336 40128 11388 40180
rect 13728 40128 13780 40180
rect 15016 40128 15068 40180
rect 21456 40128 21508 40180
rect 21824 40171 21876 40180
rect 21824 40137 21833 40171
rect 21833 40137 21867 40171
rect 21867 40137 21876 40171
rect 21824 40128 21876 40137
rect 22100 40128 22152 40180
rect 6828 40001 6842 40035
rect 6842 40001 6876 40035
rect 6876 40001 6880 40035
rect 6828 39992 6880 40001
rect 7748 40035 7800 40044
rect 7748 40001 7782 40035
rect 7782 40001 7800 40035
rect 5816 39899 5868 39908
rect 5816 39865 5825 39899
rect 5825 39865 5859 39899
rect 5859 39865 5868 39899
rect 5816 39856 5868 39865
rect 6644 39856 6696 39908
rect 6736 39856 6788 39908
rect 4620 39788 4672 39840
rect 5264 39831 5316 39840
rect 5264 39797 5273 39831
rect 5273 39797 5307 39831
rect 5307 39797 5316 39831
rect 5264 39788 5316 39797
rect 6368 39831 6420 39840
rect 6368 39797 6377 39831
rect 6377 39797 6411 39831
rect 6411 39797 6420 39831
rect 6368 39788 6420 39797
rect 7748 39992 7800 40001
rect 9864 40060 9916 40112
rect 18420 40060 18472 40112
rect 19248 40060 19300 40112
rect 8852 39831 8904 39840
rect 8852 39797 8861 39831
rect 8861 39797 8895 39831
rect 8895 39797 8904 39831
rect 8852 39788 8904 39797
rect 10968 39992 11020 40044
rect 11520 39856 11572 39908
rect 11796 40035 11848 40044
rect 11796 40001 11805 40035
rect 11805 40001 11839 40035
rect 11839 40001 11848 40035
rect 11796 39992 11848 40001
rect 12624 39992 12676 40044
rect 14556 39992 14608 40044
rect 15660 39924 15712 39976
rect 16488 39924 16540 39976
rect 11796 39856 11848 39908
rect 12624 39831 12676 39840
rect 12624 39797 12633 39831
rect 12633 39797 12667 39831
rect 12667 39797 12676 39831
rect 12624 39788 12676 39797
rect 21456 39992 21508 40044
rect 23020 40128 23072 40180
rect 23388 40128 23440 40180
rect 23756 40128 23808 40180
rect 29184 40128 29236 40180
rect 23572 40060 23624 40112
rect 22284 40035 22336 40044
rect 22284 40001 22293 40035
rect 22293 40001 22327 40035
rect 22327 40001 22336 40035
rect 22284 39992 22336 40001
rect 18328 39967 18380 39976
rect 18328 39933 18337 39967
rect 18337 39933 18371 39967
rect 18371 39933 18380 39967
rect 18328 39924 18380 39933
rect 19432 39924 19484 39976
rect 22928 39992 22980 40044
rect 20076 39856 20128 39908
rect 22192 39856 22244 39908
rect 23388 39992 23440 40044
rect 23664 39992 23716 40044
rect 28356 39992 28408 40044
rect 23848 39967 23900 39976
rect 23848 39933 23857 39967
rect 23857 39933 23891 39967
rect 23891 39933 23900 39967
rect 23848 39924 23900 39933
rect 23204 39856 23256 39908
rect 23756 39856 23808 39908
rect 25228 39788 25280 39840
rect 27620 39788 27672 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 3792 39627 3844 39636
rect 3792 39593 3801 39627
rect 3801 39593 3835 39627
rect 3835 39593 3844 39627
rect 3792 39584 3844 39593
rect 4620 39584 4672 39636
rect 5632 39627 5684 39636
rect 5632 39593 5641 39627
rect 5641 39593 5675 39627
rect 5675 39593 5684 39627
rect 5632 39584 5684 39593
rect 5356 39516 5408 39568
rect 6736 39584 6788 39636
rect 11520 39627 11572 39636
rect 11520 39593 11529 39627
rect 11529 39593 11563 39627
rect 11563 39593 11572 39627
rect 11520 39584 11572 39593
rect 14556 39584 14608 39636
rect 19340 39584 19392 39636
rect 30840 39627 30892 39636
rect 30840 39593 30849 39627
rect 30849 39593 30883 39627
rect 30883 39593 30892 39627
rect 30840 39584 30892 39593
rect 4988 39423 5040 39432
rect 4988 39389 4997 39423
rect 4997 39389 5031 39423
rect 5031 39389 5040 39423
rect 4988 39380 5040 39389
rect 5448 39448 5500 39500
rect 13452 39448 13504 39500
rect 5816 39380 5868 39432
rect 6368 39423 6420 39432
rect 6368 39389 6402 39423
rect 6402 39389 6420 39423
rect 6368 39380 6420 39389
rect 9864 39380 9916 39432
rect 6276 39312 6328 39364
rect 10048 39312 10100 39364
rect 11152 39355 11204 39364
rect 11152 39321 11161 39355
rect 11161 39321 11195 39355
rect 11195 39321 11204 39355
rect 11152 39312 11204 39321
rect 11336 39355 11388 39364
rect 11336 39321 11345 39355
rect 11345 39321 11379 39355
rect 11379 39321 11388 39355
rect 11336 39312 11388 39321
rect 11980 39312 12032 39364
rect 14556 39380 14608 39432
rect 13636 39312 13688 39364
rect 14924 39420 14976 39432
rect 14924 39386 14933 39420
rect 14933 39386 14967 39420
rect 14967 39386 14976 39420
rect 14924 39380 14976 39386
rect 16488 39380 16540 39432
rect 18328 39380 18380 39432
rect 19432 39380 19484 39432
rect 20628 39423 20680 39432
rect 20628 39389 20637 39423
rect 20637 39389 20671 39423
rect 20671 39389 20680 39423
rect 20628 39380 20680 39389
rect 23848 39380 23900 39432
rect 24400 39423 24452 39432
rect 24400 39389 24409 39423
rect 24409 39389 24443 39423
rect 24443 39389 24452 39423
rect 24400 39380 24452 39389
rect 5264 39244 5316 39296
rect 7104 39244 7156 39296
rect 8116 39244 8168 39296
rect 11244 39244 11296 39296
rect 12716 39244 12768 39296
rect 14556 39244 14608 39296
rect 16672 39287 16724 39296
rect 16672 39253 16681 39287
rect 16681 39253 16715 39287
rect 16715 39253 16724 39287
rect 16672 39244 16724 39253
rect 17776 39355 17828 39364
rect 17776 39321 17794 39355
rect 17794 39321 17828 39355
rect 17776 39312 17828 39321
rect 20260 39312 20312 39364
rect 20352 39355 20404 39364
rect 20352 39321 20370 39355
rect 20370 39321 20404 39355
rect 20352 39312 20404 39321
rect 23480 39312 23532 39364
rect 27252 39312 27304 39364
rect 27620 39312 27672 39364
rect 31576 39380 31628 39432
rect 20076 39244 20128 39296
rect 24860 39244 24912 39296
rect 28816 39244 28868 39296
rect 29000 39244 29052 39296
rect 30380 39287 30432 39296
rect 30380 39253 30389 39287
rect 30389 39253 30423 39287
rect 30423 39253 30432 39287
rect 30380 39244 30432 39253
rect 31116 39244 31168 39296
rect 31484 39244 31536 39296
rect 32036 39312 32088 39364
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 6828 39040 6880 39092
rect 8392 39040 8444 39092
rect 4160 38904 4212 38956
rect 5448 38972 5500 39024
rect 7104 39015 7156 39024
rect 7104 38981 7113 39015
rect 7113 38981 7147 39015
rect 7147 38981 7156 39015
rect 7104 38972 7156 38981
rect 4620 38836 4672 38888
rect 5080 38836 5132 38888
rect 6828 38836 6880 38888
rect 1952 38700 2004 38752
rect 3976 38700 4028 38752
rect 9864 38700 9916 38752
rect 13636 38904 13688 38956
rect 29000 38904 29052 38956
rect 30196 38904 30248 38956
rect 12716 38768 12768 38820
rect 11796 38700 11848 38752
rect 23388 38700 23440 38752
rect 26976 38700 27028 38752
rect 27620 38700 27672 38752
rect 58164 38811 58216 38820
rect 58164 38777 58173 38811
rect 58173 38777 58207 38811
rect 58207 38777 58216 38811
rect 58164 38768 58216 38777
rect 29736 38700 29788 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 4804 38496 4856 38548
rect 6276 38496 6328 38548
rect 10048 38539 10100 38548
rect 10048 38505 10057 38539
rect 10057 38505 10091 38539
rect 10091 38505 10100 38539
rect 10048 38496 10100 38505
rect 14280 38496 14332 38548
rect 23388 38496 23440 38548
rect 27252 38539 27304 38548
rect 27252 38505 27261 38539
rect 27261 38505 27295 38539
rect 27295 38505 27304 38539
rect 27252 38496 27304 38505
rect 28356 38539 28408 38548
rect 28356 38505 28365 38539
rect 28365 38505 28399 38539
rect 28399 38505 28408 38539
rect 28356 38496 28408 38505
rect 9680 38428 9732 38480
rect 10416 38428 10468 38480
rect 12624 38428 12676 38480
rect 18144 38428 18196 38480
rect 3976 38360 4028 38412
rect 4436 38360 4488 38412
rect 5356 38360 5408 38412
rect 2872 38335 2924 38344
rect 2872 38301 2881 38335
rect 2881 38301 2915 38335
rect 2915 38301 2924 38335
rect 2872 38292 2924 38301
rect 1952 38267 2004 38276
rect 1952 38233 1961 38267
rect 1961 38233 1995 38267
rect 1995 38233 2004 38267
rect 1952 38224 2004 38233
rect 1768 38199 1820 38208
rect 1768 38165 1777 38199
rect 1777 38165 1811 38199
rect 1811 38165 1820 38199
rect 1768 38156 1820 38165
rect 2688 38156 2740 38208
rect 5080 38292 5132 38344
rect 6552 38335 6604 38344
rect 6552 38301 6561 38335
rect 6561 38301 6595 38335
rect 6595 38301 6604 38335
rect 6552 38292 6604 38301
rect 8392 38335 8444 38344
rect 8392 38301 8401 38335
rect 8401 38301 8435 38335
rect 8435 38301 8444 38335
rect 8392 38292 8444 38301
rect 8852 38292 8904 38344
rect 9404 38335 9456 38344
rect 9404 38301 9413 38335
rect 9413 38301 9447 38335
rect 9447 38301 9456 38335
rect 9404 38292 9456 38301
rect 10232 38292 10284 38344
rect 20628 38403 20680 38412
rect 10968 38292 11020 38344
rect 11244 38292 11296 38344
rect 12624 38292 12676 38344
rect 20628 38369 20637 38403
rect 20637 38369 20671 38403
rect 20671 38369 20680 38403
rect 20628 38360 20680 38369
rect 13360 38335 13412 38344
rect 13360 38301 13369 38335
rect 13369 38301 13403 38335
rect 13403 38301 13412 38335
rect 13360 38292 13412 38301
rect 5356 38224 5408 38276
rect 5908 38267 5960 38276
rect 5908 38233 5917 38267
rect 5917 38233 5951 38267
rect 5951 38233 5960 38267
rect 5908 38224 5960 38233
rect 6736 38267 6788 38276
rect 6736 38233 6745 38267
rect 6745 38233 6779 38267
rect 6779 38233 6788 38267
rect 6736 38224 6788 38233
rect 4436 38156 4488 38208
rect 4620 38199 4672 38208
rect 4620 38165 4629 38199
rect 4629 38165 4663 38199
rect 4663 38165 4672 38199
rect 4620 38156 4672 38165
rect 11152 38224 11204 38276
rect 11520 38267 11572 38276
rect 11520 38233 11529 38267
rect 11529 38233 11563 38267
rect 11563 38233 11572 38267
rect 11520 38224 11572 38233
rect 13176 38267 13228 38276
rect 13176 38233 13185 38267
rect 13185 38233 13219 38267
rect 13219 38233 13228 38267
rect 13176 38224 13228 38233
rect 16672 38224 16724 38276
rect 19432 38224 19484 38276
rect 9496 38156 9548 38208
rect 27712 38335 27764 38344
rect 27712 38301 27721 38335
rect 27721 38301 27755 38335
rect 27755 38301 27764 38335
rect 27712 38292 27764 38301
rect 27988 38292 28040 38344
rect 31116 38360 31168 38412
rect 32220 38403 32272 38412
rect 32220 38369 32229 38403
rect 32229 38369 32263 38403
rect 32263 38369 32272 38403
rect 32680 38403 32732 38412
rect 32220 38360 32272 38369
rect 32680 38369 32689 38403
rect 32689 38369 32723 38403
rect 32723 38369 32732 38403
rect 32680 38360 32732 38369
rect 28908 38292 28960 38344
rect 29276 38292 29328 38344
rect 30748 38292 30800 38344
rect 31484 38292 31536 38344
rect 30104 38224 30156 38276
rect 17132 38156 17184 38208
rect 19064 38156 19116 38208
rect 27068 38156 27120 38208
rect 30472 38156 30524 38208
rect 31024 38224 31076 38276
rect 33048 38224 33100 38276
rect 31392 38156 31444 38208
rect 33876 38156 33928 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4160 37952 4212 38004
rect 5356 37995 5408 38004
rect 5356 37961 5365 37995
rect 5365 37961 5399 37995
rect 5399 37961 5408 37995
rect 5356 37952 5408 37961
rect 1768 37884 1820 37936
rect 2504 37816 2556 37868
rect 2688 37859 2740 37868
rect 2688 37825 2722 37859
rect 2722 37825 2740 37859
rect 2688 37816 2740 37825
rect 4804 37884 4856 37936
rect 6736 37952 6788 38004
rect 10232 37952 10284 38004
rect 10784 37995 10836 38004
rect 10784 37961 10793 37995
rect 10793 37961 10827 37995
rect 10827 37961 10836 37995
rect 10784 37952 10836 37961
rect 4436 37748 4488 37800
rect 5080 37816 5132 37868
rect 4804 37748 4856 37800
rect 9404 37816 9456 37868
rect 11612 37816 11664 37868
rect 13176 37952 13228 38004
rect 12164 37884 12216 37936
rect 18328 37952 18380 38004
rect 19340 37952 19392 38004
rect 27712 37952 27764 38004
rect 28908 37995 28960 38004
rect 28908 37961 28917 37995
rect 28917 37961 28951 37995
rect 28951 37961 28960 37995
rect 28908 37952 28960 37961
rect 29828 37952 29880 38004
rect 31024 37995 31076 38004
rect 11888 37859 11940 37868
rect 11888 37825 11897 37859
rect 11897 37825 11931 37859
rect 11931 37825 11940 37859
rect 11888 37816 11940 37825
rect 11980 37816 12032 37868
rect 13268 37816 13320 37868
rect 16028 37816 16080 37868
rect 17132 37859 17184 37868
rect 17132 37825 17141 37859
rect 17141 37825 17175 37859
rect 17175 37825 17184 37859
rect 17132 37816 17184 37825
rect 12624 37748 12676 37800
rect 17040 37748 17092 37800
rect 17500 37859 17552 37868
rect 17500 37825 17509 37859
rect 17509 37825 17543 37859
rect 17543 37825 17552 37859
rect 17500 37816 17552 37825
rect 18512 37816 18564 37868
rect 19064 37859 19116 37868
rect 19064 37825 19071 37859
rect 19071 37825 19116 37859
rect 19064 37816 19116 37825
rect 20076 37884 20128 37936
rect 18328 37748 18380 37800
rect 20168 37859 20220 37868
rect 20168 37825 20177 37859
rect 20177 37825 20211 37859
rect 20211 37825 20220 37859
rect 20168 37816 20220 37825
rect 20444 37884 20496 37936
rect 26516 37884 26568 37936
rect 28816 37884 28868 37936
rect 29276 37927 29328 37936
rect 24308 37816 24360 37868
rect 26240 37816 26292 37868
rect 29276 37893 29285 37927
rect 29285 37893 29319 37927
rect 29319 37893 29328 37927
rect 29276 37884 29328 37893
rect 30472 37884 30524 37936
rect 29184 37816 29236 37868
rect 30104 37816 30156 37868
rect 31024 37961 31033 37995
rect 31033 37961 31067 37995
rect 31067 37961 31076 37995
rect 31024 37952 31076 37961
rect 33048 37995 33100 38004
rect 33048 37961 33057 37995
rect 33057 37961 33091 37995
rect 33091 37961 33100 37995
rect 33048 37952 33100 37961
rect 34612 37952 34664 38004
rect 31300 37816 31352 37868
rect 31576 37816 31628 37868
rect 32588 37859 32640 37868
rect 32588 37825 32597 37859
rect 32597 37825 32631 37859
rect 32631 37825 32640 37859
rect 32588 37816 32640 37825
rect 5724 37680 5776 37732
rect 5908 37680 5960 37732
rect 11796 37680 11848 37732
rect 4712 37612 4764 37664
rect 10784 37612 10836 37664
rect 13636 37612 13688 37664
rect 13912 37680 13964 37732
rect 31024 37748 31076 37800
rect 34244 37816 34296 37868
rect 34520 37859 34572 37868
rect 34520 37825 34529 37859
rect 34529 37825 34563 37859
rect 34563 37825 34572 37859
rect 34520 37816 34572 37825
rect 21272 37680 21324 37732
rect 26516 37680 26568 37732
rect 27436 37680 27488 37732
rect 16948 37612 17000 37664
rect 17500 37612 17552 37664
rect 20996 37612 21048 37664
rect 22284 37612 22336 37664
rect 23112 37655 23164 37664
rect 23112 37621 23121 37655
rect 23121 37621 23155 37655
rect 23155 37621 23164 37655
rect 23112 37612 23164 37621
rect 25596 37655 25648 37664
rect 25596 37621 25605 37655
rect 25605 37621 25639 37655
rect 25639 37621 25648 37655
rect 25596 37612 25648 37621
rect 34152 37612 34204 37664
rect 35348 37612 35400 37664
rect 58164 37655 58216 37664
rect 58164 37621 58173 37655
rect 58173 37621 58207 37655
rect 58207 37621 58216 37655
rect 58164 37612 58216 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 20168 37451 20220 37460
rect 20168 37417 20177 37451
rect 20177 37417 20211 37451
rect 20211 37417 20220 37451
rect 20168 37408 20220 37417
rect 26240 37451 26292 37460
rect 26240 37417 26249 37451
rect 26249 37417 26283 37451
rect 26283 37417 26292 37451
rect 26240 37408 26292 37417
rect 30104 37408 30156 37460
rect 31300 37408 31352 37460
rect 32680 37408 32732 37460
rect 5724 37272 5776 37324
rect 13360 37315 13412 37324
rect 13360 37281 13369 37315
rect 13369 37281 13403 37315
rect 13403 37281 13412 37315
rect 13360 37272 13412 37281
rect 4620 37204 4672 37256
rect 7840 37247 7892 37256
rect 7012 37136 7064 37188
rect 7840 37213 7849 37247
rect 7849 37213 7883 37247
rect 7883 37213 7892 37247
rect 7840 37204 7892 37213
rect 8116 37247 8168 37256
rect 8116 37213 8125 37247
rect 8125 37213 8159 37247
rect 8159 37213 8168 37247
rect 8116 37204 8168 37213
rect 8208 37247 8260 37256
rect 8208 37213 8217 37247
rect 8217 37213 8251 37247
rect 8251 37213 8260 37247
rect 8208 37204 8260 37213
rect 11888 37204 11940 37256
rect 13268 37204 13320 37256
rect 15660 37247 15712 37256
rect 15660 37213 15669 37247
rect 15669 37213 15703 37247
rect 15703 37213 15712 37247
rect 15660 37204 15712 37213
rect 7932 37136 7984 37188
rect 11612 37136 11664 37188
rect 8300 37068 8352 37120
rect 11796 37068 11848 37120
rect 12716 37068 12768 37120
rect 13636 37136 13688 37188
rect 16672 37136 16724 37188
rect 18512 37247 18564 37256
rect 18512 37213 18526 37247
rect 18526 37213 18560 37247
rect 18560 37213 18564 37247
rect 18512 37204 18564 37213
rect 18328 37179 18380 37188
rect 15476 37068 15528 37120
rect 18328 37145 18337 37179
rect 18337 37145 18371 37179
rect 18371 37145 18380 37179
rect 18328 37136 18380 37145
rect 17040 37111 17092 37120
rect 17040 37077 17049 37111
rect 17049 37077 17083 37111
rect 17083 37077 17092 37111
rect 17040 37068 17092 37077
rect 18696 37111 18748 37120
rect 18696 37077 18705 37111
rect 18705 37077 18739 37111
rect 18739 37077 18748 37111
rect 18696 37068 18748 37077
rect 19340 37068 19392 37120
rect 20996 37204 21048 37256
rect 21916 37204 21968 37256
rect 22284 37204 22336 37256
rect 23204 37204 23256 37256
rect 24400 37247 24452 37256
rect 24400 37213 24409 37247
rect 24409 37213 24443 37247
rect 24443 37213 24452 37247
rect 24400 37204 24452 37213
rect 26516 37247 26568 37256
rect 26516 37213 26525 37247
rect 26525 37213 26559 37247
rect 26559 37213 26568 37247
rect 26516 37204 26568 37213
rect 22744 37111 22796 37120
rect 22744 37077 22753 37111
rect 22753 37077 22787 37111
rect 22787 37077 22796 37111
rect 22744 37068 22796 37077
rect 23112 37179 23164 37188
rect 23112 37145 23121 37179
rect 23121 37145 23155 37179
rect 23155 37145 23164 37179
rect 23112 37136 23164 37145
rect 24676 37179 24728 37188
rect 24676 37145 24710 37179
rect 24710 37145 24728 37179
rect 24676 37136 24728 37145
rect 24952 37136 25004 37188
rect 26700 37247 26752 37256
rect 26700 37213 26709 37247
rect 26709 37213 26743 37247
rect 26743 37213 26752 37247
rect 26700 37204 26752 37213
rect 26884 37247 26936 37256
rect 26884 37213 26893 37247
rect 26893 37213 26927 37247
rect 26927 37213 26936 37247
rect 26884 37204 26936 37213
rect 34796 37204 34848 37256
rect 35348 37247 35400 37256
rect 35348 37213 35382 37247
rect 35382 37213 35400 37247
rect 35348 37204 35400 37213
rect 30288 37136 30340 37188
rect 26240 37068 26292 37120
rect 27988 37068 28040 37120
rect 30104 37068 30156 37120
rect 35532 37068 35584 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 15476 36907 15528 36916
rect 6552 36796 6604 36848
rect 7840 36839 7892 36848
rect 7840 36805 7849 36839
rect 7849 36805 7883 36839
rect 7883 36805 7892 36839
rect 7840 36796 7892 36805
rect 5172 36728 5224 36780
rect 8208 36796 8260 36848
rect 8024 36771 8076 36780
rect 8024 36737 8033 36771
rect 8033 36737 8067 36771
rect 8067 36737 8076 36771
rect 8024 36728 8076 36737
rect 9956 36728 10008 36780
rect 12348 36728 12400 36780
rect 14740 36728 14792 36780
rect 7932 36660 7984 36712
rect 13268 36703 13320 36712
rect 13268 36669 13277 36703
rect 13277 36669 13311 36703
rect 13311 36669 13320 36703
rect 13268 36660 13320 36669
rect 12992 36592 13044 36644
rect 15476 36873 15485 36907
rect 15485 36873 15519 36907
rect 15519 36873 15528 36907
rect 15476 36864 15528 36873
rect 16672 36907 16724 36916
rect 16672 36873 16681 36907
rect 16681 36873 16715 36907
rect 16715 36873 16724 36907
rect 16672 36864 16724 36873
rect 19432 36864 19484 36916
rect 30196 36864 30248 36916
rect 32588 36864 32640 36916
rect 34520 36864 34572 36916
rect 16948 36771 17000 36780
rect 16948 36737 16957 36771
rect 16957 36737 16991 36771
rect 16991 36737 17000 36771
rect 16948 36728 17000 36737
rect 16856 36660 16908 36712
rect 17132 36771 17184 36780
rect 17132 36737 17141 36771
rect 17141 36737 17175 36771
rect 17175 36737 17184 36771
rect 18236 36796 18288 36848
rect 19064 36839 19116 36848
rect 17132 36728 17184 36737
rect 18144 36771 18196 36780
rect 18144 36737 18153 36771
rect 18153 36737 18187 36771
rect 18187 36737 18196 36771
rect 19064 36805 19073 36839
rect 19073 36805 19107 36839
rect 19107 36805 19116 36839
rect 19064 36796 19116 36805
rect 21916 36796 21968 36848
rect 24400 36796 24452 36848
rect 29000 36796 29052 36848
rect 30288 36796 30340 36848
rect 33876 36796 33928 36848
rect 34060 36796 34112 36848
rect 18144 36728 18196 36737
rect 22284 36771 22336 36780
rect 22284 36737 22293 36771
rect 22293 36737 22327 36771
rect 22327 36737 22336 36771
rect 22284 36728 22336 36737
rect 22468 36771 22520 36780
rect 22468 36737 22477 36771
rect 22477 36737 22511 36771
rect 22511 36737 22520 36771
rect 22652 36771 22704 36780
rect 22468 36728 22520 36737
rect 22652 36737 22661 36771
rect 22661 36737 22695 36771
rect 22695 36737 22704 36771
rect 22652 36728 22704 36737
rect 25688 36728 25740 36780
rect 26240 36771 26292 36780
rect 26240 36737 26249 36771
rect 26249 36737 26283 36771
rect 26283 36737 26292 36771
rect 26240 36728 26292 36737
rect 27620 36771 27672 36780
rect 27620 36737 27629 36771
rect 27629 36737 27663 36771
rect 27663 36737 27672 36771
rect 27620 36728 27672 36737
rect 27712 36728 27764 36780
rect 28908 36728 28960 36780
rect 29552 36728 29604 36780
rect 25596 36660 25648 36712
rect 30104 36728 30156 36780
rect 31300 36771 31352 36780
rect 31300 36737 31309 36771
rect 31309 36737 31343 36771
rect 31343 36737 31352 36771
rect 31300 36728 31352 36737
rect 33232 36771 33284 36780
rect 33232 36737 33241 36771
rect 33241 36737 33275 36771
rect 33275 36737 33284 36771
rect 33232 36728 33284 36737
rect 34244 36771 34296 36780
rect 34244 36737 34253 36771
rect 34253 36737 34287 36771
rect 34287 36737 34296 36771
rect 34244 36728 34296 36737
rect 35348 36771 35400 36780
rect 30564 36660 30616 36712
rect 31576 36703 31628 36712
rect 31576 36669 31585 36703
rect 31585 36669 31619 36703
rect 31619 36669 31628 36703
rect 31576 36660 31628 36669
rect 33600 36660 33652 36712
rect 18144 36592 18196 36644
rect 34428 36592 34480 36644
rect 35348 36737 35357 36771
rect 35357 36737 35391 36771
rect 35391 36737 35400 36771
rect 35348 36728 35400 36737
rect 35532 36771 35584 36780
rect 35532 36737 35541 36771
rect 35541 36737 35575 36771
rect 35575 36737 35584 36771
rect 35532 36728 35584 36737
rect 7196 36567 7248 36576
rect 7196 36533 7205 36567
rect 7205 36533 7239 36567
rect 7239 36533 7248 36567
rect 7196 36524 7248 36533
rect 7472 36524 7524 36576
rect 19432 36524 19484 36576
rect 20076 36524 20128 36576
rect 21364 36524 21416 36576
rect 22468 36524 22520 36576
rect 22652 36524 22704 36576
rect 23112 36567 23164 36576
rect 23112 36533 23121 36567
rect 23121 36533 23155 36567
rect 23155 36533 23164 36567
rect 23112 36524 23164 36533
rect 25044 36524 25096 36576
rect 29276 36524 29328 36576
rect 33692 36567 33744 36576
rect 33692 36533 33701 36567
rect 33701 36533 33735 36567
rect 33735 36533 33744 36567
rect 33692 36524 33744 36533
rect 34704 36524 34756 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 5172 36363 5224 36372
rect 5172 36329 5181 36363
rect 5181 36329 5215 36363
rect 5215 36329 5224 36363
rect 5172 36320 5224 36329
rect 7012 36363 7064 36372
rect 7012 36329 7021 36363
rect 7021 36329 7055 36363
rect 7055 36329 7064 36363
rect 7012 36320 7064 36329
rect 9496 36363 9548 36372
rect 9496 36329 9505 36363
rect 9505 36329 9539 36363
rect 9539 36329 9548 36363
rect 9496 36320 9548 36329
rect 11428 36320 11480 36372
rect 12348 36320 12400 36372
rect 14740 36363 14792 36372
rect 14740 36329 14749 36363
rect 14749 36329 14783 36363
rect 14783 36329 14792 36363
rect 14740 36320 14792 36329
rect 17132 36320 17184 36372
rect 18052 36320 18104 36372
rect 24676 36320 24728 36372
rect 26700 36320 26752 36372
rect 27712 36363 27764 36372
rect 27712 36329 27721 36363
rect 27721 36329 27755 36363
rect 27755 36329 27764 36363
rect 27712 36320 27764 36329
rect 29552 36363 29604 36372
rect 29552 36329 29561 36363
rect 29561 36329 29595 36363
rect 29595 36329 29604 36363
rect 29552 36320 29604 36329
rect 34060 36320 34112 36372
rect 24768 36252 24820 36304
rect 25688 36252 25740 36304
rect 16856 36184 16908 36236
rect 24308 36184 24360 36236
rect 2504 36116 2556 36168
rect 4620 36116 4672 36168
rect 7380 36159 7432 36168
rect 7380 36125 7389 36159
rect 7389 36125 7423 36159
rect 7423 36125 7432 36159
rect 7380 36116 7432 36125
rect 7472 36159 7524 36168
rect 7472 36125 7486 36159
rect 7486 36125 7520 36159
rect 7520 36125 7524 36159
rect 7472 36116 7524 36125
rect 8944 36116 8996 36168
rect 9864 36116 9916 36168
rect 14096 36159 14148 36168
rect 14096 36125 14105 36159
rect 14105 36125 14139 36159
rect 14139 36125 14148 36159
rect 14096 36116 14148 36125
rect 4620 35980 4672 36032
rect 6552 36023 6604 36032
rect 6552 35989 6561 36023
rect 6561 35989 6595 36023
rect 6595 35989 6604 36023
rect 6552 35980 6604 35989
rect 10324 36048 10376 36100
rect 11796 36091 11848 36100
rect 11796 36057 11805 36091
rect 11805 36057 11839 36091
rect 11839 36057 11848 36091
rect 11796 36048 11848 36057
rect 14372 36159 14424 36168
rect 14372 36125 14381 36159
rect 14381 36125 14415 36159
rect 14415 36125 14424 36159
rect 14372 36116 14424 36125
rect 15016 36116 15068 36168
rect 15476 36116 15528 36168
rect 17040 36116 17092 36168
rect 24676 36116 24728 36168
rect 24952 36159 25004 36168
rect 24952 36125 24961 36159
rect 24961 36125 24995 36159
rect 24995 36125 25004 36159
rect 24952 36116 25004 36125
rect 25044 36159 25096 36168
rect 25044 36125 25053 36159
rect 25053 36125 25087 36159
rect 25087 36125 25096 36159
rect 26884 36184 26936 36236
rect 25044 36116 25096 36125
rect 25596 36116 25648 36168
rect 27988 36159 28040 36168
rect 15660 36048 15712 36100
rect 18236 36048 18288 36100
rect 25688 36091 25740 36100
rect 25688 36057 25697 36091
rect 25697 36057 25731 36091
rect 25731 36057 25740 36091
rect 25688 36048 25740 36057
rect 27988 36125 27997 36159
rect 27997 36125 28031 36159
rect 28031 36125 28040 36159
rect 27988 36116 28040 36125
rect 30564 36184 30616 36236
rect 34796 36227 34848 36236
rect 34796 36193 34805 36227
rect 34805 36193 34839 36227
rect 34839 36193 34848 36227
rect 34796 36184 34848 36193
rect 28172 36159 28224 36168
rect 28172 36125 28181 36159
rect 28181 36125 28215 36159
rect 28215 36125 28224 36159
rect 28172 36116 28224 36125
rect 29736 36159 29788 36168
rect 27896 36048 27948 36100
rect 29736 36125 29745 36159
rect 29745 36125 29779 36159
rect 29779 36125 29788 36159
rect 29736 36116 29788 36125
rect 28908 36091 28960 36100
rect 28908 36057 28917 36091
rect 28917 36057 28951 36091
rect 28951 36057 28960 36091
rect 28908 36048 28960 36057
rect 29920 36091 29972 36100
rect 29920 36057 29929 36091
rect 29929 36057 29963 36091
rect 29963 36057 29972 36091
rect 29920 36048 29972 36057
rect 10140 35980 10192 36032
rect 11336 36023 11388 36032
rect 11336 35989 11345 36023
rect 11345 35989 11379 36023
rect 11379 35989 11388 36023
rect 11336 35980 11388 35989
rect 16948 35980 17000 36032
rect 18604 35980 18656 36032
rect 22652 35980 22704 36032
rect 23020 36023 23072 36032
rect 23020 35989 23029 36023
rect 23029 35989 23063 36023
rect 23063 35989 23072 36023
rect 23020 35980 23072 35989
rect 27160 36023 27212 36032
rect 27160 35989 27169 36023
rect 27169 35989 27203 36023
rect 27203 35989 27212 36023
rect 27160 35980 27212 35989
rect 30656 36023 30708 36032
rect 30656 35989 30665 36023
rect 30665 35989 30699 36023
rect 30699 35989 30708 36023
rect 30656 35980 30708 35989
rect 31576 35980 31628 36032
rect 33600 36116 33652 36168
rect 33784 36159 33836 36168
rect 33784 36125 33793 36159
rect 33793 36125 33827 36159
rect 33827 36125 33836 36159
rect 33784 36116 33836 36125
rect 34704 36116 34756 36168
rect 58164 36159 58216 36168
rect 58164 36125 58173 36159
rect 58173 36125 58207 36159
rect 58207 36125 58216 36159
rect 58164 36116 58216 36125
rect 34704 35980 34756 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 9772 35776 9824 35828
rect 14096 35776 14148 35828
rect 5172 35708 5224 35760
rect 4896 35640 4948 35692
rect 7472 35683 7524 35692
rect 7472 35649 7490 35683
rect 7490 35649 7524 35683
rect 7472 35640 7524 35649
rect 11060 35708 11112 35760
rect 11520 35751 11572 35760
rect 11520 35717 11529 35751
rect 11529 35717 11563 35751
rect 11563 35717 11572 35751
rect 11520 35708 11572 35717
rect 11612 35708 11664 35760
rect 9864 35640 9916 35692
rect 9956 35683 10008 35692
rect 9956 35649 9965 35683
rect 9965 35649 9999 35683
rect 9999 35649 10008 35683
rect 9956 35640 10008 35649
rect 10140 35640 10192 35692
rect 10784 35640 10836 35692
rect 10968 35640 11020 35692
rect 11704 35683 11756 35692
rect 11704 35649 11713 35683
rect 11713 35649 11747 35683
rect 11747 35649 11756 35683
rect 11704 35640 11756 35649
rect 13360 35708 13412 35760
rect 13636 35708 13688 35760
rect 27896 35776 27948 35828
rect 28172 35776 28224 35828
rect 28632 35776 28684 35828
rect 30104 35776 30156 35828
rect 30564 35776 30616 35828
rect 15016 35708 15068 35760
rect 18236 35751 18288 35760
rect 18236 35717 18245 35751
rect 18245 35717 18279 35751
rect 18279 35717 18288 35751
rect 18236 35708 18288 35717
rect 22652 35708 22704 35760
rect 29276 35708 29328 35760
rect 18052 35683 18104 35692
rect 18052 35649 18061 35683
rect 18061 35649 18095 35683
rect 18095 35649 18104 35683
rect 18052 35640 18104 35649
rect 22376 35640 22428 35692
rect 23020 35683 23072 35692
rect 23020 35649 23029 35683
rect 23029 35649 23063 35683
rect 23063 35649 23072 35683
rect 23020 35640 23072 35649
rect 23112 35683 23164 35692
rect 23112 35649 23121 35683
rect 23121 35649 23155 35683
rect 23155 35649 23164 35683
rect 23112 35640 23164 35649
rect 24860 35640 24912 35692
rect 29920 35640 29972 35692
rect 30196 35640 30248 35692
rect 8024 35572 8076 35624
rect 8944 35572 8996 35624
rect 13544 35572 13596 35624
rect 17040 35504 17092 35556
rect 29828 35504 29880 35556
rect 30472 35504 30524 35556
rect 4804 35479 4856 35488
rect 4804 35445 4813 35479
rect 4813 35445 4847 35479
rect 4847 35445 4856 35479
rect 4804 35436 4856 35445
rect 6644 35436 6696 35488
rect 10968 35436 11020 35488
rect 17960 35436 18012 35488
rect 22376 35479 22428 35488
rect 22376 35445 22385 35479
rect 22385 35445 22419 35479
rect 22419 35445 22428 35479
rect 22376 35436 22428 35445
rect 23020 35436 23072 35488
rect 24308 35436 24360 35488
rect 24676 35436 24728 35488
rect 25320 35436 25372 35488
rect 25964 35436 26016 35488
rect 30932 35479 30984 35488
rect 30932 35445 30941 35479
rect 30941 35445 30975 35479
rect 30975 35445 30984 35479
rect 30932 35436 30984 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4620 35232 4672 35284
rect 7472 35232 7524 35284
rect 18052 35232 18104 35284
rect 25964 35232 26016 35284
rect 30104 35232 30156 35284
rect 30472 35232 30524 35284
rect 3240 35096 3292 35148
rect 7380 35164 7432 35216
rect 4804 35071 4856 35080
rect 4804 35037 4813 35071
rect 4813 35037 4847 35071
rect 4847 35037 4856 35071
rect 4804 35028 4856 35037
rect 4988 35071 5040 35080
rect 4988 35037 4997 35071
rect 4997 35037 5031 35071
rect 5031 35037 5040 35071
rect 7564 35071 7616 35080
rect 4988 35028 5040 35037
rect 7564 35037 7573 35071
rect 7573 35037 7607 35071
rect 7607 35037 7616 35071
rect 7564 35028 7616 35037
rect 10416 35096 10468 35148
rect 10692 35096 10744 35148
rect 5632 34960 5684 35012
rect 6644 35003 6696 35012
rect 6644 34969 6653 35003
rect 6653 34969 6687 35003
rect 6687 34969 6696 35003
rect 6644 34960 6696 34969
rect 6092 34892 6144 34944
rect 6828 34892 6880 34944
rect 9588 35028 9640 35080
rect 10784 35071 10836 35080
rect 10784 35037 10793 35071
rect 10793 35037 10827 35071
rect 10827 35037 10836 35071
rect 10784 35028 10836 35037
rect 10968 35071 11020 35080
rect 10968 35037 10977 35071
rect 10977 35037 11011 35071
rect 11011 35037 11020 35071
rect 10968 35028 11020 35037
rect 11980 35096 12032 35148
rect 16948 35096 17000 35148
rect 11336 35028 11388 35080
rect 12808 35071 12860 35080
rect 12808 35037 12817 35071
rect 12817 35037 12851 35071
rect 12851 35037 12860 35071
rect 12808 35028 12860 35037
rect 12992 35028 13044 35080
rect 10968 34892 11020 34944
rect 11612 34892 11664 34944
rect 12532 34892 12584 34944
rect 13544 34960 13596 35012
rect 14924 34892 14976 34944
rect 22100 35164 22152 35216
rect 20812 35096 20864 35148
rect 17316 35071 17368 35080
rect 17316 35037 17325 35071
rect 17325 35037 17359 35071
rect 17359 35037 17368 35071
rect 17316 35028 17368 35037
rect 22100 35028 22152 35080
rect 22192 35071 22244 35080
rect 22192 35037 22201 35071
rect 22201 35037 22235 35071
rect 22235 35037 22244 35071
rect 22192 35028 22244 35037
rect 23112 35028 23164 35080
rect 27528 35028 27580 35080
rect 30932 35028 30984 35080
rect 32036 35028 32088 35080
rect 32680 35096 32732 35148
rect 58164 35071 58216 35080
rect 58164 35037 58173 35071
rect 58173 35037 58207 35071
rect 58207 35037 58216 35071
rect 58164 35028 58216 35037
rect 17592 35003 17644 35012
rect 17592 34969 17626 35003
rect 17626 34969 17644 35003
rect 17592 34960 17644 34969
rect 18236 34960 18288 35012
rect 18696 34960 18748 35012
rect 21088 34960 21140 35012
rect 24768 35003 24820 35012
rect 24768 34969 24777 35003
rect 24777 34969 24811 35003
rect 24811 34969 24820 35003
rect 24768 34960 24820 34969
rect 25504 34960 25556 35012
rect 29920 35003 29972 35012
rect 29920 34969 29929 35003
rect 29929 34969 29963 35003
rect 29963 34969 29972 35003
rect 29920 34960 29972 34969
rect 19432 34892 19484 34944
rect 21548 34935 21600 34944
rect 21548 34901 21557 34935
rect 21557 34901 21591 34935
rect 21591 34901 21600 34935
rect 21548 34892 21600 34901
rect 25044 34892 25096 34944
rect 31116 34892 31168 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 6644 34688 6696 34740
rect 8484 34688 8536 34740
rect 8852 34688 8904 34740
rect 10324 34731 10376 34740
rect 10324 34697 10333 34731
rect 10333 34697 10367 34731
rect 10367 34697 10376 34731
rect 10324 34688 10376 34697
rect 10692 34688 10744 34740
rect 11704 34688 11756 34740
rect 5080 34620 5132 34672
rect 2504 34595 2556 34604
rect 2504 34561 2513 34595
rect 2513 34561 2547 34595
rect 2547 34561 2556 34595
rect 2504 34552 2556 34561
rect 2780 34595 2832 34604
rect 2780 34561 2814 34595
rect 2814 34561 2832 34595
rect 2780 34552 2832 34561
rect 5632 34552 5684 34604
rect 8300 34620 8352 34672
rect 10416 34620 10468 34672
rect 8208 34595 8260 34604
rect 8208 34561 8218 34595
rect 8218 34561 8252 34595
rect 8252 34561 8260 34595
rect 8208 34552 8260 34561
rect 8484 34595 8536 34604
rect 8484 34561 8490 34595
rect 8490 34561 8524 34595
rect 8524 34561 8536 34595
rect 8484 34552 8536 34561
rect 9680 34552 9732 34604
rect 9956 34552 10008 34604
rect 10232 34552 10284 34604
rect 7564 34484 7616 34536
rect 7748 34484 7800 34536
rect 4988 34416 5040 34468
rect 10784 34595 10836 34604
rect 10784 34561 10798 34595
rect 10798 34561 10832 34595
rect 10832 34561 10836 34595
rect 10784 34552 10836 34561
rect 10968 34595 11020 34604
rect 10968 34561 10977 34595
rect 10977 34561 11011 34595
rect 11011 34561 11020 34595
rect 10968 34552 11020 34561
rect 11612 34552 11664 34604
rect 13544 34663 13596 34672
rect 13544 34629 13553 34663
rect 13553 34629 13587 34663
rect 13587 34629 13596 34663
rect 13544 34620 13596 34629
rect 13728 34688 13780 34740
rect 16948 34731 17000 34740
rect 16948 34697 16957 34731
rect 16957 34697 16991 34731
rect 16991 34697 17000 34731
rect 16948 34688 17000 34697
rect 17592 34688 17644 34740
rect 15476 34620 15528 34672
rect 18328 34688 18380 34740
rect 18052 34620 18104 34672
rect 20168 34688 20220 34740
rect 11428 34484 11480 34536
rect 12992 34484 13044 34536
rect 16948 34552 17000 34604
rect 17868 34595 17920 34604
rect 17868 34561 17877 34595
rect 17877 34561 17911 34595
rect 17911 34561 17920 34595
rect 17868 34552 17920 34561
rect 17960 34595 18012 34604
rect 17960 34561 17969 34595
rect 17969 34561 18003 34595
rect 18003 34561 18012 34595
rect 17960 34552 18012 34561
rect 18144 34595 18196 34604
rect 18144 34561 18153 34595
rect 18153 34561 18187 34595
rect 18187 34561 18196 34595
rect 19800 34620 19852 34672
rect 18144 34552 18196 34561
rect 19248 34595 19300 34604
rect 19248 34561 19262 34595
rect 19262 34561 19296 34595
rect 19296 34561 19300 34595
rect 19248 34552 19300 34561
rect 19524 34552 19576 34604
rect 20076 34595 20128 34604
rect 20076 34561 20085 34595
rect 20085 34561 20119 34595
rect 20119 34561 20128 34595
rect 20076 34552 20128 34561
rect 3148 34348 3200 34400
rect 11244 34416 11296 34468
rect 19432 34484 19484 34536
rect 20260 34595 20312 34604
rect 20260 34561 20269 34595
rect 20269 34561 20303 34595
rect 20303 34561 20312 34595
rect 24676 34688 24728 34740
rect 25504 34731 25556 34740
rect 25504 34697 25513 34731
rect 25513 34697 25547 34731
rect 25547 34697 25556 34731
rect 25504 34688 25556 34697
rect 33784 34688 33836 34740
rect 21548 34620 21600 34672
rect 24952 34620 25004 34672
rect 20260 34552 20312 34561
rect 21916 34552 21968 34604
rect 24400 34552 24452 34604
rect 25044 34595 25096 34604
rect 25044 34561 25053 34595
rect 25053 34561 25087 34595
rect 25087 34561 25096 34595
rect 25044 34552 25096 34561
rect 30104 34620 30156 34672
rect 35716 34620 35768 34672
rect 25228 34595 25280 34604
rect 25228 34561 25237 34595
rect 25237 34561 25271 34595
rect 25271 34561 25280 34595
rect 25228 34552 25280 34561
rect 26056 34552 26108 34604
rect 20444 34484 20496 34536
rect 21548 34484 21600 34536
rect 29644 34484 29696 34536
rect 30656 34552 30708 34604
rect 31760 34552 31812 34604
rect 30196 34484 30248 34536
rect 9864 34348 9916 34400
rect 11704 34348 11756 34400
rect 27160 34416 27212 34468
rect 22836 34348 22888 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 2780 34144 2832 34196
rect 7380 34144 7432 34196
rect 10784 34144 10836 34196
rect 11244 34144 11296 34196
rect 11980 34187 12032 34196
rect 11980 34153 11989 34187
rect 11989 34153 12023 34187
rect 12023 34153 12032 34187
rect 11980 34144 12032 34153
rect 14372 34144 14424 34196
rect 2872 33983 2924 33992
rect 2872 33949 2881 33983
rect 2881 33949 2915 33983
rect 2915 33949 2924 33983
rect 2872 33940 2924 33949
rect 3148 33940 3200 33992
rect 4068 33983 4120 33992
rect 4068 33949 4077 33983
rect 4077 33949 4111 33983
rect 4111 33949 4120 33983
rect 4068 33940 4120 33949
rect 6828 34076 6880 34128
rect 9680 34076 9732 34128
rect 4344 33940 4396 33992
rect 3792 33847 3844 33856
rect 3792 33813 3801 33847
rect 3801 33813 3835 33847
rect 3835 33813 3844 33847
rect 3792 33804 3844 33813
rect 4068 33804 4120 33856
rect 4160 33804 4212 33856
rect 11704 34008 11756 34060
rect 11336 33940 11388 33992
rect 9588 33872 9640 33924
rect 11060 33872 11112 33924
rect 5724 33804 5776 33856
rect 17316 34008 17368 34060
rect 16396 33940 16448 33992
rect 17592 33940 17644 33992
rect 17868 34144 17920 34196
rect 20076 34187 20128 34196
rect 20076 34153 20085 34187
rect 20085 34153 20119 34187
rect 20119 34153 20128 34187
rect 20076 34144 20128 34153
rect 22100 34144 22152 34196
rect 27896 34144 27948 34196
rect 28356 34144 28408 34196
rect 17868 33983 17920 33992
rect 17868 33949 17877 33983
rect 17877 33949 17911 33983
rect 17911 33949 17920 33983
rect 17868 33940 17920 33949
rect 18144 33940 18196 33992
rect 19340 33940 19392 33992
rect 19800 33940 19852 33992
rect 21548 33940 21600 33992
rect 22008 33940 22060 33992
rect 24400 33983 24452 33992
rect 24400 33949 24409 33983
rect 24409 33949 24443 33983
rect 24443 33949 24452 33983
rect 24400 33940 24452 33949
rect 24584 33983 24636 33992
rect 24584 33949 24593 33983
rect 24593 33949 24627 33983
rect 24627 33949 24636 33983
rect 24584 33940 24636 33949
rect 24952 34008 25004 34060
rect 33600 34008 33652 34060
rect 14372 33872 14424 33924
rect 15568 33847 15620 33856
rect 15568 33813 15577 33847
rect 15577 33813 15611 33847
rect 15611 33813 15620 33847
rect 15568 33804 15620 33813
rect 19064 33872 19116 33924
rect 19524 33872 19576 33924
rect 22744 33915 22796 33924
rect 22744 33881 22753 33915
rect 22753 33881 22787 33915
rect 22787 33881 22796 33915
rect 22744 33872 22796 33881
rect 18512 33804 18564 33856
rect 19248 33804 19300 33856
rect 22100 33804 22152 33856
rect 23296 33872 23348 33924
rect 23756 33872 23808 33924
rect 27528 33940 27580 33992
rect 29920 33940 29972 33992
rect 30104 33940 30156 33992
rect 30748 33940 30800 33992
rect 31760 33940 31812 33992
rect 32036 33940 32088 33992
rect 33784 33983 33836 33992
rect 33784 33949 33793 33983
rect 33793 33949 33827 33983
rect 33827 33949 33836 33983
rect 33784 33940 33836 33949
rect 34612 33940 34664 33992
rect 27712 33872 27764 33924
rect 30012 33915 30064 33924
rect 30012 33881 30021 33915
rect 30021 33881 30055 33915
rect 30055 33881 30064 33915
rect 30012 33872 30064 33881
rect 32220 33915 32272 33924
rect 32220 33881 32254 33915
rect 32254 33881 32272 33915
rect 32220 33872 32272 33881
rect 35716 33940 35768 33992
rect 25044 33847 25096 33856
rect 25044 33813 25053 33847
rect 25053 33813 25087 33847
rect 25087 33813 25096 33847
rect 25044 33804 25096 33813
rect 29092 33804 29144 33856
rect 30472 33804 30524 33856
rect 33324 33847 33376 33856
rect 33324 33813 33333 33847
rect 33333 33813 33367 33847
rect 33367 33813 33376 33847
rect 33324 33804 33376 33813
rect 34980 33804 35032 33856
rect 35992 33804 36044 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4344 33643 4396 33652
rect 4344 33609 4353 33643
rect 4353 33609 4387 33643
rect 4387 33609 4396 33643
rect 4344 33600 4396 33609
rect 8208 33643 8260 33652
rect 8208 33609 8217 33643
rect 8217 33609 8251 33643
rect 8251 33609 8260 33643
rect 8208 33600 8260 33609
rect 11244 33600 11296 33652
rect 2228 33396 2280 33448
rect 6368 33532 6420 33584
rect 3792 33464 3844 33516
rect 5632 33464 5684 33516
rect 10416 33532 10468 33584
rect 15476 33532 15528 33584
rect 15568 33532 15620 33584
rect 16304 33532 16356 33584
rect 17868 33600 17920 33652
rect 19064 33643 19116 33652
rect 19064 33609 19073 33643
rect 19073 33609 19107 33643
rect 19107 33609 19116 33643
rect 19064 33600 19116 33609
rect 17592 33532 17644 33584
rect 18604 33532 18656 33584
rect 6920 33464 6972 33516
rect 12348 33464 12400 33516
rect 16488 33464 16540 33516
rect 5356 33396 5408 33448
rect 14556 33439 14608 33448
rect 14556 33405 14565 33439
rect 14565 33405 14599 33439
rect 14599 33405 14608 33439
rect 14556 33396 14608 33405
rect 15660 33396 15712 33448
rect 17960 33464 18012 33516
rect 19340 33532 19392 33584
rect 23480 33532 23532 33584
rect 24768 33600 24820 33652
rect 27712 33643 27764 33652
rect 27712 33609 27721 33643
rect 27721 33609 27755 33643
rect 27755 33609 27764 33643
rect 27712 33600 27764 33609
rect 19708 33464 19760 33516
rect 24400 33507 24452 33516
rect 17132 33396 17184 33448
rect 24400 33473 24409 33507
rect 24409 33473 24443 33507
rect 24443 33473 24452 33507
rect 24400 33464 24452 33473
rect 24952 33532 25004 33584
rect 24768 33507 24820 33516
rect 24768 33473 24777 33507
rect 24777 33473 24811 33507
rect 24811 33473 24820 33507
rect 24768 33464 24820 33473
rect 25136 33396 25188 33448
rect 27160 33464 27212 33516
rect 30564 33600 30616 33652
rect 30104 33532 30156 33584
rect 28356 33507 28408 33516
rect 28356 33473 28365 33507
rect 28365 33473 28399 33507
rect 28399 33473 28408 33507
rect 28356 33464 28408 33473
rect 29092 33464 29144 33516
rect 30196 33464 30248 33516
rect 30472 33507 30524 33516
rect 30472 33473 30476 33507
rect 30476 33473 30510 33507
rect 30510 33473 30524 33507
rect 30472 33464 30524 33473
rect 26240 33328 26292 33380
rect 30380 33396 30432 33448
rect 34152 33600 34204 33652
rect 33600 33464 33652 33516
rect 34060 33507 34112 33516
rect 34060 33473 34069 33507
rect 34069 33473 34103 33507
rect 34103 33473 34112 33507
rect 34060 33464 34112 33473
rect 31852 33396 31904 33448
rect 34428 33464 34480 33516
rect 36268 33464 36320 33516
rect 34520 33396 34572 33448
rect 34980 33396 35032 33448
rect 58164 33371 58216 33380
rect 58164 33337 58173 33371
rect 58173 33337 58207 33371
rect 58207 33337 58216 33371
rect 58164 33328 58216 33337
rect 17592 33260 17644 33312
rect 18236 33260 18288 33312
rect 19708 33303 19760 33312
rect 19708 33269 19717 33303
rect 19717 33269 19751 33303
rect 19751 33269 19760 33303
rect 19708 33260 19760 33269
rect 27160 33303 27212 33312
rect 27160 33269 27169 33303
rect 27169 33269 27203 33303
rect 27203 33269 27212 33303
rect 27160 33260 27212 33269
rect 29368 33260 29420 33312
rect 30380 33260 30432 33312
rect 30840 33260 30892 33312
rect 34520 33260 34572 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 6920 33056 6972 33108
rect 13820 33056 13872 33108
rect 18052 33056 18104 33108
rect 24584 33056 24636 33108
rect 24860 33056 24912 33108
rect 25136 33099 25188 33108
rect 25136 33065 25145 33099
rect 25145 33065 25179 33099
rect 25179 33065 25188 33099
rect 25136 33056 25188 33065
rect 15844 32988 15896 33040
rect 7932 32920 7984 32972
rect 16396 32920 16448 32972
rect 7472 32895 7524 32904
rect 7472 32861 7481 32895
rect 7481 32861 7515 32895
rect 7515 32861 7524 32895
rect 7472 32852 7524 32861
rect 8208 32852 8260 32904
rect 14096 32895 14148 32904
rect 14096 32861 14105 32895
rect 14105 32861 14139 32895
rect 14139 32861 14148 32895
rect 14096 32852 14148 32861
rect 14924 32852 14976 32904
rect 16304 32895 16356 32904
rect 16304 32861 16314 32895
rect 16314 32861 16348 32895
rect 16348 32861 16356 32895
rect 16304 32852 16356 32861
rect 16488 32895 16540 32904
rect 16488 32861 16497 32895
rect 16497 32861 16531 32895
rect 16531 32861 16540 32895
rect 16488 32852 16540 32861
rect 17132 32920 17184 32972
rect 23756 32988 23808 33040
rect 24216 32988 24268 33040
rect 32220 33056 32272 33108
rect 34060 33056 34112 33108
rect 34612 33056 34664 33108
rect 34796 33056 34848 33108
rect 30196 32988 30248 33040
rect 35900 33056 35952 33108
rect 17592 32895 17644 32904
rect 17592 32861 17622 32895
rect 17622 32861 17644 32895
rect 17592 32852 17644 32861
rect 17684 32895 17736 32904
rect 17684 32861 17693 32895
rect 17693 32861 17727 32895
rect 17727 32861 17736 32895
rect 18604 32920 18656 32972
rect 29184 32920 29236 32972
rect 23480 32895 23532 32904
rect 17684 32852 17736 32861
rect 4068 32716 4120 32768
rect 6552 32716 6604 32768
rect 7380 32716 7432 32768
rect 8208 32716 8260 32768
rect 14464 32784 14516 32836
rect 23480 32861 23489 32895
rect 23489 32861 23523 32895
rect 23523 32861 23532 32895
rect 23480 32852 23532 32861
rect 26240 32895 26292 32904
rect 26240 32861 26258 32895
rect 26258 32861 26292 32895
rect 26516 32895 26568 32904
rect 26240 32852 26292 32861
rect 26516 32861 26525 32895
rect 26525 32861 26559 32895
rect 26559 32861 26568 32895
rect 29736 32895 29788 32904
rect 26516 32852 26568 32861
rect 19708 32784 19760 32836
rect 23664 32827 23716 32836
rect 15200 32716 15252 32768
rect 17868 32716 17920 32768
rect 18420 32716 18472 32768
rect 23664 32793 23673 32827
rect 23673 32793 23707 32827
rect 23707 32793 23716 32827
rect 23664 32784 23716 32793
rect 23572 32716 23624 32768
rect 29736 32861 29745 32895
rect 29745 32861 29779 32895
rect 29779 32861 29788 32895
rect 29736 32852 29788 32861
rect 34428 32920 34480 32972
rect 29000 32784 29052 32836
rect 29276 32784 29328 32836
rect 30196 32784 30248 32836
rect 31024 32852 31076 32904
rect 31484 32852 31536 32904
rect 31300 32784 31352 32836
rect 31852 32784 31904 32836
rect 32496 32852 32548 32904
rect 33600 32852 33652 32904
rect 33784 32895 33836 32904
rect 33784 32861 33793 32895
rect 33793 32861 33827 32895
rect 33827 32861 33836 32895
rect 33784 32852 33836 32861
rect 34520 32852 34572 32904
rect 35992 32895 36044 32904
rect 35992 32861 36010 32895
rect 36010 32861 36044 32895
rect 36268 32895 36320 32904
rect 35992 32852 36044 32861
rect 36268 32861 36277 32895
rect 36277 32861 36311 32895
rect 36311 32861 36320 32895
rect 36268 32852 36320 32861
rect 27528 32716 27580 32768
rect 30656 32759 30708 32768
rect 30656 32725 30665 32759
rect 30665 32725 30699 32759
rect 30699 32725 30708 32759
rect 30656 32716 30708 32725
rect 30932 32716 30984 32768
rect 31484 32716 31536 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 7472 32512 7524 32564
rect 9772 32512 9824 32564
rect 10876 32512 10928 32564
rect 14188 32512 14240 32564
rect 14464 32555 14516 32564
rect 14464 32521 14473 32555
rect 14473 32521 14507 32555
rect 14507 32521 14516 32555
rect 14464 32512 14516 32521
rect 17316 32512 17368 32564
rect 8944 32444 8996 32496
rect 12624 32444 12676 32496
rect 13084 32444 13136 32496
rect 13452 32444 13504 32496
rect 2228 32419 2280 32428
rect 2228 32385 2237 32419
rect 2237 32385 2271 32419
rect 2271 32385 2280 32419
rect 2228 32376 2280 32385
rect 2320 32376 2372 32428
rect 6368 32419 6420 32428
rect 6368 32385 6377 32419
rect 6377 32385 6411 32419
rect 6411 32385 6420 32419
rect 6368 32376 6420 32385
rect 6460 32376 6512 32428
rect 8208 32376 8260 32428
rect 11060 32376 11112 32428
rect 12900 32376 12952 32428
rect 13820 32419 13872 32428
rect 13820 32385 13829 32419
rect 13829 32385 13863 32419
rect 13863 32385 13872 32419
rect 13820 32376 13872 32385
rect 14372 32444 14424 32496
rect 15200 32444 15252 32496
rect 15384 32444 15436 32496
rect 17592 32444 17644 32496
rect 12072 32308 12124 32360
rect 14188 32419 14240 32428
rect 14188 32385 14197 32419
rect 14197 32385 14231 32419
rect 14231 32385 14240 32419
rect 14188 32376 14240 32385
rect 14556 32376 14608 32428
rect 14924 32419 14976 32428
rect 14924 32385 14933 32419
rect 14933 32385 14967 32419
rect 14967 32385 14976 32419
rect 14924 32376 14976 32385
rect 15568 32376 15620 32428
rect 17132 32419 17184 32428
rect 17132 32385 17141 32419
rect 17141 32385 17175 32419
rect 17175 32385 17184 32419
rect 17132 32376 17184 32385
rect 18604 32512 18656 32564
rect 23664 32512 23716 32564
rect 24124 32555 24176 32564
rect 24124 32521 24133 32555
rect 24133 32521 24167 32555
rect 24167 32521 24176 32555
rect 24124 32512 24176 32521
rect 18512 32444 18564 32496
rect 25044 32444 25096 32496
rect 19248 32376 19300 32428
rect 19432 32376 19484 32428
rect 16948 32308 17000 32360
rect 17316 32308 17368 32360
rect 17592 32308 17644 32360
rect 21180 32308 21232 32360
rect 24032 32376 24084 32428
rect 26516 32376 26568 32428
rect 29736 32512 29788 32564
rect 29920 32555 29972 32564
rect 29920 32521 29929 32555
rect 29929 32521 29963 32555
rect 29963 32521 29972 32555
rect 29920 32512 29972 32521
rect 32312 32512 32364 32564
rect 36268 32555 36320 32564
rect 36268 32521 36277 32555
rect 36277 32521 36311 32555
rect 36311 32521 36320 32555
rect 36268 32512 36320 32521
rect 29092 32444 29144 32496
rect 32496 32487 32548 32496
rect 32496 32453 32505 32487
rect 32505 32453 32539 32487
rect 32539 32453 32548 32487
rect 32496 32444 32548 32453
rect 22192 32308 22244 32360
rect 28816 32376 28868 32428
rect 29644 32376 29696 32428
rect 31760 32376 31812 32428
rect 32220 32376 32272 32428
rect 33324 32376 33376 32428
rect 30196 32308 30248 32360
rect 3608 32215 3660 32224
rect 3608 32181 3617 32215
rect 3617 32181 3651 32215
rect 3651 32181 3660 32215
rect 3608 32172 3660 32181
rect 6736 32172 6788 32224
rect 17040 32240 17092 32292
rect 23480 32240 23532 32292
rect 27436 32240 27488 32292
rect 8116 32172 8168 32224
rect 10140 32172 10192 32224
rect 13360 32172 13412 32224
rect 27712 32172 27764 32224
rect 29000 32240 29052 32292
rect 30288 32240 30340 32292
rect 31208 32172 31260 32224
rect 58164 32215 58216 32224
rect 58164 32181 58173 32215
rect 58173 32181 58207 32215
rect 58207 32181 58216 32215
rect 58164 32172 58216 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2320 31968 2372 32020
rect 6368 31968 6420 32020
rect 3240 31900 3292 31952
rect 7288 31968 7340 32020
rect 11796 31968 11848 32020
rect 12072 31968 12124 32020
rect 14924 31968 14976 32020
rect 17132 31968 17184 32020
rect 20628 31968 20680 32020
rect 27160 31968 27212 32020
rect 29000 31968 29052 32020
rect 30012 31968 30064 32020
rect 11060 31900 11112 31952
rect 14188 31943 14240 31952
rect 14188 31909 14197 31943
rect 14197 31909 14231 31943
rect 14231 31909 14240 31943
rect 14188 31900 14240 31909
rect 17316 31900 17368 31952
rect 22284 31900 22336 31952
rect 28540 31900 28592 31952
rect 30748 31968 30800 32020
rect 31208 31968 31260 32020
rect 36452 31968 36504 32020
rect 36268 31900 36320 31952
rect 11428 31875 11480 31884
rect 11428 31841 11437 31875
rect 11437 31841 11471 31875
rect 11471 31841 11480 31875
rect 11428 31832 11480 31841
rect 17960 31832 18012 31884
rect 24400 31832 24452 31884
rect 24676 31832 24728 31884
rect 24952 31875 25004 31884
rect 24952 31841 24961 31875
rect 24961 31841 24995 31875
rect 24995 31841 25004 31875
rect 24952 31832 25004 31841
rect 37556 31875 37608 31884
rect 2688 31807 2740 31816
rect 2688 31773 2697 31807
rect 2697 31773 2731 31807
rect 2731 31773 2740 31807
rect 2688 31764 2740 31773
rect 4988 31764 5040 31816
rect 7288 31764 7340 31816
rect 7564 31764 7616 31816
rect 12808 31764 12860 31816
rect 16672 31764 16724 31816
rect 22100 31807 22152 31816
rect 22100 31773 22109 31807
rect 22109 31773 22143 31807
rect 22143 31773 22152 31807
rect 22100 31764 22152 31773
rect 25228 31807 25280 31816
rect 25228 31773 25237 31807
rect 25237 31773 25271 31807
rect 25271 31773 25280 31807
rect 25228 31764 25280 31773
rect 30840 31807 30892 31816
rect 30840 31773 30858 31807
rect 30858 31773 30892 31807
rect 30840 31764 30892 31773
rect 32312 31764 32364 31816
rect 36268 31807 36320 31816
rect 2780 31696 2832 31748
rect 5632 31696 5684 31748
rect 8116 31739 8168 31748
rect 8116 31705 8125 31739
rect 8125 31705 8159 31739
rect 8159 31705 8168 31739
rect 8116 31696 8168 31705
rect 9680 31696 9732 31748
rect 3332 31628 3384 31680
rect 12900 31628 12952 31680
rect 22468 31671 22520 31680
rect 22468 31637 22477 31671
rect 22477 31637 22511 31671
rect 22511 31637 22520 31671
rect 22468 31628 22520 31637
rect 22652 31696 22704 31748
rect 22836 31696 22888 31748
rect 23664 31696 23716 31748
rect 35992 31696 36044 31748
rect 36268 31773 36277 31807
rect 36277 31773 36311 31807
rect 36311 31773 36320 31807
rect 36268 31764 36320 31773
rect 36176 31696 36228 31748
rect 36452 31764 36504 31816
rect 37556 31841 37565 31875
rect 37565 31841 37599 31875
rect 37599 31841 37608 31875
rect 37556 31832 37608 31841
rect 22928 31628 22980 31680
rect 38936 31671 38988 31680
rect 38936 31637 38945 31671
rect 38945 31637 38979 31671
rect 38979 31637 38988 31671
rect 38936 31628 38988 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 2780 31424 2832 31476
rect 5264 31424 5316 31476
rect 5632 31467 5684 31476
rect 5632 31433 5641 31467
rect 5641 31433 5675 31467
rect 5675 31433 5684 31467
rect 5632 31424 5684 31433
rect 7288 31424 7340 31476
rect 9680 31467 9732 31476
rect 9680 31433 9689 31467
rect 9689 31433 9723 31467
rect 9723 31433 9732 31467
rect 9680 31424 9732 31433
rect 3608 31356 3660 31408
rect 4068 31356 4120 31408
rect 2780 31331 2832 31340
rect 2780 31297 2789 31331
rect 2789 31297 2823 31331
rect 2823 31297 2832 31331
rect 6828 31356 6880 31408
rect 2780 31288 2832 31297
rect 7104 31331 7156 31340
rect 7104 31297 7113 31331
rect 7113 31297 7147 31331
rect 7147 31297 7156 31331
rect 7104 31288 7156 31297
rect 10232 31424 10284 31476
rect 10876 31467 10928 31476
rect 10876 31433 10885 31467
rect 10885 31433 10919 31467
rect 10919 31433 10928 31467
rect 10876 31424 10928 31433
rect 12808 31424 12860 31476
rect 13268 31424 13320 31476
rect 16304 31424 16356 31476
rect 24400 31424 24452 31476
rect 5908 31220 5960 31272
rect 7472 31331 7524 31340
rect 7472 31297 7481 31331
rect 7481 31297 7515 31331
rect 7515 31297 7524 31331
rect 7472 31288 7524 31297
rect 8576 31220 8628 31272
rect 9588 31220 9640 31272
rect 10140 31331 10192 31340
rect 10140 31297 10149 31331
rect 10149 31297 10183 31331
rect 10183 31297 10192 31331
rect 10140 31288 10192 31297
rect 10784 31288 10836 31340
rect 11704 31331 11756 31340
rect 11704 31297 11713 31331
rect 11713 31297 11747 31331
rect 11747 31297 11756 31331
rect 11704 31288 11756 31297
rect 11888 31331 11940 31340
rect 11888 31297 11897 31331
rect 11897 31297 11931 31331
rect 11931 31297 11940 31331
rect 11888 31288 11940 31297
rect 13360 31331 13412 31340
rect 13360 31297 13369 31331
rect 13369 31297 13403 31331
rect 13403 31297 13412 31331
rect 13360 31288 13412 31297
rect 13728 31288 13780 31340
rect 14280 31288 14332 31340
rect 15016 31220 15068 31272
rect 13176 31152 13228 31204
rect 7656 31084 7708 31136
rect 10416 31084 10468 31136
rect 12440 31127 12492 31136
rect 12440 31093 12449 31127
rect 12449 31093 12483 31127
rect 12483 31093 12492 31127
rect 12440 31084 12492 31093
rect 13728 31084 13780 31136
rect 14924 31084 14976 31136
rect 15660 31288 15712 31340
rect 15476 31152 15528 31204
rect 15568 31084 15620 31136
rect 19432 31288 19484 31340
rect 22282 31331 22334 31340
rect 22282 31297 22293 31331
rect 22293 31297 22327 31331
rect 22327 31297 22334 31331
rect 22282 31288 22334 31297
rect 19248 31220 19300 31272
rect 20812 31220 20864 31272
rect 22468 31331 22520 31340
rect 22468 31297 22482 31331
rect 22482 31297 22516 31331
rect 22516 31297 22520 31331
rect 22468 31288 22520 31297
rect 22560 31220 22612 31272
rect 15936 31152 15988 31204
rect 24308 31356 24360 31408
rect 29552 31424 29604 31476
rect 29920 31424 29972 31476
rect 32220 31424 32272 31476
rect 36268 31424 36320 31476
rect 30932 31356 30984 31408
rect 31116 31399 31168 31408
rect 31116 31365 31125 31399
rect 31125 31365 31159 31399
rect 31159 31365 31168 31399
rect 31116 31356 31168 31365
rect 33600 31356 33652 31408
rect 38936 31356 38988 31408
rect 23664 31288 23716 31340
rect 29920 31288 29972 31340
rect 30196 31331 30248 31340
rect 30196 31297 30205 31331
rect 30205 31297 30239 31331
rect 30239 31297 30248 31331
rect 30196 31288 30248 31297
rect 30380 31288 30432 31340
rect 31208 31331 31260 31340
rect 16304 31084 16356 31136
rect 18788 31084 18840 31136
rect 31208 31297 31217 31331
rect 31217 31297 31251 31331
rect 31251 31297 31260 31331
rect 31208 31288 31260 31297
rect 31392 31331 31444 31340
rect 31392 31297 31401 31331
rect 31401 31297 31435 31331
rect 31435 31297 31444 31331
rect 31392 31288 31444 31297
rect 33140 31288 33192 31340
rect 35348 31288 35400 31340
rect 37280 31288 37332 31340
rect 33508 31220 33560 31272
rect 30104 31152 30156 31204
rect 20904 31127 20956 31136
rect 20904 31093 20913 31127
rect 20913 31093 20947 31127
rect 20947 31093 20956 31127
rect 20904 31084 20956 31093
rect 22008 31127 22060 31136
rect 22008 31093 22017 31127
rect 22017 31093 22051 31127
rect 22051 31093 22060 31127
rect 22008 31084 22060 31093
rect 23664 31084 23716 31136
rect 25412 31084 25464 31136
rect 29460 31127 29512 31136
rect 29460 31093 29469 31127
rect 29469 31093 29503 31127
rect 29503 31093 29512 31127
rect 29460 31084 29512 31093
rect 31024 31084 31076 31136
rect 31116 31084 31168 31136
rect 31944 31084 31996 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 5908 30923 5960 30932
rect 5908 30889 5917 30923
rect 5917 30889 5951 30923
rect 5951 30889 5960 30923
rect 5908 30880 5960 30889
rect 6460 30880 6512 30932
rect 7932 30880 7984 30932
rect 11796 30880 11848 30932
rect 17040 30880 17092 30932
rect 20260 30880 20312 30932
rect 6828 30812 6880 30864
rect 3792 30676 3844 30728
rect 5632 30676 5684 30728
rect 6644 30719 6696 30728
rect 6644 30685 6653 30719
rect 6653 30685 6687 30719
rect 6687 30685 6696 30719
rect 6644 30676 6696 30685
rect 7564 30744 7616 30796
rect 7104 30676 7156 30728
rect 9680 30744 9732 30796
rect 13452 30744 13504 30796
rect 11060 30676 11112 30728
rect 12900 30719 12952 30728
rect 12900 30685 12909 30719
rect 12909 30685 12943 30719
rect 12943 30685 12952 30719
rect 12900 30676 12952 30685
rect 12992 30719 13044 30728
rect 12992 30685 13025 30719
rect 13025 30685 13044 30719
rect 12992 30676 13044 30685
rect 2780 30651 2832 30660
rect 2780 30617 2789 30651
rect 2789 30617 2823 30651
rect 2823 30617 2832 30651
rect 2780 30608 2832 30617
rect 4896 30608 4948 30660
rect 6276 30608 6328 30660
rect 6920 30608 6972 30660
rect 12440 30608 12492 30660
rect 12532 30608 12584 30660
rect 14280 30812 14332 30864
rect 16764 30812 16816 30864
rect 17316 30812 17368 30864
rect 18328 30812 18380 30864
rect 19248 30812 19300 30864
rect 14096 30744 14148 30796
rect 14832 30787 14884 30796
rect 14832 30753 14841 30787
rect 14841 30753 14875 30787
rect 14875 30753 14884 30787
rect 14832 30744 14884 30753
rect 29552 30880 29604 30932
rect 24400 30855 24452 30864
rect 24400 30821 24409 30855
rect 24409 30821 24443 30855
rect 24443 30821 24452 30855
rect 24400 30812 24452 30821
rect 14924 30676 14976 30728
rect 16488 30676 16540 30728
rect 17040 30719 17092 30728
rect 17040 30685 17049 30719
rect 17049 30685 17083 30719
rect 17083 30685 17092 30719
rect 17040 30676 17092 30685
rect 16672 30651 16724 30660
rect 2596 30540 2648 30592
rect 14004 30540 14056 30592
rect 14924 30540 14976 30592
rect 16672 30617 16681 30651
rect 16681 30617 16715 30651
rect 16715 30617 16724 30651
rect 16672 30608 16724 30617
rect 20444 30676 20496 30728
rect 21732 30719 21784 30728
rect 18512 30651 18564 30660
rect 16212 30583 16264 30592
rect 16212 30549 16221 30583
rect 16221 30549 16255 30583
rect 16255 30549 16264 30583
rect 16212 30540 16264 30549
rect 17316 30540 17368 30592
rect 18512 30617 18521 30651
rect 18521 30617 18555 30651
rect 18555 30617 18564 30651
rect 18512 30608 18564 30617
rect 21732 30685 21741 30719
rect 21741 30685 21775 30719
rect 21775 30685 21784 30719
rect 21732 30676 21784 30685
rect 22008 30719 22060 30728
rect 22008 30685 22042 30719
rect 22042 30685 22060 30719
rect 22008 30676 22060 30685
rect 24676 30676 24728 30728
rect 25136 30719 25188 30728
rect 25136 30685 25145 30719
rect 25145 30685 25179 30719
rect 25179 30685 25188 30719
rect 25136 30676 25188 30685
rect 25237 30719 25289 30728
rect 27528 30787 27580 30796
rect 25237 30685 25256 30719
rect 25256 30685 25289 30719
rect 25237 30676 25289 30685
rect 27528 30753 27537 30787
rect 27537 30753 27571 30787
rect 27571 30753 27580 30787
rect 27528 30744 27580 30753
rect 30932 30880 30984 30932
rect 33784 30880 33836 30932
rect 30380 30719 30432 30728
rect 30380 30685 30389 30719
rect 30389 30685 30423 30719
rect 30423 30685 30432 30719
rect 30380 30676 30432 30685
rect 31116 30676 31168 30728
rect 31300 30744 31352 30796
rect 32312 30787 32364 30796
rect 32312 30753 32321 30787
rect 32321 30753 32355 30787
rect 32355 30753 32364 30787
rect 32312 30744 32364 30753
rect 22100 30608 22152 30660
rect 30012 30608 30064 30660
rect 18604 30540 18656 30592
rect 22192 30540 22244 30592
rect 22928 30540 22980 30592
rect 23664 30583 23716 30592
rect 23664 30549 23673 30583
rect 23673 30549 23707 30583
rect 23707 30549 23716 30583
rect 23664 30540 23716 30549
rect 24952 30540 25004 30592
rect 30196 30583 30248 30592
rect 30196 30549 30205 30583
rect 30205 30549 30239 30583
rect 30239 30549 30248 30583
rect 30196 30540 30248 30549
rect 31208 30540 31260 30592
rect 31576 30719 31628 30728
rect 31576 30685 31585 30719
rect 31585 30685 31619 30719
rect 31619 30685 31628 30719
rect 31576 30676 31628 30685
rect 34612 30676 34664 30728
rect 35716 30744 35768 30796
rect 35900 30719 35952 30728
rect 35900 30685 35909 30719
rect 35909 30685 35943 30719
rect 35943 30685 35952 30719
rect 35900 30676 35952 30685
rect 37556 30744 37608 30796
rect 58164 30719 58216 30728
rect 58164 30685 58173 30719
rect 58173 30685 58207 30719
rect 58207 30685 58216 30719
rect 58164 30676 58216 30685
rect 35348 30608 35400 30660
rect 32312 30540 32364 30592
rect 32404 30540 32456 30592
rect 32956 30540 33008 30592
rect 36176 30540 36228 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 11888 30336 11940 30388
rect 14832 30336 14884 30388
rect 4896 30268 4948 30320
rect 6368 30268 6420 30320
rect 6828 30268 6880 30320
rect 2228 30200 2280 30252
rect 2504 30200 2556 30252
rect 5264 30200 5316 30252
rect 7656 30200 7708 30252
rect 15752 30268 15804 30320
rect 16212 30268 16264 30320
rect 12348 30200 12400 30252
rect 14004 30200 14056 30252
rect 15292 30243 15344 30252
rect 15292 30209 15299 30243
rect 15299 30209 15344 30243
rect 15292 30200 15344 30209
rect 9956 30132 10008 30184
rect 16488 30200 16540 30252
rect 16672 30336 16724 30388
rect 17040 30336 17092 30388
rect 18328 30268 18380 30320
rect 17960 30243 18012 30252
rect 17960 30209 17994 30243
rect 17994 30209 18012 30243
rect 18512 30336 18564 30388
rect 19156 30336 19208 30388
rect 19432 30336 19484 30388
rect 29460 30336 29512 30388
rect 30840 30336 30892 30388
rect 31208 30336 31260 30388
rect 17960 30200 18012 30209
rect 21640 30268 21692 30320
rect 22100 30268 22152 30320
rect 24124 30268 24176 30320
rect 25136 30268 25188 30320
rect 3792 30107 3844 30116
rect 3792 30073 3801 30107
rect 3801 30073 3835 30107
rect 3835 30073 3844 30107
rect 3792 30064 3844 30073
rect 3516 29996 3568 30048
rect 6368 30039 6420 30048
rect 6368 30005 6377 30039
rect 6377 30005 6411 30039
rect 6411 30005 6420 30039
rect 6368 29996 6420 30005
rect 10784 29996 10836 30048
rect 19248 30132 19300 30184
rect 20352 30200 20404 30252
rect 20444 30200 20496 30252
rect 20904 30200 20956 30252
rect 21824 30200 21876 30252
rect 22284 30200 22336 30252
rect 22744 30243 22796 30252
rect 21640 30132 21692 30184
rect 22744 30209 22753 30243
rect 22753 30209 22787 30243
rect 22787 30209 22796 30243
rect 22744 30200 22796 30209
rect 24032 30200 24084 30252
rect 24952 30200 25004 30252
rect 25412 30243 25464 30252
rect 14004 30064 14056 30116
rect 15844 30064 15896 30116
rect 19892 30064 19944 30116
rect 21456 30064 21508 30116
rect 25412 30209 25414 30243
rect 25414 30209 25448 30243
rect 25448 30209 25464 30243
rect 25412 30200 25464 30209
rect 25504 30200 25556 30252
rect 27896 30200 27948 30252
rect 28632 30200 28684 30252
rect 30656 30268 30708 30320
rect 32220 30311 32272 30320
rect 32220 30277 32229 30311
rect 32229 30277 32263 30311
rect 32263 30277 32272 30311
rect 32220 30268 32272 30277
rect 32312 30268 32364 30320
rect 33600 30311 33652 30320
rect 33600 30277 33609 30311
rect 33609 30277 33643 30311
rect 33643 30277 33652 30311
rect 33600 30268 33652 30277
rect 34428 30336 34480 30388
rect 33968 30268 34020 30320
rect 34612 30311 34664 30320
rect 34612 30277 34621 30311
rect 34621 30277 34655 30311
rect 34655 30277 34664 30311
rect 34612 30268 34664 30277
rect 28908 30243 28960 30252
rect 28908 30209 28917 30243
rect 28917 30209 28951 30243
rect 28951 30209 28960 30243
rect 28908 30200 28960 30209
rect 30288 30200 30340 30252
rect 30564 30200 30616 30252
rect 32404 30243 32456 30252
rect 32404 30209 32413 30243
rect 32413 30209 32447 30243
rect 32447 30209 32456 30243
rect 32404 30200 32456 30209
rect 33508 30243 33560 30252
rect 33508 30209 33517 30243
rect 33517 30209 33551 30243
rect 33551 30209 33560 30243
rect 33876 30243 33928 30252
rect 33508 30200 33560 30209
rect 33876 30209 33885 30243
rect 33885 30209 33919 30243
rect 33919 30209 33928 30243
rect 33876 30200 33928 30209
rect 34336 30200 34388 30252
rect 27436 30132 27488 30184
rect 30012 30132 30064 30184
rect 34060 30132 34112 30184
rect 34796 30200 34848 30252
rect 25964 30107 26016 30116
rect 25964 30073 25973 30107
rect 25973 30073 26007 30107
rect 26007 30073 26016 30107
rect 25964 30064 26016 30073
rect 28264 30064 28316 30116
rect 31576 30064 31628 30116
rect 32220 30064 32272 30116
rect 16396 29996 16448 30048
rect 22376 29996 22428 30048
rect 25504 29996 25556 30048
rect 27896 30039 27948 30048
rect 27896 30005 27905 30039
rect 27905 30005 27939 30039
rect 27939 30005 27948 30039
rect 27896 29996 27948 30005
rect 28448 30039 28500 30048
rect 28448 30005 28457 30039
rect 28457 30005 28491 30039
rect 28491 30005 28500 30039
rect 28448 29996 28500 30005
rect 33600 29996 33652 30048
rect 34336 30039 34388 30048
rect 34336 30005 34345 30039
rect 34345 30005 34379 30039
rect 34379 30005 34388 30039
rect 34336 29996 34388 30005
rect 35900 30243 35952 30252
rect 35900 30209 35909 30243
rect 35909 30209 35943 30243
rect 35943 30209 35952 30243
rect 35900 30200 35952 30209
rect 37280 30311 37332 30320
rect 37280 30277 37289 30311
rect 37289 30277 37323 30311
rect 37323 30277 37332 30311
rect 37280 30268 37332 30277
rect 36176 30243 36228 30252
rect 36176 30209 36185 30243
rect 36185 30209 36219 30243
rect 36219 30209 36228 30243
rect 36176 30200 36228 30209
rect 36360 30200 36412 30252
rect 37464 30243 37516 30252
rect 37464 30209 37473 30243
rect 37473 30209 37507 30243
rect 37507 30209 37516 30243
rect 37464 30200 37516 30209
rect 36360 29996 36412 30048
rect 39672 29996 39724 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2504 29792 2556 29844
rect 8944 29792 8996 29844
rect 11704 29792 11756 29844
rect 11980 29835 12032 29844
rect 11980 29801 11989 29835
rect 11989 29801 12023 29835
rect 12023 29801 12032 29835
rect 11980 29792 12032 29801
rect 15476 29835 15528 29844
rect 15476 29801 15485 29835
rect 15485 29801 15519 29835
rect 15519 29801 15528 29835
rect 15476 29792 15528 29801
rect 17960 29792 18012 29844
rect 2596 29724 2648 29776
rect 2320 29588 2372 29640
rect 14188 29724 14240 29776
rect 2780 29631 2832 29640
rect 2780 29597 2789 29631
rect 2789 29597 2823 29631
rect 2823 29597 2832 29631
rect 2780 29588 2832 29597
rect 3424 29588 3476 29640
rect 3608 29588 3660 29640
rect 4712 29656 4764 29708
rect 9956 29699 10008 29708
rect 9956 29665 9965 29699
rect 9965 29665 9999 29699
rect 9999 29665 10008 29699
rect 9956 29656 10008 29665
rect 5632 29588 5684 29640
rect 9312 29631 9364 29640
rect 9312 29597 9321 29631
rect 9321 29597 9355 29631
rect 9355 29597 9364 29631
rect 9312 29588 9364 29597
rect 12164 29588 12216 29640
rect 13176 29588 13228 29640
rect 14924 29588 14976 29640
rect 15752 29588 15804 29640
rect 16948 29588 17000 29640
rect 3240 29520 3292 29572
rect 4344 29563 4396 29572
rect 4344 29529 4353 29563
rect 4353 29529 4387 29563
rect 4387 29529 4396 29563
rect 4344 29520 4396 29529
rect 7748 29520 7800 29572
rect 10692 29520 10744 29572
rect 10968 29520 11020 29572
rect 12624 29520 12676 29572
rect 18604 29588 18656 29640
rect 18880 29588 18932 29640
rect 20352 29792 20404 29844
rect 21548 29835 21600 29844
rect 21548 29801 21557 29835
rect 21557 29801 21591 29835
rect 21591 29801 21600 29835
rect 21548 29792 21600 29801
rect 23296 29792 23348 29844
rect 20812 29724 20864 29776
rect 18788 29520 18840 29572
rect 19432 29520 19484 29572
rect 19892 29520 19944 29572
rect 20352 29520 20404 29572
rect 21180 29588 21232 29640
rect 21456 29588 21508 29640
rect 22192 29631 22244 29640
rect 22192 29597 22201 29631
rect 22201 29597 22235 29631
rect 22235 29597 22244 29631
rect 22192 29588 22244 29597
rect 22284 29588 22336 29640
rect 21640 29520 21692 29572
rect 24860 29724 24912 29776
rect 24676 29631 24728 29640
rect 24676 29597 24685 29631
rect 24685 29597 24719 29631
rect 24719 29597 24728 29631
rect 24676 29588 24728 29597
rect 24860 29631 24912 29640
rect 24860 29597 24869 29631
rect 24869 29597 24903 29631
rect 24903 29597 24912 29631
rect 24860 29588 24912 29597
rect 25412 29792 25464 29844
rect 28356 29792 28408 29844
rect 28908 29792 28960 29844
rect 31300 29792 31352 29844
rect 34244 29792 34296 29844
rect 33140 29724 33192 29776
rect 27528 29656 27580 29708
rect 28264 29588 28316 29640
rect 28540 29588 28592 29640
rect 29092 29656 29144 29708
rect 29736 29631 29788 29640
rect 29736 29597 29745 29631
rect 29745 29597 29779 29631
rect 29779 29597 29788 29631
rect 29736 29588 29788 29597
rect 29828 29631 29880 29640
rect 29828 29597 29837 29631
rect 29837 29597 29871 29631
rect 29871 29597 29880 29631
rect 29828 29588 29880 29597
rect 30748 29631 30800 29640
rect 25228 29520 25280 29572
rect 29920 29563 29972 29572
rect 29920 29529 29929 29563
rect 29929 29529 29963 29563
rect 29963 29529 29972 29563
rect 29920 29520 29972 29529
rect 30380 29520 30432 29572
rect 30748 29597 30757 29631
rect 30757 29597 30791 29631
rect 30791 29597 30800 29631
rect 30748 29588 30800 29597
rect 33508 29588 33560 29640
rect 33968 29631 34020 29640
rect 33968 29597 33977 29631
rect 33977 29597 34011 29631
rect 34011 29597 34020 29631
rect 33968 29588 34020 29597
rect 34520 29588 34572 29640
rect 35348 29792 35400 29844
rect 35440 29724 35492 29776
rect 36176 29656 36228 29708
rect 37464 29588 37516 29640
rect 39304 29631 39356 29640
rect 39304 29597 39313 29631
rect 39313 29597 39347 29631
rect 39347 29597 39356 29631
rect 39304 29588 39356 29597
rect 58164 29631 58216 29640
rect 58164 29597 58173 29631
rect 58173 29597 58207 29631
rect 58207 29597 58216 29631
rect 58164 29588 58216 29597
rect 36728 29520 36780 29572
rect 4896 29452 4948 29504
rect 6920 29452 6972 29504
rect 8024 29452 8076 29504
rect 14188 29495 14240 29504
rect 14188 29461 14197 29495
rect 14197 29461 14231 29495
rect 14231 29461 14240 29495
rect 14188 29452 14240 29461
rect 22928 29452 22980 29504
rect 25044 29452 25096 29504
rect 25780 29495 25832 29504
rect 25780 29461 25789 29495
rect 25789 29461 25823 29495
rect 25823 29461 25832 29495
rect 25780 29452 25832 29461
rect 29552 29495 29604 29504
rect 29552 29461 29561 29495
rect 29561 29461 29595 29495
rect 29595 29461 29604 29495
rect 29552 29452 29604 29461
rect 33416 29452 33468 29504
rect 34152 29452 34204 29504
rect 36636 29495 36688 29504
rect 36636 29461 36645 29495
rect 36645 29461 36679 29495
rect 36679 29461 36688 29495
rect 36636 29452 36688 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 2964 29112 3016 29164
rect 3148 29155 3200 29164
rect 3148 29121 3157 29155
rect 3157 29121 3191 29155
rect 3191 29121 3200 29155
rect 3148 29112 3200 29121
rect 3516 29180 3568 29232
rect 4344 29180 4396 29232
rect 9312 29248 9364 29300
rect 10968 29291 11020 29300
rect 5540 29223 5592 29232
rect 3424 29155 3476 29164
rect 3424 29121 3433 29155
rect 3433 29121 3467 29155
rect 3467 29121 3476 29155
rect 3424 29112 3476 29121
rect 3792 29112 3844 29164
rect 5264 29155 5316 29164
rect 1952 29044 2004 29096
rect 5264 29121 5273 29155
rect 5273 29121 5307 29155
rect 5307 29121 5316 29155
rect 5264 29112 5316 29121
rect 5540 29189 5549 29223
rect 5549 29189 5583 29223
rect 5583 29189 5592 29223
rect 5540 29180 5592 29189
rect 8392 29180 8444 29232
rect 9680 29180 9732 29232
rect 10968 29257 10977 29291
rect 10977 29257 11011 29291
rect 11011 29257 11020 29291
rect 10968 29248 11020 29257
rect 18788 29291 18840 29300
rect 18788 29257 18797 29291
rect 18797 29257 18831 29291
rect 18831 29257 18840 29291
rect 18788 29248 18840 29257
rect 19248 29248 19300 29300
rect 20444 29291 20496 29300
rect 20444 29257 20453 29291
rect 20453 29257 20487 29291
rect 20487 29257 20496 29291
rect 20444 29248 20496 29257
rect 21456 29248 21508 29300
rect 24860 29248 24912 29300
rect 26056 29248 26108 29300
rect 5632 29155 5684 29164
rect 5632 29121 5641 29155
rect 5641 29121 5675 29155
rect 5675 29121 5684 29155
rect 5632 29112 5684 29121
rect 6828 29112 6880 29164
rect 9036 29112 9088 29164
rect 9864 29112 9916 29164
rect 13268 29180 13320 29232
rect 14924 29223 14976 29232
rect 13452 29155 13504 29164
rect 2780 28951 2832 28960
rect 2780 28917 2789 28951
rect 2789 28917 2823 28951
rect 2823 28917 2832 28951
rect 10416 29044 10468 29096
rect 4988 28976 5040 29028
rect 13452 29121 13461 29155
rect 13461 29121 13495 29155
rect 13495 29121 13504 29155
rect 13452 29112 13504 29121
rect 14924 29189 14933 29223
rect 14933 29189 14967 29223
rect 14967 29189 14976 29223
rect 14924 29180 14976 29189
rect 15384 29180 15436 29232
rect 23296 29180 23348 29232
rect 23388 29180 23440 29232
rect 25780 29180 25832 29232
rect 29000 29248 29052 29300
rect 30104 29248 30156 29300
rect 33140 29248 33192 29300
rect 36728 29291 36780 29300
rect 36728 29257 36737 29291
rect 36737 29257 36771 29291
rect 36771 29257 36780 29291
rect 36728 29248 36780 29257
rect 37464 29248 37516 29300
rect 34428 29180 34480 29232
rect 35440 29223 35492 29232
rect 35440 29189 35449 29223
rect 35449 29189 35483 29223
rect 35483 29189 35492 29223
rect 35440 29180 35492 29189
rect 13728 29112 13780 29164
rect 15108 29155 15160 29164
rect 15108 29121 15117 29155
rect 15117 29121 15151 29155
rect 15151 29121 15160 29155
rect 15108 29112 15160 29121
rect 19156 29112 19208 29164
rect 19340 29112 19392 29164
rect 14464 29044 14516 29096
rect 20076 29112 20128 29164
rect 21640 29112 21692 29164
rect 24032 29155 24084 29164
rect 24032 29121 24041 29155
rect 24041 29121 24075 29155
rect 24075 29121 24084 29155
rect 24032 29112 24084 29121
rect 24952 29044 25004 29096
rect 25504 29112 25556 29164
rect 13176 29019 13228 29028
rect 13176 28985 13185 29019
rect 13185 28985 13219 29019
rect 13219 28985 13228 29019
rect 13176 28976 13228 28985
rect 13452 28976 13504 29028
rect 14188 28976 14240 29028
rect 15384 28976 15436 29028
rect 18880 28976 18932 29028
rect 20352 28976 20404 29028
rect 22560 28976 22612 29028
rect 22836 28976 22888 29028
rect 25688 29019 25740 29028
rect 25688 28985 25697 29019
rect 25697 28985 25731 29019
rect 25731 28985 25740 29019
rect 25688 28976 25740 28985
rect 27620 28976 27672 29028
rect 29736 29112 29788 29164
rect 33508 29155 33560 29164
rect 33508 29121 33517 29155
rect 33517 29121 33551 29155
rect 33551 29121 33560 29155
rect 33508 29112 33560 29121
rect 35348 29112 35400 29164
rect 36084 29155 36136 29164
rect 36084 29121 36093 29155
rect 36093 29121 36127 29155
rect 36127 29121 36136 29155
rect 39672 29223 39724 29232
rect 39672 29189 39690 29223
rect 39690 29189 39724 29223
rect 39672 29180 39724 29189
rect 36084 29112 36136 29121
rect 30840 29087 30892 29096
rect 30840 29053 30849 29087
rect 30849 29053 30883 29087
rect 30883 29053 30892 29087
rect 30840 29044 30892 29053
rect 34152 29044 34204 29096
rect 36176 29044 36228 29096
rect 36636 29112 36688 29164
rect 30288 28976 30340 29028
rect 31760 28976 31812 29028
rect 2780 28908 2832 28917
rect 6644 28908 6696 28960
rect 9220 28951 9272 28960
rect 9220 28917 9229 28951
rect 9229 28917 9263 28951
rect 9263 28917 9272 28951
rect 9220 28908 9272 28917
rect 10416 28908 10468 28960
rect 15292 28951 15344 28960
rect 15292 28917 15301 28951
rect 15301 28917 15335 28951
rect 15335 28917 15344 28951
rect 15292 28908 15344 28917
rect 16212 28908 16264 28960
rect 19340 28908 19392 28960
rect 21640 28908 21692 28960
rect 26424 28951 26476 28960
rect 26424 28917 26433 28951
rect 26433 28917 26467 28951
rect 26467 28917 26476 28951
rect 26424 28908 26476 28917
rect 38752 28908 38804 28960
rect 39304 28908 39356 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2320 28704 2372 28756
rect 2872 28747 2924 28756
rect 2872 28713 2881 28747
rect 2881 28713 2915 28747
rect 2915 28713 2924 28747
rect 2872 28704 2924 28713
rect 9036 28747 9088 28756
rect 9036 28713 9045 28747
rect 9045 28713 9079 28747
rect 9079 28713 9088 28747
rect 9036 28704 9088 28713
rect 13728 28704 13780 28756
rect 14464 28747 14516 28756
rect 14464 28713 14473 28747
rect 14473 28713 14507 28747
rect 14507 28713 14516 28747
rect 14464 28704 14516 28713
rect 5632 28636 5684 28688
rect 11704 28636 11756 28688
rect 8392 28611 8444 28620
rect 8392 28577 8401 28611
rect 8401 28577 8435 28611
rect 8435 28577 8444 28611
rect 8392 28568 8444 28577
rect 9588 28568 9640 28620
rect 8300 28543 8352 28552
rect 8300 28509 8309 28543
rect 8309 28509 8343 28543
rect 8343 28509 8352 28543
rect 8300 28500 8352 28509
rect 9404 28543 9456 28552
rect 2964 28364 3016 28416
rect 4620 28364 4672 28416
rect 9404 28509 9413 28543
rect 9413 28509 9447 28543
rect 9447 28509 9456 28543
rect 9404 28500 9456 28509
rect 9496 28543 9548 28552
rect 9496 28509 9505 28543
rect 9505 28509 9539 28543
rect 9539 28509 9548 28543
rect 9496 28500 9548 28509
rect 10784 28500 10836 28552
rect 15660 28704 15712 28756
rect 19432 28704 19484 28756
rect 20444 28747 20496 28756
rect 20444 28713 20453 28747
rect 20453 28713 20487 28747
rect 20487 28713 20496 28747
rect 20444 28704 20496 28713
rect 24768 28747 24820 28756
rect 24768 28713 24777 28747
rect 24777 28713 24811 28747
rect 24811 28713 24820 28747
rect 24768 28704 24820 28713
rect 26976 28747 27028 28756
rect 26976 28713 26985 28747
rect 26985 28713 27019 28747
rect 27019 28713 27028 28747
rect 26976 28704 27028 28713
rect 29092 28704 29144 28756
rect 30840 28704 30892 28756
rect 15292 28636 15344 28688
rect 36176 28636 36228 28688
rect 30380 28611 30432 28620
rect 12532 28500 12584 28552
rect 12808 28543 12860 28552
rect 12808 28509 12817 28543
rect 12817 28509 12851 28543
rect 12851 28509 12860 28543
rect 12808 28500 12860 28509
rect 10416 28364 10468 28416
rect 14924 28543 14976 28552
rect 14924 28509 14933 28543
rect 14933 28509 14967 28543
rect 14967 28509 14976 28543
rect 14924 28500 14976 28509
rect 30380 28577 30389 28611
rect 30389 28577 30423 28611
rect 30423 28577 30432 28611
rect 30380 28568 30432 28577
rect 33968 28568 34020 28620
rect 13544 28432 13596 28484
rect 15384 28500 15436 28552
rect 15568 28500 15620 28552
rect 21456 28543 21508 28552
rect 21456 28509 21465 28543
rect 21465 28509 21499 28543
rect 21499 28509 21508 28543
rect 21640 28543 21692 28552
rect 21456 28500 21508 28509
rect 21640 28509 21649 28543
rect 21649 28509 21683 28543
rect 21683 28509 21692 28543
rect 21640 28500 21692 28509
rect 21824 28543 21876 28552
rect 21824 28509 21833 28543
rect 21833 28509 21867 28543
rect 21867 28509 21876 28543
rect 21824 28500 21876 28509
rect 26424 28543 26476 28552
rect 16212 28475 16264 28484
rect 11520 28364 11572 28416
rect 12992 28407 13044 28416
rect 12992 28373 13001 28407
rect 13001 28373 13035 28407
rect 13035 28373 13044 28407
rect 12992 28364 13044 28373
rect 13084 28364 13136 28416
rect 16212 28441 16221 28475
rect 16221 28441 16255 28475
rect 16255 28441 16264 28475
rect 16212 28432 16264 28441
rect 18236 28432 18288 28484
rect 18420 28432 18472 28484
rect 15568 28407 15620 28416
rect 15568 28373 15577 28407
rect 15577 28373 15611 28407
rect 15611 28373 15620 28407
rect 15568 28364 15620 28373
rect 20996 28364 21048 28416
rect 23572 28432 23624 28484
rect 26424 28509 26433 28543
rect 26433 28509 26467 28543
rect 26467 28509 26476 28543
rect 27160 28543 27212 28552
rect 26424 28500 26476 28509
rect 27160 28509 27169 28543
rect 27169 28509 27203 28543
rect 27203 28509 27212 28543
rect 27160 28500 27212 28509
rect 27620 28543 27672 28552
rect 27620 28509 27629 28543
rect 27629 28509 27663 28543
rect 27663 28509 27672 28543
rect 27620 28500 27672 28509
rect 28448 28500 28500 28552
rect 27068 28432 27120 28484
rect 23388 28364 23440 28416
rect 25504 28407 25556 28416
rect 25504 28373 25513 28407
rect 25513 28373 25547 28407
rect 25547 28373 25556 28407
rect 25504 28364 25556 28373
rect 26700 28364 26752 28416
rect 31576 28500 31628 28552
rect 34152 28500 34204 28552
rect 35440 28568 35492 28620
rect 35532 28500 35584 28552
rect 36084 28500 36136 28552
rect 36360 28543 36412 28552
rect 36360 28509 36369 28543
rect 36369 28509 36403 28543
rect 36403 28509 36412 28543
rect 36360 28500 36412 28509
rect 38752 28543 38804 28552
rect 34428 28432 34480 28484
rect 35992 28432 36044 28484
rect 38752 28509 38761 28543
rect 38761 28509 38795 28543
rect 38795 28509 38804 28543
rect 38752 28500 38804 28509
rect 34612 28364 34664 28416
rect 36176 28364 36228 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 5264 28160 5316 28212
rect 8484 28203 8536 28212
rect 8484 28169 8493 28203
rect 8493 28169 8527 28203
rect 8527 28169 8536 28203
rect 8484 28160 8536 28169
rect 9496 28160 9548 28212
rect 13084 28160 13136 28212
rect 2780 28135 2832 28144
rect 2780 28101 2814 28135
rect 2814 28101 2832 28135
rect 2780 28092 2832 28101
rect 6368 28092 6420 28144
rect 8944 28135 8996 28144
rect 6644 28067 6696 28076
rect 6644 28033 6653 28067
rect 6653 28033 6687 28067
rect 6687 28033 6696 28067
rect 6644 28024 6696 28033
rect 6736 28067 6788 28076
rect 6736 28033 6746 28067
rect 6746 28033 6780 28067
rect 6780 28033 6788 28067
rect 6920 28067 6972 28076
rect 6736 28024 6788 28033
rect 6920 28033 6929 28067
rect 6929 28033 6963 28067
rect 6963 28033 6972 28067
rect 6920 28024 6972 28033
rect 7472 28024 7524 28076
rect 8944 28101 8953 28135
rect 8953 28101 8987 28135
rect 8987 28101 8996 28135
rect 8944 28092 8996 28101
rect 9220 28092 9272 28144
rect 9588 28092 9640 28144
rect 11980 28092 12032 28144
rect 15108 28160 15160 28212
rect 16212 28160 16264 28212
rect 2412 27956 2464 28008
rect 9404 28024 9456 28076
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 12992 28024 13044 28076
rect 14832 28092 14884 28144
rect 22284 28135 22336 28144
rect 9312 27956 9364 28008
rect 11152 27956 11204 28008
rect 12348 27956 12400 28008
rect 14004 28067 14056 28076
rect 14004 28033 14018 28067
rect 14018 28033 14052 28067
rect 14052 28033 14056 28067
rect 14004 28024 14056 28033
rect 15568 28024 15620 28076
rect 22284 28101 22293 28135
rect 22293 28101 22327 28135
rect 22327 28101 22336 28135
rect 22284 28092 22336 28101
rect 19340 28024 19392 28076
rect 20076 28024 20128 28076
rect 21456 28024 21508 28076
rect 23756 28160 23808 28212
rect 33692 28160 33744 28212
rect 35992 28160 36044 28212
rect 36360 28203 36412 28212
rect 36360 28169 36369 28203
rect 36369 28169 36403 28203
rect 36403 28169 36412 28203
rect 36360 28160 36412 28169
rect 36176 28135 36228 28144
rect 36176 28101 36185 28135
rect 36185 28101 36219 28135
rect 36219 28101 36228 28135
rect 36176 28092 36228 28101
rect 26884 28024 26936 28076
rect 29736 28024 29788 28076
rect 9312 27820 9364 27872
rect 9864 27820 9916 27872
rect 14924 27888 14976 27940
rect 16672 27956 16724 28008
rect 30748 28024 30800 28076
rect 32772 28024 32824 28076
rect 34152 28067 34204 28076
rect 34152 28033 34161 28067
rect 34161 28033 34195 28067
rect 34195 28033 34204 28067
rect 34152 28024 34204 28033
rect 34428 28024 34480 28076
rect 34704 28024 34756 28076
rect 35348 28024 35400 28076
rect 31576 27999 31628 28008
rect 15016 27820 15068 27872
rect 17776 27888 17828 27940
rect 20076 27888 20128 27940
rect 22652 27888 22704 27940
rect 16856 27863 16908 27872
rect 16856 27829 16865 27863
rect 16865 27829 16899 27863
rect 16899 27829 16908 27863
rect 16856 27820 16908 27829
rect 17960 27820 18012 27872
rect 27896 27888 27948 27940
rect 31576 27965 31585 27999
rect 31585 27965 31619 27999
rect 31619 27965 31628 27999
rect 31576 27956 31628 27965
rect 58164 27931 58216 27940
rect 58164 27897 58173 27931
rect 58173 27897 58207 27931
rect 58207 27897 58216 27931
rect 58164 27888 58216 27897
rect 25044 27820 25096 27872
rect 29460 27863 29512 27872
rect 29460 27829 29469 27863
rect 29469 27829 29503 27863
rect 29503 27829 29512 27863
rect 29460 27820 29512 27829
rect 30012 27820 30064 27872
rect 30288 27820 30340 27872
rect 33508 27820 33560 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 11704 27616 11756 27668
rect 13544 27659 13596 27668
rect 7748 27548 7800 27600
rect 13544 27625 13553 27659
rect 13553 27625 13587 27659
rect 13587 27625 13596 27659
rect 13544 27616 13596 27625
rect 16856 27616 16908 27668
rect 14004 27548 14056 27600
rect 16764 27548 16816 27600
rect 4988 27455 5040 27464
rect 4988 27421 4997 27455
rect 4997 27421 5031 27455
rect 5031 27421 5040 27455
rect 4988 27412 5040 27421
rect 5356 27455 5408 27464
rect 3976 27344 4028 27396
rect 5356 27421 5365 27455
rect 5365 27421 5399 27455
rect 5399 27421 5408 27455
rect 5356 27412 5408 27421
rect 5448 27412 5500 27464
rect 7472 27480 7524 27532
rect 8300 27480 8352 27532
rect 6736 27412 6788 27464
rect 9496 27455 9548 27464
rect 9496 27421 9505 27455
rect 9505 27421 9539 27455
rect 9539 27421 9548 27455
rect 9496 27412 9548 27421
rect 10232 27480 10284 27532
rect 12164 27523 12216 27532
rect 12164 27489 12173 27523
rect 12173 27489 12207 27523
rect 12207 27489 12216 27523
rect 12164 27480 12216 27489
rect 29460 27616 29512 27668
rect 32772 27616 32824 27668
rect 33784 27616 33836 27668
rect 34428 27616 34480 27668
rect 35992 27659 36044 27668
rect 35992 27625 36001 27659
rect 36001 27625 36035 27659
rect 36035 27625 36044 27659
rect 35992 27616 36044 27625
rect 20260 27591 20312 27600
rect 20260 27557 20269 27591
rect 20269 27557 20303 27591
rect 20303 27557 20312 27591
rect 20260 27548 20312 27557
rect 5172 27344 5224 27396
rect 6920 27344 6972 27396
rect 7380 27387 7432 27396
rect 7380 27353 7389 27387
rect 7389 27353 7423 27387
rect 7423 27353 7432 27387
rect 7380 27344 7432 27353
rect 7472 27344 7524 27396
rect 10232 27344 10284 27396
rect 2504 27276 2556 27328
rect 3332 27276 3384 27328
rect 5632 27276 5684 27328
rect 8668 27276 8720 27328
rect 13176 27412 13228 27464
rect 12900 27344 12952 27396
rect 17040 27412 17092 27464
rect 17776 27412 17828 27464
rect 15384 27387 15436 27396
rect 15384 27353 15393 27387
rect 15393 27353 15427 27387
rect 15427 27353 15436 27387
rect 15384 27344 15436 27353
rect 15752 27344 15804 27396
rect 17500 27344 17552 27396
rect 24032 27548 24084 27600
rect 24768 27480 24820 27532
rect 24952 27412 25004 27464
rect 25044 27455 25096 27464
rect 25044 27421 25053 27455
rect 25053 27421 25087 27455
rect 25087 27421 25096 27455
rect 25228 27455 25280 27464
rect 25044 27412 25096 27421
rect 25228 27421 25237 27455
rect 25237 27421 25271 27455
rect 25271 27421 25280 27455
rect 25228 27412 25280 27421
rect 29736 27480 29788 27532
rect 21732 27344 21784 27396
rect 24032 27344 24084 27396
rect 27620 27412 27672 27464
rect 28448 27344 28500 27396
rect 30932 27412 30984 27464
rect 33140 27548 33192 27600
rect 34152 27548 34204 27600
rect 32772 27387 32824 27396
rect 32772 27353 32781 27387
rect 32781 27353 32815 27387
rect 32815 27353 32824 27387
rect 32772 27344 32824 27353
rect 32956 27455 33008 27464
rect 32956 27421 32965 27455
rect 32965 27421 32999 27455
rect 32999 27421 33008 27455
rect 32956 27412 33008 27421
rect 33232 27412 33284 27464
rect 34428 27412 34480 27464
rect 33692 27344 33744 27396
rect 24492 27319 24544 27328
rect 24492 27285 24501 27319
rect 24501 27285 24535 27319
rect 24535 27285 24544 27319
rect 24492 27276 24544 27285
rect 28540 27276 28592 27328
rect 32404 27319 32456 27328
rect 32404 27285 32413 27319
rect 32413 27285 32447 27319
rect 32447 27285 32456 27319
rect 32404 27276 32456 27285
rect 32588 27276 32640 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 3148 27072 3200 27124
rect 5080 27072 5132 27124
rect 6736 27072 6788 27124
rect 7932 27072 7984 27124
rect 9496 27115 9548 27124
rect 2504 26936 2556 26988
rect 3240 26979 3292 26988
rect 3240 26945 3249 26979
rect 3249 26945 3283 26979
rect 3283 26945 3292 26979
rect 3240 26936 3292 26945
rect 3884 26979 3936 26988
rect 3884 26945 3893 26979
rect 3893 26945 3927 26979
rect 3927 26945 3936 26979
rect 3884 26936 3936 26945
rect 4068 26979 4120 26988
rect 4068 26945 4077 26979
rect 4077 26945 4111 26979
rect 4111 26945 4120 26979
rect 4068 26936 4120 26945
rect 4896 26979 4948 26988
rect 4896 26945 4905 26979
rect 4905 26945 4939 26979
rect 4939 26945 4948 26979
rect 4896 26936 4948 26945
rect 5172 26979 5224 26988
rect 5172 26945 5181 26979
rect 5181 26945 5215 26979
rect 5215 26945 5224 26979
rect 5172 26936 5224 26945
rect 5448 26936 5500 26988
rect 6736 26936 6788 26988
rect 7196 26936 7248 26988
rect 7932 26936 7984 26988
rect 9496 27081 9505 27115
rect 9505 27081 9539 27115
rect 9539 27081 9548 27115
rect 9496 27072 9548 27081
rect 16212 27072 16264 27124
rect 17224 27072 17276 27124
rect 17776 27072 17828 27124
rect 20812 27072 20864 27124
rect 23756 27072 23808 27124
rect 29368 27072 29420 27124
rect 30932 27115 30984 27124
rect 30932 27081 30941 27115
rect 30941 27081 30975 27115
rect 30975 27081 30984 27115
rect 30932 27072 30984 27081
rect 10232 27004 10284 27056
rect 8668 26979 8720 26988
rect 8668 26945 8677 26979
rect 8677 26945 8711 26979
rect 8711 26945 8720 26979
rect 8668 26936 8720 26945
rect 9036 26936 9088 26988
rect 10876 26936 10928 26988
rect 12532 26936 12584 26988
rect 12808 26936 12860 26988
rect 17684 26936 17736 26988
rect 21732 27004 21784 27056
rect 25412 27004 25464 27056
rect 29552 27004 29604 27056
rect 31760 27004 31812 27056
rect 36084 27072 36136 27124
rect 19248 26979 19300 26988
rect 19248 26945 19282 26979
rect 19282 26945 19300 26979
rect 19248 26936 19300 26945
rect 20812 26936 20864 26988
rect 9588 26868 9640 26920
rect 11152 26868 11204 26920
rect 12900 26911 12952 26920
rect 12900 26877 12909 26911
rect 12909 26877 12943 26911
rect 12943 26877 12952 26911
rect 12900 26868 12952 26877
rect 13636 26868 13688 26920
rect 20168 26868 20220 26920
rect 20444 26868 20496 26920
rect 20904 26868 20956 26920
rect 22468 26936 22520 26988
rect 24032 26979 24084 26988
rect 24032 26945 24041 26979
rect 24041 26945 24075 26979
rect 24075 26945 24084 26979
rect 24032 26936 24084 26945
rect 25320 26979 25372 26988
rect 25320 26945 25354 26979
rect 25354 26945 25372 26979
rect 25320 26936 25372 26945
rect 26424 26936 26476 26988
rect 29644 26936 29696 26988
rect 32588 26979 32640 26988
rect 32588 26945 32597 26979
rect 32597 26945 32631 26979
rect 32631 26945 32640 26979
rect 32588 26936 32640 26945
rect 12164 26800 12216 26852
rect 21916 26800 21968 26852
rect 2780 26732 2832 26784
rect 6828 26732 6880 26784
rect 19340 26732 19392 26784
rect 20444 26732 20496 26784
rect 21180 26775 21232 26784
rect 21180 26741 21189 26775
rect 21189 26741 21223 26775
rect 21223 26741 21232 26775
rect 21180 26732 21232 26741
rect 22008 26732 22060 26784
rect 27620 26868 27672 26920
rect 30288 26868 30340 26920
rect 32772 26979 32824 26988
rect 32772 26945 32781 26979
rect 32781 26945 32815 26979
rect 32815 26945 32824 26979
rect 32772 26936 32824 26945
rect 34152 26979 34204 26988
rect 34152 26945 34161 26979
rect 34161 26945 34195 26979
rect 34195 26945 34204 26979
rect 34152 26936 34204 26945
rect 34428 26936 34480 26988
rect 34520 26936 34572 26988
rect 35440 26936 35492 26988
rect 33968 26868 34020 26920
rect 34152 26800 34204 26852
rect 23112 26732 23164 26784
rect 26240 26732 26292 26784
rect 29276 26775 29328 26784
rect 29276 26741 29285 26775
rect 29285 26741 29319 26775
rect 29319 26741 29328 26775
rect 29276 26732 29328 26741
rect 33232 26732 33284 26784
rect 34520 26775 34572 26784
rect 34520 26741 34529 26775
rect 34529 26741 34563 26775
rect 34563 26741 34572 26775
rect 34520 26732 34572 26741
rect 39948 26732 40000 26784
rect 58164 26775 58216 26784
rect 58164 26741 58173 26775
rect 58173 26741 58207 26775
rect 58207 26741 58216 26775
rect 58164 26732 58216 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3976 26460 4028 26512
rect 2872 26367 2924 26376
rect 2872 26333 2881 26367
rect 2881 26333 2915 26367
rect 2915 26333 2924 26367
rect 2872 26324 2924 26333
rect 2872 26188 2924 26240
rect 3240 26367 3292 26376
rect 3240 26333 3249 26367
rect 3249 26333 3283 26367
rect 3283 26333 3292 26367
rect 3240 26324 3292 26333
rect 4068 26324 4120 26376
rect 7380 26528 7432 26580
rect 9680 26528 9732 26580
rect 12348 26528 12400 26580
rect 17500 26528 17552 26580
rect 19248 26528 19300 26580
rect 22468 26571 22520 26580
rect 6920 26460 6972 26512
rect 7656 26460 7708 26512
rect 10600 26460 10652 26512
rect 22468 26537 22477 26571
rect 22477 26537 22511 26571
rect 22511 26537 22520 26571
rect 22468 26528 22520 26537
rect 24676 26528 24728 26580
rect 25320 26571 25372 26580
rect 6736 26324 6788 26376
rect 9772 26392 9824 26444
rect 5632 26256 5684 26308
rect 3148 26188 3200 26240
rect 3608 26188 3660 26240
rect 6184 26299 6236 26308
rect 6184 26265 6193 26299
rect 6193 26265 6227 26299
rect 6227 26265 6236 26299
rect 7472 26324 7524 26376
rect 7932 26324 7984 26376
rect 9404 26367 9456 26376
rect 9404 26333 9413 26367
rect 9413 26333 9447 26367
rect 9447 26333 9456 26367
rect 9404 26324 9456 26333
rect 9588 26367 9640 26376
rect 9588 26333 9597 26367
rect 9597 26333 9631 26367
rect 9631 26333 9640 26367
rect 9588 26324 9640 26333
rect 6184 26256 6236 26265
rect 8116 26256 8168 26308
rect 8208 26256 8260 26308
rect 10324 26324 10376 26376
rect 16764 26392 16816 26444
rect 24308 26460 24360 26512
rect 25044 26460 25096 26512
rect 10876 26256 10928 26308
rect 16580 26324 16632 26376
rect 14096 26256 14148 26308
rect 17040 26367 17092 26376
rect 17040 26333 17049 26367
rect 17049 26333 17083 26367
rect 17083 26333 17092 26367
rect 17040 26324 17092 26333
rect 17776 26324 17828 26376
rect 18236 26367 18288 26376
rect 17316 26256 17368 26308
rect 18236 26333 18245 26367
rect 18245 26333 18279 26367
rect 18279 26333 18288 26367
rect 18236 26324 18288 26333
rect 18144 26256 18196 26308
rect 6276 26188 6328 26240
rect 6552 26188 6604 26240
rect 18052 26188 18104 26240
rect 18696 26324 18748 26376
rect 21824 26367 21876 26376
rect 20812 26299 20864 26308
rect 20812 26265 20821 26299
rect 20821 26265 20855 26299
rect 20855 26265 20864 26299
rect 20812 26256 20864 26265
rect 21824 26333 21833 26367
rect 21833 26333 21867 26367
rect 21867 26333 21876 26367
rect 21824 26324 21876 26333
rect 21987 26367 22039 26376
rect 21987 26333 21996 26367
rect 21996 26333 22030 26367
rect 22030 26333 22039 26367
rect 21987 26324 22039 26333
rect 22100 26367 22152 26376
rect 22100 26333 22109 26367
rect 22109 26333 22143 26367
rect 22143 26333 22152 26367
rect 24492 26392 24544 26444
rect 25320 26537 25329 26571
rect 25329 26537 25363 26571
rect 25363 26537 25372 26571
rect 25320 26528 25372 26537
rect 26424 26571 26476 26580
rect 26424 26537 26433 26571
rect 26433 26537 26467 26571
rect 26467 26537 26476 26571
rect 26424 26528 26476 26537
rect 29460 26528 29512 26580
rect 29644 26571 29696 26580
rect 29644 26537 29653 26571
rect 29653 26537 29687 26571
rect 29687 26537 29696 26571
rect 29644 26528 29696 26537
rect 30104 26571 30156 26580
rect 30104 26537 30113 26571
rect 30113 26537 30147 26571
rect 30147 26537 30156 26571
rect 30104 26528 30156 26537
rect 33968 26528 34020 26580
rect 32220 26503 32272 26512
rect 32220 26469 32229 26503
rect 32229 26469 32263 26503
rect 32263 26469 32272 26503
rect 32220 26460 32272 26469
rect 32772 26460 32824 26512
rect 35440 26528 35492 26580
rect 22100 26324 22152 26333
rect 24676 26367 24728 26376
rect 24676 26333 24685 26367
rect 24685 26333 24719 26367
rect 24719 26333 24728 26367
rect 24676 26324 24728 26333
rect 24860 26367 24912 26376
rect 24860 26333 24869 26367
rect 24869 26333 24903 26367
rect 24903 26333 24912 26367
rect 24860 26324 24912 26333
rect 22468 26256 22520 26308
rect 22100 26188 22152 26240
rect 24768 26188 24820 26240
rect 25688 26324 25740 26376
rect 26976 26324 27028 26376
rect 32956 26367 33008 26376
rect 32956 26333 32965 26367
rect 32965 26333 32999 26367
rect 32999 26333 33008 26367
rect 32956 26324 33008 26333
rect 36912 26460 36964 26512
rect 33784 26392 33836 26444
rect 33876 26435 33928 26444
rect 33876 26401 33885 26435
rect 33885 26401 33919 26435
rect 33919 26401 33928 26435
rect 33876 26392 33928 26401
rect 34428 26392 34480 26444
rect 33324 26367 33376 26376
rect 33324 26333 33333 26367
rect 33333 26333 33367 26367
rect 33367 26333 33376 26367
rect 33324 26324 33376 26333
rect 34520 26324 34572 26376
rect 37096 26324 37148 26376
rect 38752 26324 38804 26376
rect 39948 26324 40000 26376
rect 26332 26256 26384 26308
rect 29276 26256 29328 26308
rect 39764 26256 39816 26308
rect 39856 26299 39908 26308
rect 39856 26265 39865 26299
rect 39865 26265 39899 26299
rect 39899 26265 39908 26299
rect 39856 26256 39908 26265
rect 32772 26231 32824 26240
rect 32772 26197 32781 26231
rect 32781 26197 32815 26231
rect 32815 26197 32824 26231
rect 32772 26188 32824 26197
rect 40408 26188 40460 26240
rect 40776 26231 40828 26240
rect 40776 26197 40785 26231
rect 40785 26197 40819 26231
rect 40819 26197 40828 26231
rect 40776 26188 40828 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 3976 26027 4028 26036
rect 3976 25993 3985 26027
rect 3985 25993 4019 26027
rect 4019 25993 4028 26027
rect 3976 25984 4028 25993
rect 6368 25984 6420 26036
rect 8208 25984 8260 26036
rect 9036 26027 9088 26036
rect 9036 25993 9045 26027
rect 9045 25993 9079 26027
rect 9079 25993 9088 26027
rect 10600 26027 10652 26036
rect 9036 25984 9088 25993
rect 10600 25993 10609 26027
rect 10609 25993 10643 26027
rect 10643 25993 10652 26027
rect 10600 25984 10652 25993
rect 13452 25984 13504 26036
rect 17684 26027 17736 26036
rect 17684 25993 17693 26027
rect 17693 25993 17727 26027
rect 17727 25993 17736 26027
rect 17684 25984 17736 25993
rect 18236 25984 18288 26036
rect 2872 25959 2924 25968
rect 2872 25925 2906 25959
rect 2906 25925 2924 25959
rect 2872 25916 2924 25925
rect 6092 25916 6144 25968
rect 10324 25916 10376 25968
rect 6368 25891 6420 25900
rect 6368 25857 6377 25891
rect 6377 25857 6411 25891
rect 6411 25857 6420 25891
rect 6368 25848 6420 25857
rect 6552 25891 6604 25900
rect 6552 25857 6561 25891
rect 6561 25857 6595 25891
rect 6595 25857 6604 25891
rect 6552 25848 6604 25857
rect 2412 25780 2464 25832
rect 3608 25780 3660 25832
rect 6736 25891 6788 25900
rect 6736 25857 6745 25891
rect 6745 25857 6779 25891
rect 6779 25857 6788 25891
rect 6736 25848 6788 25857
rect 12808 25848 12860 25900
rect 14096 25848 14148 25900
rect 15752 25891 15804 25900
rect 15752 25857 15761 25891
rect 15761 25857 15795 25891
rect 15795 25857 15804 25891
rect 15752 25848 15804 25857
rect 17500 25848 17552 25900
rect 18420 25916 18472 25968
rect 18604 25916 18656 25968
rect 18052 25891 18104 25900
rect 18052 25857 18061 25891
rect 18061 25857 18095 25891
rect 18095 25857 18104 25891
rect 18052 25848 18104 25857
rect 7840 25780 7892 25832
rect 9404 25780 9456 25832
rect 13820 25780 13872 25832
rect 13912 25780 13964 25832
rect 21824 25984 21876 26036
rect 25228 25984 25280 26036
rect 26976 26027 27028 26036
rect 20444 25916 20496 25968
rect 19248 25848 19300 25900
rect 19432 25848 19484 25900
rect 11336 25712 11388 25764
rect 16028 25712 16080 25764
rect 19248 25712 19300 25764
rect 20904 25891 20956 25900
rect 20904 25857 20913 25891
rect 20913 25857 20947 25891
rect 20947 25857 20956 25891
rect 20904 25848 20956 25857
rect 21640 25848 21692 25900
rect 21824 25891 21876 25900
rect 21824 25857 21833 25891
rect 21833 25857 21867 25891
rect 21867 25857 21876 25891
rect 21824 25848 21876 25857
rect 22468 25916 22520 25968
rect 25688 25916 25740 25968
rect 22100 25891 22152 25900
rect 22100 25857 22109 25891
rect 22109 25857 22143 25891
rect 22143 25857 22152 25891
rect 22100 25848 22152 25857
rect 26976 25993 26985 26027
rect 26985 25993 27019 26027
rect 27019 25993 27028 26027
rect 26976 25984 27028 25993
rect 30104 25984 30156 26036
rect 31576 25984 31628 26036
rect 32772 25984 32824 26036
rect 33692 25984 33744 26036
rect 26332 25916 26384 25968
rect 33232 25959 33284 25968
rect 33232 25925 33266 25959
rect 33266 25925 33284 25959
rect 33232 25916 33284 25925
rect 28540 25848 28592 25900
rect 28632 25848 28684 25900
rect 40592 25891 40644 25900
rect 24124 25780 24176 25832
rect 31300 25780 31352 25832
rect 39948 25823 40000 25832
rect 25504 25712 25556 25764
rect 31208 25712 31260 25764
rect 7012 25687 7064 25696
rect 7012 25653 7021 25687
rect 7021 25653 7055 25687
rect 7055 25653 7064 25687
rect 7012 25644 7064 25653
rect 12808 25644 12860 25696
rect 15568 25644 15620 25696
rect 22468 25687 22520 25696
rect 22468 25653 22477 25687
rect 22477 25653 22511 25687
rect 22511 25653 22520 25687
rect 22468 25644 22520 25653
rect 27620 25644 27672 25696
rect 30748 25644 30800 25696
rect 39948 25789 39957 25823
rect 39957 25789 39991 25823
rect 39991 25789 40000 25823
rect 39948 25780 40000 25789
rect 40592 25857 40601 25891
rect 40601 25857 40635 25891
rect 40635 25857 40644 25891
rect 40592 25848 40644 25857
rect 40500 25780 40552 25832
rect 37280 25712 37332 25764
rect 38568 25755 38620 25764
rect 38568 25721 38577 25755
rect 38577 25721 38611 25755
rect 38611 25721 38620 25755
rect 38568 25712 38620 25721
rect 40224 25712 40276 25764
rect 40776 25891 40828 25900
rect 40776 25857 40785 25891
rect 40785 25857 40819 25891
rect 40819 25857 40828 25891
rect 40776 25848 40828 25857
rect 33140 25644 33192 25696
rect 36360 25644 36412 25696
rect 37372 25687 37424 25696
rect 37372 25653 37381 25687
rect 37381 25653 37415 25687
rect 37415 25653 37424 25687
rect 37372 25644 37424 25653
rect 39304 25644 39356 25696
rect 40592 25644 40644 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 6184 25440 6236 25492
rect 8576 25440 8628 25492
rect 18052 25440 18104 25492
rect 2412 25236 2464 25288
rect 6368 25279 6420 25288
rect 6368 25245 6377 25279
rect 6377 25245 6411 25279
rect 6411 25245 6420 25279
rect 6368 25236 6420 25245
rect 7012 25236 7064 25288
rect 8576 25236 8628 25288
rect 17960 25372 18012 25424
rect 18236 25372 18288 25424
rect 9956 25304 10008 25356
rect 10324 25304 10376 25356
rect 11060 25304 11112 25356
rect 12164 25304 12216 25356
rect 9772 25236 9824 25288
rect 9864 25279 9916 25288
rect 9864 25245 9873 25279
rect 9873 25245 9907 25279
rect 9907 25245 9916 25279
rect 9864 25236 9916 25245
rect 5908 25211 5960 25220
rect 5908 25177 5917 25211
rect 5917 25177 5951 25211
rect 5951 25177 5960 25211
rect 5908 25168 5960 25177
rect 7288 25168 7340 25220
rect 13360 25236 13412 25288
rect 15936 25236 15988 25288
rect 8576 25100 8628 25152
rect 14096 25143 14148 25152
rect 14096 25109 14105 25143
rect 14105 25109 14139 25143
rect 14139 25109 14148 25143
rect 14096 25100 14148 25109
rect 14832 25100 14884 25152
rect 15568 25168 15620 25220
rect 16028 25168 16080 25220
rect 16948 25211 17000 25220
rect 16948 25177 16957 25211
rect 16957 25177 16991 25211
rect 16991 25177 17000 25211
rect 16948 25168 17000 25177
rect 18144 25236 18196 25288
rect 24860 25440 24912 25492
rect 31300 25483 31352 25492
rect 31300 25449 31309 25483
rect 31309 25449 31343 25483
rect 31343 25449 31352 25483
rect 31300 25440 31352 25449
rect 39304 25483 39356 25492
rect 39304 25449 39313 25483
rect 39313 25449 39347 25483
rect 39347 25449 39356 25483
rect 39304 25440 39356 25449
rect 39764 25440 39816 25492
rect 29828 25372 29880 25424
rect 30380 25372 30432 25424
rect 19340 25236 19392 25288
rect 21732 25236 21784 25288
rect 24952 25236 25004 25288
rect 26332 25236 26384 25288
rect 29828 25279 29880 25288
rect 29828 25245 29837 25279
rect 29837 25245 29871 25279
rect 29871 25245 29880 25279
rect 29828 25236 29880 25245
rect 20168 25168 20220 25220
rect 22468 25168 22520 25220
rect 26240 25168 26292 25220
rect 29736 25168 29788 25220
rect 30656 25236 30708 25288
rect 15844 25100 15896 25152
rect 18604 25100 18656 25152
rect 19156 25100 19208 25152
rect 19340 25143 19392 25152
rect 19340 25109 19349 25143
rect 19349 25109 19383 25143
rect 19383 25109 19392 25143
rect 19340 25100 19392 25109
rect 20444 25100 20496 25152
rect 21640 25143 21692 25152
rect 21640 25109 21649 25143
rect 21649 25109 21683 25143
rect 21683 25109 21692 25143
rect 21640 25100 21692 25109
rect 22836 25100 22888 25152
rect 28264 25100 28316 25152
rect 29644 25100 29696 25152
rect 30012 25100 30064 25152
rect 37096 25347 37148 25356
rect 37096 25313 37105 25347
rect 37105 25313 37139 25347
rect 37139 25313 37148 25347
rect 37096 25304 37148 25313
rect 40224 25440 40276 25492
rect 33140 25236 33192 25288
rect 34060 25236 34112 25288
rect 37372 25236 37424 25288
rect 38936 25279 38988 25288
rect 32036 25168 32088 25220
rect 37648 25168 37700 25220
rect 32496 25100 32548 25152
rect 35624 25100 35676 25152
rect 38936 25245 38945 25279
rect 38945 25245 38979 25279
rect 38979 25245 38988 25279
rect 38936 25236 38988 25245
rect 39856 25236 39908 25288
rect 40132 25279 40184 25288
rect 40132 25245 40141 25279
rect 40141 25245 40175 25279
rect 40175 25245 40184 25279
rect 40132 25236 40184 25245
rect 58164 25279 58216 25288
rect 38568 25168 38620 25220
rect 40408 25168 40460 25220
rect 58164 25245 58173 25279
rect 58173 25245 58207 25279
rect 58207 25245 58216 25279
rect 58164 25236 58216 25245
rect 40500 25100 40552 25152
rect 40868 25100 40920 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 3884 24939 3936 24948
rect 3884 24905 3893 24939
rect 3893 24905 3927 24939
rect 3927 24905 3936 24939
rect 3884 24896 3936 24905
rect 5908 24896 5960 24948
rect 7288 24896 7340 24948
rect 2780 24803 2832 24812
rect 2780 24769 2814 24803
rect 2814 24769 2832 24803
rect 2780 24760 2832 24769
rect 5724 24760 5776 24812
rect 7196 24760 7248 24812
rect 9036 24803 9088 24812
rect 9036 24769 9045 24803
rect 9045 24769 9079 24803
rect 9079 24769 9088 24803
rect 9036 24760 9088 24769
rect 9588 24760 9640 24812
rect 2412 24692 2464 24744
rect 10324 24803 10376 24812
rect 7196 24624 7248 24676
rect 9680 24599 9732 24608
rect 9680 24565 9689 24599
rect 9689 24565 9723 24599
rect 9723 24565 9732 24599
rect 9680 24556 9732 24565
rect 9956 24624 10008 24676
rect 10324 24769 10333 24803
rect 10333 24769 10367 24803
rect 10367 24769 10376 24803
rect 10324 24760 10376 24769
rect 13728 24803 13780 24812
rect 12440 24692 12492 24744
rect 13728 24769 13737 24803
rect 13737 24769 13771 24803
rect 13771 24769 13780 24803
rect 13728 24760 13780 24769
rect 14372 24760 14424 24812
rect 16580 24760 16632 24812
rect 19156 24803 19208 24812
rect 19156 24769 19190 24803
rect 19190 24769 19208 24803
rect 19156 24760 19208 24769
rect 27528 24896 27580 24948
rect 32404 24896 32456 24948
rect 32496 24896 32548 24948
rect 40132 24896 40184 24948
rect 40868 24896 40920 24948
rect 21732 24760 21784 24812
rect 22100 24760 22152 24812
rect 22744 24803 22796 24812
rect 22744 24769 22753 24803
rect 22753 24769 22787 24803
rect 22787 24769 22796 24803
rect 22744 24760 22796 24769
rect 22836 24803 22888 24812
rect 22836 24769 22881 24803
rect 22881 24769 22888 24803
rect 22836 24760 22888 24769
rect 23020 24803 23072 24812
rect 23020 24769 23029 24803
rect 23029 24769 23063 24803
rect 23063 24769 23072 24803
rect 23020 24760 23072 24769
rect 14188 24692 14240 24744
rect 10140 24624 10192 24676
rect 12624 24624 12676 24676
rect 12256 24556 12308 24608
rect 13176 24556 13228 24608
rect 17776 24692 17828 24744
rect 15200 24556 15252 24608
rect 16488 24624 16540 24676
rect 15844 24599 15896 24608
rect 15844 24565 15853 24599
rect 15853 24565 15887 24599
rect 15887 24565 15896 24599
rect 15844 24556 15896 24565
rect 16304 24556 16356 24608
rect 20904 24692 20956 24744
rect 24676 24760 24728 24812
rect 25044 24803 25096 24812
rect 25044 24769 25053 24803
rect 25053 24769 25087 24803
rect 25087 24769 25096 24803
rect 25044 24760 25096 24769
rect 24768 24692 24820 24744
rect 19892 24624 19944 24676
rect 18512 24556 18564 24608
rect 20076 24556 20128 24608
rect 20444 24624 20496 24676
rect 21640 24624 21692 24676
rect 27988 24828 28040 24880
rect 29000 24828 29052 24880
rect 29736 24828 29788 24880
rect 30104 24760 30156 24812
rect 30656 24803 30708 24812
rect 30656 24769 30665 24803
rect 30665 24769 30699 24803
rect 30699 24769 30708 24803
rect 30656 24760 30708 24769
rect 30748 24760 30800 24812
rect 21548 24556 21600 24608
rect 22192 24556 22244 24608
rect 25504 24599 25556 24608
rect 25504 24565 25513 24599
rect 25513 24565 25547 24599
rect 25547 24565 25556 24599
rect 25504 24556 25556 24565
rect 28264 24599 28316 24608
rect 28264 24565 28273 24599
rect 28273 24565 28307 24599
rect 28307 24565 28316 24599
rect 28264 24556 28316 24565
rect 28816 24599 28868 24608
rect 28816 24565 28825 24599
rect 28825 24565 28859 24599
rect 28859 24565 28868 24599
rect 28816 24556 28868 24565
rect 28908 24556 28960 24608
rect 32036 24692 32088 24744
rect 33968 24803 34020 24812
rect 33968 24769 33977 24803
rect 33977 24769 34011 24803
rect 34011 24769 34020 24803
rect 33968 24760 34020 24769
rect 35716 24735 35768 24744
rect 35716 24701 35725 24735
rect 35725 24701 35759 24735
rect 35759 24701 35768 24735
rect 35716 24692 35768 24701
rect 35624 24624 35676 24676
rect 38936 24760 38988 24812
rect 39764 24803 39816 24812
rect 39764 24769 39782 24803
rect 39782 24769 39816 24803
rect 39764 24760 39816 24769
rect 39948 24760 40000 24812
rect 37648 24735 37700 24744
rect 37648 24701 37657 24735
rect 37657 24701 37691 24735
rect 37691 24701 37700 24735
rect 37648 24692 37700 24701
rect 33876 24556 33928 24608
rect 36084 24556 36136 24608
rect 38660 24599 38712 24608
rect 38660 24565 38669 24599
rect 38669 24565 38703 24599
rect 38703 24565 38712 24599
rect 38660 24556 38712 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 9956 24352 10008 24404
rect 11888 24352 11940 24404
rect 14372 24395 14424 24404
rect 14372 24361 14381 24395
rect 14381 24361 14415 24395
rect 14415 24361 14424 24395
rect 14372 24352 14424 24361
rect 11060 24216 11112 24268
rect 13544 24284 13596 24336
rect 13728 24284 13780 24336
rect 15568 24284 15620 24336
rect 9680 24148 9732 24200
rect 11244 24148 11296 24200
rect 11888 24191 11940 24200
rect 11888 24157 11897 24191
rect 11897 24157 11931 24191
rect 11931 24157 11940 24191
rect 11888 24148 11940 24157
rect 12072 24191 12124 24200
rect 12072 24157 12081 24191
rect 12081 24157 12115 24191
rect 12115 24157 12124 24191
rect 12072 24148 12124 24157
rect 12256 24191 12308 24200
rect 12256 24157 12265 24191
rect 12265 24157 12299 24191
rect 12299 24157 12308 24191
rect 12256 24148 12308 24157
rect 12440 24148 12492 24200
rect 13912 24216 13964 24268
rect 13176 24191 13228 24200
rect 13176 24157 13185 24191
rect 13185 24157 13219 24191
rect 13219 24157 13228 24191
rect 13176 24148 13228 24157
rect 13360 24191 13412 24200
rect 13360 24157 13369 24191
rect 13369 24157 13403 24191
rect 13403 24157 13412 24191
rect 14648 24191 14700 24200
rect 13360 24148 13412 24157
rect 14648 24157 14657 24191
rect 14657 24157 14691 24191
rect 14691 24157 14700 24191
rect 14648 24148 14700 24157
rect 14832 24191 14884 24200
rect 14832 24157 14846 24191
rect 14846 24157 14880 24191
rect 14880 24157 14884 24191
rect 14832 24148 14884 24157
rect 15936 24352 15988 24404
rect 18236 24352 18288 24404
rect 16948 24284 17000 24336
rect 20904 24284 20956 24336
rect 18052 24216 18104 24268
rect 18420 24191 18472 24200
rect 18420 24157 18429 24191
rect 18429 24157 18463 24191
rect 18463 24157 18472 24191
rect 18420 24148 18472 24157
rect 19892 24148 19944 24200
rect 21916 24284 21968 24336
rect 21548 24216 21600 24268
rect 7840 24123 7892 24132
rect 7840 24089 7849 24123
rect 7849 24089 7883 24123
rect 7883 24089 7892 24123
rect 7840 24080 7892 24089
rect 10140 24080 10192 24132
rect 9036 24012 9088 24064
rect 9956 24012 10008 24064
rect 11244 24012 11296 24064
rect 11612 24055 11664 24064
rect 11612 24021 11621 24055
rect 11621 24021 11655 24055
rect 11655 24021 11664 24055
rect 11612 24012 11664 24021
rect 12900 24012 12952 24064
rect 13912 24012 13964 24064
rect 18236 24080 18288 24132
rect 19248 24080 19300 24132
rect 21456 24191 21508 24200
rect 21456 24157 21465 24191
rect 21465 24157 21499 24191
rect 21499 24157 21508 24191
rect 21456 24148 21508 24157
rect 16580 24055 16632 24064
rect 16580 24021 16589 24055
rect 16589 24021 16623 24055
rect 16623 24021 16632 24055
rect 16580 24012 16632 24021
rect 20904 24012 20956 24064
rect 21272 24080 21324 24132
rect 21456 24012 21508 24064
rect 22100 24148 22152 24200
rect 22560 24284 22612 24336
rect 21916 24055 21968 24064
rect 21916 24021 21925 24055
rect 21925 24021 21959 24055
rect 21959 24021 21968 24055
rect 21916 24012 21968 24021
rect 22744 24080 22796 24132
rect 24124 24012 24176 24064
rect 25044 24352 25096 24404
rect 26792 24352 26844 24404
rect 30012 24352 30064 24404
rect 30104 24352 30156 24404
rect 28264 24284 28316 24336
rect 30656 24327 30708 24336
rect 27804 24216 27856 24268
rect 28632 24216 28684 24268
rect 24952 24191 25004 24200
rect 24952 24157 24961 24191
rect 24961 24157 24995 24191
rect 24995 24157 25004 24191
rect 24952 24148 25004 24157
rect 25412 24191 25464 24200
rect 25412 24157 25421 24191
rect 25421 24157 25455 24191
rect 25455 24157 25464 24191
rect 25412 24148 25464 24157
rect 27620 24148 27672 24200
rect 28816 24191 28868 24200
rect 25504 24080 25556 24132
rect 28816 24157 28825 24191
rect 28825 24157 28859 24191
rect 28859 24157 28868 24191
rect 28816 24148 28868 24157
rect 30656 24293 30665 24327
rect 30665 24293 30699 24327
rect 30699 24293 30708 24327
rect 30656 24284 30708 24293
rect 29092 24216 29144 24268
rect 38660 24216 38712 24268
rect 27804 24123 27856 24132
rect 27804 24089 27813 24123
rect 27813 24089 27847 24123
rect 27847 24089 27856 24123
rect 27804 24080 27856 24089
rect 27988 24123 28040 24132
rect 27988 24089 27997 24123
rect 27997 24089 28031 24123
rect 28031 24089 28040 24123
rect 28632 24123 28684 24132
rect 27988 24080 28040 24089
rect 28632 24089 28641 24123
rect 28641 24089 28675 24123
rect 28675 24089 28684 24123
rect 28632 24080 28684 24089
rect 41052 24191 41104 24200
rect 26792 24055 26844 24064
rect 26792 24021 26801 24055
rect 26801 24021 26835 24055
rect 26835 24021 26844 24055
rect 26792 24012 26844 24021
rect 28172 24012 28224 24064
rect 41052 24157 41061 24191
rect 41061 24157 41095 24191
rect 41095 24157 41104 24191
rect 41052 24148 41104 24157
rect 58164 24191 58216 24200
rect 58164 24157 58173 24191
rect 58173 24157 58207 24191
rect 58207 24157 58216 24191
rect 58164 24148 58216 24157
rect 39856 24080 39908 24132
rect 29920 24012 29972 24064
rect 40408 24055 40460 24064
rect 40408 24021 40417 24055
rect 40417 24021 40451 24055
rect 40451 24021 40460 24055
rect 40408 24012 40460 24021
rect 41144 24012 41196 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 9772 23808 9824 23860
rect 12072 23808 12124 23860
rect 2228 23715 2280 23724
rect 2228 23681 2237 23715
rect 2237 23681 2271 23715
rect 2271 23681 2280 23715
rect 2228 23672 2280 23681
rect 3240 23672 3292 23724
rect 7840 23672 7892 23724
rect 11060 23740 11112 23792
rect 13728 23808 13780 23860
rect 14188 23851 14240 23860
rect 14188 23817 14197 23851
rect 14197 23817 14231 23851
rect 14231 23817 14240 23851
rect 14188 23808 14240 23817
rect 14648 23851 14700 23860
rect 14648 23817 14657 23851
rect 14657 23817 14691 23851
rect 14691 23817 14700 23851
rect 14648 23808 14700 23817
rect 18236 23851 18288 23860
rect 18236 23817 18245 23851
rect 18245 23817 18279 23851
rect 18279 23817 18288 23851
rect 18236 23808 18288 23817
rect 18604 23808 18656 23860
rect 8576 23715 8628 23724
rect 8576 23681 8610 23715
rect 8610 23681 8628 23715
rect 8576 23672 8628 23681
rect 10140 23672 10192 23724
rect 11980 23715 12032 23724
rect 7012 23604 7064 23656
rect 9588 23604 9640 23656
rect 11980 23681 11989 23715
rect 11989 23681 12023 23715
rect 12023 23681 12032 23715
rect 11980 23672 12032 23681
rect 15200 23740 15252 23792
rect 12900 23672 12952 23724
rect 13544 23672 13596 23724
rect 20628 23740 20680 23792
rect 21272 23740 21324 23792
rect 21732 23740 21784 23792
rect 22744 23783 22796 23792
rect 22744 23749 22753 23783
rect 22753 23749 22787 23783
rect 22787 23749 22796 23783
rect 22744 23740 22796 23749
rect 17960 23672 18012 23724
rect 21456 23672 21508 23724
rect 23112 23740 23164 23792
rect 24308 23783 24360 23792
rect 24308 23749 24317 23783
rect 24317 23749 24351 23783
rect 24351 23749 24360 23783
rect 24308 23740 24360 23749
rect 27988 23808 28040 23860
rect 32496 23851 32548 23860
rect 32496 23817 32505 23851
rect 32505 23817 32539 23851
rect 32539 23817 32548 23851
rect 32496 23808 32548 23817
rect 33140 23808 33192 23860
rect 39948 23808 40000 23860
rect 23020 23715 23072 23724
rect 23020 23681 23029 23715
rect 23029 23681 23063 23715
rect 23063 23681 23072 23715
rect 23020 23672 23072 23681
rect 25596 23715 25648 23724
rect 25596 23681 25605 23715
rect 25605 23681 25639 23715
rect 25639 23681 25648 23715
rect 25596 23672 25648 23681
rect 27620 23740 27672 23792
rect 28908 23740 28960 23792
rect 2596 23511 2648 23520
rect 2596 23477 2605 23511
rect 2605 23477 2639 23511
rect 2639 23477 2648 23511
rect 2596 23468 2648 23477
rect 10140 23468 10192 23520
rect 11888 23468 11940 23520
rect 17776 23536 17828 23588
rect 14648 23468 14700 23520
rect 22560 23536 22612 23588
rect 24676 23604 24728 23656
rect 23756 23536 23808 23588
rect 24124 23536 24176 23588
rect 24768 23536 24820 23588
rect 29644 23715 29696 23724
rect 30656 23740 30708 23792
rect 33508 23740 33560 23792
rect 34336 23740 34388 23792
rect 29644 23681 29662 23715
rect 29662 23681 29696 23715
rect 29644 23672 29696 23681
rect 35532 23672 35584 23724
rect 35992 23715 36044 23724
rect 35992 23681 36001 23715
rect 36001 23681 36035 23715
rect 36035 23681 36044 23715
rect 35992 23672 36044 23681
rect 36268 23672 36320 23724
rect 36912 23672 36964 23724
rect 33508 23647 33560 23656
rect 33508 23613 33517 23647
rect 33517 23613 33551 23647
rect 33551 23613 33560 23647
rect 33508 23604 33560 23613
rect 30012 23536 30064 23588
rect 33324 23536 33376 23588
rect 25872 23468 25924 23520
rect 33692 23511 33744 23520
rect 33692 23477 33701 23511
rect 33701 23477 33735 23511
rect 33735 23477 33744 23511
rect 33692 23468 33744 23477
rect 40868 23715 40920 23724
rect 40868 23681 40877 23715
rect 40877 23681 40911 23715
rect 40911 23681 40920 23715
rect 40868 23672 40920 23681
rect 40684 23604 40736 23656
rect 41144 23672 41196 23724
rect 41236 23715 41288 23724
rect 41236 23681 41245 23715
rect 41245 23681 41279 23715
rect 41279 23681 41288 23715
rect 41236 23672 41288 23681
rect 41052 23468 41104 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2964 23196 3016 23248
rect 3792 23128 3844 23180
rect 11336 23264 11388 23316
rect 11980 23264 12032 23316
rect 2688 23103 2740 23112
rect 2688 23069 2697 23103
rect 2697 23069 2731 23103
rect 2731 23069 2740 23103
rect 2688 23060 2740 23069
rect 7288 23103 7340 23112
rect 1584 22992 1636 23044
rect 7288 23069 7297 23103
rect 7297 23069 7331 23103
rect 7331 23069 7340 23103
rect 7288 23060 7340 23069
rect 11060 23060 11112 23112
rect 11612 23060 11664 23112
rect 12624 23060 12676 23112
rect 13820 23128 13872 23180
rect 14372 23128 14424 23180
rect 16304 23264 16356 23316
rect 16856 23307 16908 23316
rect 16856 23273 16865 23307
rect 16865 23273 16899 23307
rect 16899 23273 16908 23307
rect 16856 23264 16908 23273
rect 20260 23264 20312 23316
rect 14832 23103 14884 23112
rect 11704 22992 11756 23044
rect 14832 23069 14841 23103
rect 14841 23069 14875 23103
rect 14875 23069 14884 23103
rect 14832 23060 14884 23069
rect 14924 23060 14976 23112
rect 21364 23264 21416 23316
rect 22468 23264 22520 23316
rect 29644 23307 29696 23316
rect 29644 23273 29653 23307
rect 29653 23273 29687 23307
rect 29687 23273 29696 23307
rect 29644 23264 29696 23273
rect 29920 23264 29972 23316
rect 33876 23264 33928 23316
rect 39764 23264 39816 23316
rect 40868 23264 40920 23316
rect 16120 23060 16172 23112
rect 22560 23103 22612 23112
rect 15844 22992 15896 23044
rect 17960 22992 18012 23044
rect 20076 22992 20128 23044
rect 22560 23069 22569 23103
rect 22569 23069 22603 23103
rect 22603 23069 22612 23103
rect 22560 23060 22612 23069
rect 22652 22992 22704 23044
rect 25412 23128 25464 23180
rect 34060 23171 34112 23180
rect 34060 23137 34069 23171
rect 34069 23137 34103 23171
rect 34103 23137 34112 23171
rect 34060 23128 34112 23137
rect 35716 23128 35768 23180
rect 25872 23103 25924 23112
rect 25872 23069 25906 23103
rect 25906 23069 25924 23103
rect 25872 23060 25924 23069
rect 26240 23060 26292 23112
rect 34244 23060 34296 23112
rect 40776 23196 40828 23248
rect 2320 22967 2372 22976
rect 2320 22933 2329 22967
rect 2329 22933 2363 22967
rect 2363 22933 2372 22967
rect 2320 22924 2372 22933
rect 3792 22967 3844 22976
rect 3792 22933 3801 22967
rect 3801 22933 3835 22967
rect 3835 22933 3844 22967
rect 3792 22924 3844 22933
rect 9864 22924 9916 22976
rect 14740 22924 14792 22976
rect 15384 22967 15436 22976
rect 15384 22933 15393 22967
rect 15393 22933 15427 22967
rect 15427 22933 15436 22967
rect 15384 22924 15436 22933
rect 19340 22924 19392 22976
rect 22468 22924 22520 22976
rect 23756 22967 23808 22976
rect 23756 22933 23765 22967
rect 23765 22933 23799 22967
rect 23799 22933 23808 22967
rect 28816 22992 28868 23044
rect 31944 22992 31996 23044
rect 32036 23035 32088 23044
rect 32036 23001 32045 23035
rect 32045 23001 32079 23035
rect 32079 23001 32088 23035
rect 32036 22992 32088 23001
rect 23756 22924 23808 22933
rect 26332 22924 26384 22976
rect 27344 22924 27396 22976
rect 32220 22967 32272 22976
rect 32220 22933 32229 22967
rect 32229 22933 32263 22967
rect 32263 22933 32272 22967
rect 32220 22924 32272 22933
rect 33232 22992 33284 23044
rect 36176 23035 36228 23044
rect 36176 23001 36210 23035
rect 36210 23001 36228 23035
rect 40408 23103 40460 23112
rect 40408 23069 40417 23103
rect 40417 23069 40451 23103
rect 40451 23069 40460 23103
rect 40408 23060 40460 23069
rect 41144 23060 41196 23112
rect 36176 22992 36228 23001
rect 40684 22992 40736 23044
rect 36728 22924 36780 22976
rect 37280 22967 37332 22976
rect 37280 22933 37289 22967
rect 37289 22933 37323 22967
rect 37323 22933 37332 22967
rect 37280 22924 37332 22933
rect 40408 22924 40460 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 1584 22763 1636 22772
rect 1584 22729 1593 22763
rect 1593 22729 1627 22763
rect 1627 22729 1636 22763
rect 1584 22720 1636 22729
rect 2320 22652 2372 22704
rect 5172 22652 5224 22704
rect 6000 22720 6052 22772
rect 10416 22720 10468 22772
rect 2412 22627 2464 22636
rect 2412 22593 2421 22627
rect 2421 22593 2455 22627
rect 2455 22593 2464 22627
rect 2412 22584 2464 22593
rect 2228 22516 2280 22568
rect 6368 22584 6420 22636
rect 6920 22627 6972 22636
rect 6920 22593 6954 22627
rect 6954 22593 6972 22627
rect 6920 22584 6972 22593
rect 11980 22652 12032 22704
rect 8668 22627 8720 22636
rect 8668 22593 8677 22627
rect 8677 22593 8711 22627
rect 8711 22593 8720 22627
rect 8668 22584 8720 22593
rect 9220 22584 9272 22636
rect 10324 22584 10376 22636
rect 8116 22516 8168 22568
rect 11704 22627 11756 22636
rect 11704 22593 11713 22627
rect 11713 22593 11747 22627
rect 11747 22593 11756 22627
rect 11704 22584 11756 22593
rect 11888 22627 11940 22636
rect 11888 22593 11897 22627
rect 11897 22593 11931 22627
rect 11931 22593 11940 22627
rect 11888 22584 11940 22593
rect 11060 22516 11112 22568
rect 16120 22763 16172 22772
rect 16120 22729 16129 22763
rect 16129 22729 16163 22763
rect 16163 22729 16172 22763
rect 16120 22720 16172 22729
rect 14188 22652 14240 22704
rect 14924 22652 14976 22704
rect 18604 22720 18656 22772
rect 18788 22720 18840 22772
rect 20168 22720 20220 22772
rect 23756 22720 23808 22772
rect 24952 22720 25004 22772
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 16488 22584 16540 22636
rect 18788 22584 18840 22636
rect 23940 22652 23992 22704
rect 20904 22627 20956 22636
rect 20904 22593 20913 22627
rect 20913 22593 20947 22627
rect 20947 22593 20956 22627
rect 20904 22584 20956 22593
rect 22192 22627 22244 22636
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 24124 22627 24176 22636
rect 24124 22593 24133 22627
rect 24133 22593 24167 22627
rect 24167 22593 24176 22627
rect 24124 22584 24176 22593
rect 24768 22584 24820 22636
rect 25596 22720 25648 22772
rect 25872 22652 25924 22704
rect 27804 22720 27856 22772
rect 27344 22652 27396 22704
rect 33048 22720 33100 22772
rect 33232 22763 33284 22772
rect 33232 22729 33241 22763
rect 33241 22729 33275 22763
rect 33275 22729 33284 22763
rect 33232 22720 33284 22729
rect 33692 22763 33744 22772
rect 33692 22729 33701 22763
rect 33701 22729 33735 22763
rect 33735 22729 33744 22763
rect 33692 22720 33744 22729
rect 36176 22720 36228 22772
rect 32128 22652 32180 22704
rect 32220 22652 32272 22704
rect 34060 22695 34112 22704
rect 16672 22559 16724 22568
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 4620 22380 4672 22432
rect 6368 22380 6420 22432
rect 14832 22448 14884 22500
rect 16304 22448 16356 22500
rect 20076 22491 20128 22500
rect 20076 22457 20085 22491
rect 20085 22457 20119 22491
rect 20119 22457 20128 22491
rect 20076 22448 20128 22457
rect 20628 22448 20680 22500
rect 21364 22448 21416 22500
rect 23572 22516 23624 22568
rect 24676 22516 24728 22568
rect 28172 22584 28224 22636
rect 28908 22516 28960 22568
rect 8392 22380 8444 22432
rect 10324 22423 10376 22432
rect 10324 22389 10333 22423
rect 10333 22389 10367 22423
rect 10367 22389 10376 22423
rect 10324 22380 10376 22389
rect 12900 22380 12952 22432
rect 14464 22380 14516 22432
rect 14740 22380 14792 22432
rect 21088 22380 21140 22432
rect 21640 22380 21692 22432
rect 23664 22448 23716 22500
rect 31392 22627 31444 22636
rect 31392 22593 31401 22627
rect 31401 22593 31435 22627
rect 31435 22593 31444 22627
rect 31392 22584 31444 22593
rect 32312 22584 32364 22636
rect 32864 22627 32916 22636
rect 32864 22593 32873 22627
rect 32873 22593 32907 22627
rect 32907 22593 32916 22627
rect 32864 22584 32916 22593
rect 33140 22584 33192 22636
rect 34060 22661 34069 22695
rect 34069 22661 34103 22695
rect 34103 22661 34112 22695
rect 34060 22652 34112 22661
rect 37280 22652 37332 22704
rect 38568 22652 38620 22704
rect 33968 22627 34020 22636
rect 33968 22593 33977 22627
rect 33977 22593 34011 22627
rect 34011 22593 34020 22627
rect 34244 22627 34296 22636
rect 33968 22584 34020 22593
rect 34244 22593 34253 22627
rect 34253 22593 34287 22627
rect 34287 22593 34296 22627
rect 34244 22584 34296 22593
rect 33784 22448 33836 22500
rect 22560 22380 22612 22432
rect 28080 22380 28132 22432
rect 32956 22380 33008 22432
rect 33140 22380 33192 22432
rect 35624 22627 35676 22636
rect 35624 22593 35633 22627
rect 35633 22593 35667 22627
rect 35667 22593 35676 22627
rect 35624 22584 35676 22593
rect 36360 22627 36412 22636
rect 36360 22593 36369 22627
rect 36369 22593 36403 22627
rect 36403 22593 36412 22627
rect 36360 22584 36412 22593
rect 36728 22627 36780 22636
rect 36268 22448 36320 22500
rect 36728 22593 36737 22627
rect 36737 22593 36771 22627
rect 36771 22593 36780 22627
rect 36728 22584 36780 22593
rect 37004 22584 37056 22636
rect 38476 22584 38528 22636
rect 38936 22584 38988 22636
rect 39764 22516 39816 22568
rect 40408 22448 40460 22500
rect 58164 22491 58216 22500
rect 58164 22457 58173 22491
rect 58173 22457 58207 22491
rect 58207 22457 58216 22491
rect 58164 22448 58216 22457
rect 35992 22380 36044 22432
rect 40316 22380 40368 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3240 22219 3292 22228
rect 3240 22185 3249 22219
rect 3249 22185 3283 22219
rect 3283 22185 3292 22219
rect 3240 22176 3292 22185
rect 8116 22176 8168 22228
rect 8668 22176 8720 22228
rect 14924 22219 14976 22228
rect 6092 22040 6144 22092
rect 2872 21972 2924 22024
rect 6368 22015 6420 22024
rect 2136 21947 2188 21956
rect 2136 21913 2170 21947
rect 2170 21913 2188 21947
rect 2136 21904 2188 21913
rect 3700 21904 3752 21956
rect 4160 21904 4212 21956
rect 5080 21904 5132 21956
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 6552 22015 6604 22024
rect 6552 21981 6561 22015
rect 6561 21981 6595 22015
rect 6595 21981 6604 22015
rect 6920 22040 6972 22092
rect 14924 22185 14933 22219
rect 14933 22185 14967 22219
rect 14967 22185 14976 22219
rect 14924 22176 14976 22185
rect 15200 22176 15252 22228
rect 16580 22176 16632 22228
rect 17684 22176 17736 22228
rect 18788 22176 18840 22228
rect 10324 22108 10376 22160
rect 12808 22108 12860 22160
rect 6552 21972 6604 21981
rect 7012 21972 7064 22024
rect 7288 22015 7340 22024
rect 7288 21981 7297 22015
rect 7297 21981 7331 22015
rect 7331 21981 7340 22015
rect 7288 21972 7340 21981
rect 7472 22015 7524 22024
rect 7472 21981 7481 22015
rect 7481 21981 7515 22015
rect 7515 21981 7524 22015
rect 7472 21972 7524 21981
rect 6920 21904 6972 21956
rect 8392 21972 8444 22024
rect 9956 21972 10008 22024
rect 11060 21972 11112 22024
rect 5172 21879 5224 21888
rect 5172 21845 5181 21879
rect 5181 21845 5215 21879
rect 5215 21845 5224 21879
rect 5172 21836 5224 21845
rect 6736 21836 6788 21888
rect 8300 21904 8352 21956
rect 10048 21947 10100 21956
rect 10048 21913 10057 21947
rect 10057 21913 10091 21947
rect 10091 21913 10100 21947
rect 15844 22040 15896 22092
rect 15200 21972 15252 22024
rect 17592 22108 17644 22160
rect 20812 22176 20864 22228
rect 20996 22176 21048 22228
rect 22008 22176 22060 22228
rect 24308 22176 24360 22228
rect 28908 22176 28960 22228
rect 16120 21972 16172 22024
rect 16304 22015 16356 22024
rect 16304 21981 16313 22015
rect 16313 21981 16347 22015
rect 16347 21981 16356 22015
rect 16304 21972 16356 21981
rect 17132 22040 17184 22092
rect 16948 21972 17000 22024
rect 17224 22015 17276 22024
rect 17224 21981 17233 22015
rect 17233 21981 17267 22015
rect 17267 21981 17276 22015
rect 17224 21972 17276 21981
rect 17500 21972 17552 22024
rect 18052 22015 18104 22024
rect 18052 21981 18061 22015
rect 18061 21981 18095 22015
rect 18095 21981 18104 22015
rect 18052 21972 18104 21981
rect 19340 22040 19392 22092
rect 22652 22108 22704 22160
rect 10048 21904 10100 21913
rect 7932 21879 7984 21888
rect 7932 21845 7941 21879
rect 7941 21845 7975 21879
rect 7975 21845 7984 21879
rect 7932 21836 7984 21845
rect 10600 21836 10652 21888
rect 11704 21836 11756 21888
rect 15660 21879 15712 21888
rect 15660 21845 15669 21879
rect 15669 21845 15703 21879
rect 15703 21845 15712 21879
rect 16948 21879 17000 21888
rect 15660 21836 15712 21845
rect 16948 21845 16957 21879
rect 16957 21845 16991 21879
rect 16991 21845 17000 21879
rect 16948 21836 17000 21845
rect 18604 21972 18656 22024
rect 20812 22040 20864 22092
rect 22376 22040 22428 22092
rect 21916 21972 21968 22024
rect 22560 21972 22612 22024
rect 23572 22040 23624 22092
rect 25964 22040 26016 22092
rect 23480 22015 23532 22024
rect 23480 21981 23489 22015
rect 23489 21981 23523 22015
rect 23523 21981 23532 22015
rect 23480 21972 23532 21981
rect 20720 21904 20772 21956
rect 18420 21836 18472 21888
rect 19064 21836 19116 21888
rect 20260 21879 20312 21888
rect 20260 21845 20269 21879
rect 20269 21845 20303 21879
rect 20303 21845 20312 21879
rect 22100 21904 22152 21956
rect 24308 21972 24360 22024
rect 26608 21972 26660 22024
rect 29920 22040 29972 22092
rect 31392 22040 31444 22092
rect 29276 21972 29328 22024
rect 32036 21972 32088 22024
rect 33048 21972 33100 22024
rect 33324 22040 33376 22092
rect 33416 22015 33468 22024
rect 23020 21879 23072 21888
rect 20260 21836 20312 21845
rect 23020 21845 23029 21879
rect 23029 21845 23063 21879
rect 23063 21845 23072 21879
rect 23020 21836 23072 21845
rect 23664 21836 23716 21888
rect 26884 21879 26936 21888
rect 26884 21845 26893 21879
rect 26893 21845 26927 21879
rect 26927 21845 26936 21879
rect 26884 21836 26936 21845
rect 27712 21904 27764 21956
rect 32128 21947 32180 21956
rect 32128 21913 32137 21947
rect 32137 21913 32171 21947
rect 32171 21913 32180 21947
rect 32128 21904 32180 21913
rect 33416 21981 33425 22015
rect 33425 21981 33459 22015
rect 33459 21981 33468 22015
rect 33416 21972 33468 21981
rect 35992 22015 36044 22024
rect 35992 21981 36001 22015
rect 36001 21981 36035 22015
rect 36035 21981 36044 22015
rect 35992 21972 36044 21981
rect 36084 22015 36136 22024
rect 36084 21981 36093 22015
rect 36093 21981 36127 22015
rect 36127 21981 36136 22015
rect 36084 21972 36136 21981
rect 37188 21972 37240 22024
rect 40040 21972 40092 22024
rect 33692 21904 33744 21956
rect 36268 21904 36320 21956
rect 40316 22015 40368 22021
rect 40316 21981 40325 22015
rect 40325 21981 40359 22015
rect 40359 21981 40368 22015
rect 40500 22015 40552 22024
rect 40316 21969 40368 21981
rect 40500 21981 40509 22015
rect 40509 21981 40543 22015
rect 40543 21981 40552 22015
rect 40500 21972 40552 21981
rect 35532 21836 35584 21888
rect 39856 21879 39908 21888
rect 39856 21845 39865 21879
rect 39865 21845 39899 21879
rect 39899 21845 39908 21879
rect 39856 21836 39908 21845
rect 40224 21836 40276 21888
rect 40960 21836 41012 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 2136 21632 2188 21684
rect 3700 21675 3752 21684
rect 3700 21641 3709 21675
rect 3709 21641 3743 21675
rect 3743 21641 3752 21675
rect 3700 21632 3752 21641
rect 2780 21564 2832 21616
rect 6092 21632 6144 21684
rect 6184 21632 6236 21684
rect 14648 21632 14700 21684
rect 15936 21632 15988 21684
rect 16304 21632 16356 21684
rect 18052 21632 18104 21684
rect 2596 21496 2648 21548
rect 3976 21539 4028 21548
rect 3976 21505 3985 21539
rect 3985 21505 4019 21539
rect 4019 21505 4028 21539
rect 3976 21496 4028 21505
rect 4620 21564 4672 21616
rect 5080 21564 5132 21616
rect 5172 21564 5224 21616
rect 6920 21496 6972 21548
rect 7932 21564 7984 21616
rect 8300 21607 8352 21616
rect 8300 21573 8309 21607
rect 8309 21573 8343 21607
rect 8343 21573 8352 21607
rect 8300 21564 8352 21573
rect 10140 21607 10192 21616
rect 10140 21573 10149 21607
rect 10149 21573 10183 21607
rect 10183 21573 10192 21607
rect 10140 21564 10192 21573
rect 16396 21564 16448 21616
rect 16948 21607 17000 21616
rect 16948 21573 16982 21607
rect 16982 21573 17000 21607
rect 16948 21564 17000 21573
rect 20720 21632 20772 21684
rect 25964 21632 26016 21684
rect 27712 21632 27764 21684
rect 28816 21632 28868 21684
rect 29644 21632 29696 21684
rect 32036 21632 32088 21684
rect 21824 21564 21876 21616
rect 23020 21564 23072 21616
rect 23940 21564 23992 21616
rect 10048 21539 10100 21548
rect 10048 21505 10057 21539
rect 10057 21505 10091 21539
rect 10091 21505 10100 21539
rect 10048 21496 10100 21505
rect 11060 21496 11112 21548
rect 15384 21539 15436 21548
rect 15384 21505 15393 21539
rect 15393 21505 15427 21539
rect 15427 21505 15436 21539
rect 15384 21496 15436 21505
rect 8300 21428 8352 21480
rect 14004 21428 14056 21480
rect 16304 21496 16356 21548
rect 16488 21496 16540 21548
rect 17224 21496 17276 21548
rect 20444 21496 20496 21548
rect 21548 21496 21600 21548
rect 26700 21496 26752 21548
rect 8116 21360 8168 21412
rect 12440 21360 12492 21412
rect 13636 21360 13688 21412
rect 2504 21292 2556 21344
rect 3240 21335 3292 21344
rect 3240 21301 3249 21335
rect 3249 21301 3283 21335
rect 3283 21301 3292 21335
rect 3240 21292 3292 21301
rect 11428 21292 11480 21344
rect 14280 21335 14332 21344
rect 14280 21301 14289 21335
rect 14289 21301 14323 21335
rect 14323 21301 14332 21335
rect 14280 21292 14332 21301
rect 20444 21403 20496 21412
rect 20444 21369 20453 21403
rect 20453 21369 20487 21403
rect 20487 21369 20496 21403
rect 20444 21360 20496 21369
rect 22560 21360 22612 21412
rect 16948 21292 17000 21344
rect 17592 21292 17644 21344
rect 18052 21335 18104 21344
rect 18052 21301 18061 21335
rect 18061 21301 18095 21335
rect 18095 21301 18104 21335
rect 18052 21292 18104 21301
rect 22192 21335 22244 21344
rect 22192 21301 22201 21335
rect 22201 21301 22235 21335
rect 22235 21301 22244 21335
rect 22192 21292 22244 21301
rect 23204 21292 23256 21344
rect 26608 21428 26660 21480
rect 27436 21428 27488 21480
rect 28080 21539 28132 21548
rect 28080 21505 28089 21539
rect 28089 21505 28123 21539
rect 28123 21505 28132 21539
rect 28264 21539 28316 21548
rect 28080 21496 28132 21505
rect 28264 21505 28273 21539
rect 28273 21505 28307 21539
rect 28307 21505 28316 21539
rect 28264 21496 28316 21505
rect 28448 21496 28500 21548
rect 34612 21632 34664 21684
rect 33600 21564 33652 21616
rect 39856 21564 39908 21616
rect 29000 21428 29052 21480
rect 29644 21428 29696 21480
rect 33140 21496 33192 21548
rect 29828 21471 29880 21480
rect 29828 21437 29837 21471
rect 29837 21437 29871 21471
rect 29871 21437 29880 21471
rect 29828 21428 29880 21437
rect 31852 21428 31904 21480
rect 39948 21471 40000 21480
rect 39948 21437 39957 21471
rect 39957 21437 39991 21471
rect 39991 21437 40000 21471
rect 39948 21428 40000 21437
rect 37280 21360 37332 21412
rect 27252 21292 27304 21344
rect 29736 21335 29788 21344
rect 29736 21301 29745 21335
rect 29745 21301 29779 21335
rect 29779 21301 29788 21335
rect 29736 21292 29788 21301
rect 32956 21335 33008 21344
rect 32956 21301 32965 21335
rect 32965 21301 32999 21335
rect 32999 21301 33008 21335
rect 32956 21292 33008 21301
rect 35900 21335 35952 21344
rect 35900 21301 35909 21335
rect 35909 21301 35943 21335
rect 35943 21301 35952 21335
rect 35900 21292 35952 21301
rect 36360 21292 36412 21344
rect 37832 21292 37884 21344
rect 38568 21335 38620 21344
rect 38568 21301 38577 21335
rect 38577 21301 38611 21335
rect 38611 21301 38620 21335
rect 38568 21292 38620 21301
rect 58164 21335 58216 21344
rect 58164 21301 58173 21335
rect 58173 21301 58207 21335
rect 58207 21301 58216 21335
rect 58164 21292 58216 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 7472 21088 7524 21140
rect 10692 21088 10744 21140
rect 16488 21088 16540 21140
rect 17500 21088 17552 21140
rect 23480 21088 23532 21140
rect 26332 21088 26384 21140
rect 26700 21088 26752 21140
rect 32036 21088 32088 21140
rect 35900 21088 35952 21140
rect 6644 21020 6696 21072
rect 8116 21063 8168 21072
rect 8116 21029 8125 21063
rect 8125 21029 8159 21063
rect 8159 21029 8168 21063
rect 8116 21020 8168 21029
rect 11612 21063 11664 21072
rect 11612 21029 11621 21063
rect 11621 21029 11655 21063
rect 11655 21029 11664 21063
rect 11612 21020 11664 21029
rect 13912 21020 13964 21072
rect 16304 21020 16356 21072
rect 21456 21020 21508 21072
rect 6000 20927 6052 20936
rect 6000 20893 6009 20927
rect 6009 20893 6043 20927
rect 6043 20893 6052 20927
rect 6000 20884 6052 20893
rect 6184 20927 6236 20936
rect 6184 20893 6193 20927
rect 6193 20893 6227 20927
rect 6227 20893 6236 20927
rect 6184 20884 6236 20893
rect 13452 20952 13504 21004
rect 18144 20952 18196 21004
rect 13360 20884 13412 20936
rect 13912 20884 13964 20936
rect 14280 20884 14332 20936
rect 17592 20884 17644 20936
rect 18052 20884 18104 20936
rect 19340 20884 19392 20936
rect 8392 20816 8444 20868
rect 10968 20816 11020 20868
rect 14004 20816 14056 20868
rect 16028 20816 16080 20868
rect 17960 20859 18012 20868
rect 17960 20825 17969 20859
rect 17969 20825 18003 20859
rect 18003 20825 18012 20859
rect 17960 20816 18012 20825
rect 20168 20816 20220 20868
rect 21272 20816 21324 20868
rect 24768 21020 24820 21072
rect 22100 20952 22152 21004
rect 22192 20816 22244 20868
rect 23112 20927 23164 20936
rect 23112 20893 23121 20927
rect 23121 20893 23155 20927
rect 23155 20893 23164 20927
rect 23112 20884 23164 20893
rect 23572 20884 23624 20936
rect 27160 20952 27212 21004
rect 29184 20952 29236 21004
rect 26608 20927 26660 20936
rect 26608 20893 26617 20927
rect 26617 20893 26651 20927
rect 26651 20893 26660 20927
rect 26608 20884 26660 20893
rect 27252 20884 27304 20936
rect 23480 20816 23532 20868
rect 24584 20859 24636 20868
rect 24584 20825 24593 20859
rect 24593 20825 24627 20859
rect 24627 20825 24636 20859
rect 24584 20816 24636 20825
rect 26976 20816 27028 20868
rect 13268 20748 13320 20800
rect 16948 20748 17000 20800
rect 21732 20748 21784 20800
rect 22836 20748 22888 20800
rect 23388 20791 23440 20800
rect 23388 20757 23397 20791
rect 23397 20757 23431 20791
rect 23431 20757 23440 20791
rect 23388 20748 23440 20757
rect 25228 20791 25280 20800
rect 25228 20757 25237 20791
rect 25237 20757 25271 20791
rect 25271 20757 25280 20791
rect 25228 20748 25280 20757
rect 26240 20748 26292 20800
rect 26884 20748 26936 20800
rect 29184 20816 29236 20868
rect 27252 20748 27304 20800
rect 28448 20791 28500 20800
rect 28448 20757 28457 20791
rect 28457 20757 28491 20791
rect 28491 20757 28500 20791
rect 28448 20748 28500 20757
rect 29000 20748 29052 20800
rect 29828 20748 29880 20800
rect 30104 20791 30156 20800
rect 30104 20757 30113 20791
rect 30113 20757 30147 20791
rect 30147 20757 30156 20791
rect 30104 20748 30156 20757
rect 30380 20748 30432 20800
rect 32220 20791 32272 20800
rect 32220 20757 32229 20791
rect 32229 20757 32263 20791
rect 32263 20757 32272 20791
rect 32220 20748 32272 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 3056 20476 3108 20528
rect 11244 20544 11296 20596
rect 11612 20544 11664 20596
rect 11888 20544 11940 20596
rect 14004 20587 14056 20596
rect 14004 20553 14013 20587
rect 14013 20553 14047 20587
rect 14047 20553 14056 20587
rect 14004 20544 14056 20553
rect 16028 20587 16080 20596
rect 16028 20553 16037 20587
rect 16037 20553 16071 20587
rect 16071 20553 16080 20587
rect 16028 20544 16080 20553
rect 16948 20587 17000 20596
rect 16948 20553 16957 20587
rect 16957 20553 16991 20587
rect 16991 20553 17000 20587
rect 16948 20544 17000 20553
rect 4804 20451 4856 20460
rect 4804 20417 4813 20451
rect 4813 20417 4847 20451
rect 4847 20417 4856 20451
rect 16488 20476 16540 20528
rect 4804 20408 4856 20417
rect 12716 20408 12768 20460
rect 13360 20408 13412 20460
rect 15752 20408 15804 20460
rect 18788 20476 18840 20528
rect 19248 20451 19300 20460
rect 19248 20417 19260 20451
rect 19260 20417 19294 20451
rect 19294 20417 19300 20451
rect 19248 20408 19300 20417
rect 19432 20451 19484 20460
rect 20812 20476 20864 20528
rect 22652 20587 22704 20596
rect 22652 20553 22661 20587
rect 22661 20553 22695 20587
rect 22695 20553 22704 20587
rect 22652 20544 22704 20553
rect 23112 20544 23164 20596
rect 26976 20587 27028 20596
rect 25228 20476 25280 20528
rect 26976 20553 26985 20587
rect 26985 20553 27019 20587
rect 27019 20553 27028 20587
rect 26976 20544 27028 20553
rect 29736 20587 29788 20596
rect 29736 20553 29745 20587
rect 29745 20553 29779 20587
rect 29779 20553 29788 20587
rect 29736 20544 29788 20553
rect 19432 20417 19477 20451
rect 19477 20417 19484 20451
rect 19432 20408 19484 20417
rect 15568 20272 15620 20324
rect 17960 20272 18012 20324
rect 20168 20340 20220 20392
rect 20444 20451 20496 20460
rect 20444 20417 20453 20451
rect 20453 20417 20487 20451
rect 20487 20417 20496 20451
rect 20628 20451 20680 20460
rect 20444 20408 20496 20417
rect 20628 20417 20636 20451
rect 20636 20417 20670 20451
rect 20670 20417 20680 20451
rect 20628 20408 20680 20417
rect 20904 20408 20956 20460
rect 22100 20451 22152 20460
rect 22100 20417 22109 20451
rect 22109 20417 22143 20451
rect 22143 20417 22152 20451
rect 22100 20408 22152 20417
rect 23112 20451 23164 20460
rect 23112 20417 23121 20451
rect 23121 20417 23155 20451
rect 23155 20417 23164 20451
rect 23112 20408 23164 20417
rect 23388 20451 23440 20460
rect 23388 20417 23422 20451
rect 23422 20417 23440 20451
rect 23388 20408 23440 20417
rect 23848 20408 23900 20460
rect 25872 20451 25924 20460
rect 25872 20417 25881 20451
rect 25881 20417 25915 20451
rect 25915 20417 25924 20451
rect 25872 20408 25924 20417
rect 27068 20408 27120 20460
rect 27252 20451 27304 20460
rect 27252 20417 27261 20451
rect 27261 20417 27295 20451
rect 27295 20417 27304 20451
rect 27252 20408 27304 20417
rect 21916 20340 21968 20392
rect 20444 20272 20496 20324
rect 26884 20272 26936 20324
rect 27436 20272 27488 20324
rect 7932 20204 7984 20256
rect 8392 20204 8444 20256
rect 17592 20247 17644 20256
rect 17592 20213 17601 20247
rect 17601 20213 17635 20247
rect 17635 20213 17644 20247
rect 17592 20204 17644 20213
rect 17868 20247 17920 20256
rect 17868 20213 17877 20247
rect 17877 20213 17911 20247
rect 17911 20213 17920 20247
rect 17868 20204 17920 20213
rect 18788 20204 18840 20256
rect 19892 20204 19944 20256
rect 20076 20247 20128 20256
rect 20076 20213 20085 20247
rect 20085 20213 20119 20247
rect 20119 20213 20128 20247
rect 20076 20204 20128 20213
rect 24584 20204 24636 20256
rect 27896 20408 27948 20460
rect 28632 20408 28684 20460
rect 29368 20451 29420 20460
rect 29368 20417 29377 20451
rect 29377 20417 29411 20451
rect 29411 20417 29420 20451
rect 29368 20408 29420 20417
rect 29552 20451 29604 20460
rect 29552 20417 29561 20451
rect 29561 20417 29595 20451
rect 29595 20417 29604 20451
rect 36912 20544 36964 20596
rect 37280 20587 37332 20596
rect 37280 20553 37289 20587
rect 37289 20553 37323 20587
rect 37323 20553 37332 20587
rect 37280 20544 37332 20553
rect 30656 20519 30708 20528
rect 30656 20485 30665 20519
rect 30665 20485 30699 20519
rect 30699 20485 30708 20519
rect 30656 20476 30708 20485
rect 29552 20408 29604 20417
rect 32312 20408 32364 20460
rect 30472 20383 30524 20392
rect 30472 20349 30481 20383
rect 30481 20349 30515 20383
rect 30515 20349 30524 20383
rect 30472 20340 30524 20349
rect 32680 20451 32732 20460
rect 32680 20417 32689 20451
rect 32689 20417 32723 20451
rect 32723 20417 32732 20451
rect 32680 20408 32732 20417
rect 32864 20408 32916 20460
rect 27896 20204 27948 20256
rect 28264 20204 28316 20256
rect 30380 20247 30432 20256
rect 30380 20213 30389 20247
rect 30389 20213 30423 20247
rect 30423 20213 30432 20247
rect 30380 20204 30432 20213
rect 33048 20272 33100 20324
rect 32864 20204 32916 20256
rect 34244 20204 34296 20256
rect 36268 20408 36320 20460
rect 37188 20408 37240 20460
rect 37832 20451 37884 20460
rect 37096 20340 37148 20392
rect 37832 20417 37841 20451
rect 37841 20417 37875 20451
rect 37875 20417 37884 20451
rect 37832 20408 37884 20417
rect 39580 20408 39632 20460
rect 39764 20408 39816 20460
rect 39948 20340 40000 20392
rect 40684 20204 40736 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7196 20000 7248 20052
rect 12716 20043 12768 20052
rect 12716 20009 12725 20043
rect 12725 20009 12759 20043
rect 12759 20009 12768 20043
rect 12716 20000 12768 20009
rect 15568 20043 15620 20052
rect 15568 20009 15577 20043
rect 15577 20009 15611 20043
rect 15611 20009 15620 20043
rect 15568 20000 15620 20009
rect 22100 20000 22152 20052
rect 23572 20000 23624 20052
rect 33048 20043 33100 20052
rect 33048 20009 33057 20043
rect 33057 20009 33091 20043
rect 33091 20009 33100 20043
rect 33048 20000 33100 20009
rect 36912 20000 36964 20052
rect 39580 20000 39632 20052
rect 3240 19932 3292 19984
rect 9404 19932 9456 19984
rect 18052 19932 18104 19984
rect 26332 19932 26384 19984
rect 27160 19932 27212 19984
rect 36728 19932 36780 19984
rect 2596 19839 2648 19848
rect 2596 19805 2605 19839
rect 2605 19805 2639 19839
rect 2639 19805 2648 19839
rect 2596 19796 2648 19805
rect 4804 19796 4856 19848
rect 8300 19796 8352 19848
rect 11336 19796 11388 19848
rect 12440 19864 12492 19916
rect 11704 19839 11756 19848
rect 11704 19805 11713 19839
rect 11713 19805 11747 19839
rect 11747 19805 11756 19839
rect 11704 19796 11756 19805
rect 11888 19839 11940 19848
rect 11888 19805 11897 19839
rect 11897 19805 11931 19839
rect 11931 19805 11940 19839
rect 11888 19796 11940 19805
rect 12164 19796 12216 19848
rect 12716 19796 12768 19848
rect 13268 19796 13320 19848
rect 13452 19796 13504 19848
rect 14188 19796 14240 19848
rect 16120 19864 16172 19916
rect 15752 19839 15804 19848
rect 15752 19805 15761 19839
rect 15761 19805 15795 19839
rect 15795 19805 15804 19839
rect 15752 19796 15804 19805
rect 15844 19839 15896 19848
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 20352 19864 20404 19916
rect 15844 19796 15896 19805
rect 6000 19728 6052 19780
rect 19340 19728 19392 19780
rect 19892 19796 19944 19848
rect 20168 19839 20220 19848
rect 20168 19805 20182 19839
rect 20182 19805 20216 19839
rect 20216 19805 20220 19839
rect 20168 19796 20220 19805
rect 21180 19796 21232 19848
rect 29920 19907 29972 19916
rect 29920 19873 29929 19907
rect 29929 19873 29963 19907
rect 29963 19873 29972 19907
rect 29920 19864 29972 19873
rect 30840 19864 30892 19916
rect 31392 19864 31444 19916
rect 35992 19864 36044 19916
rect 40408 19864 40460 19916
rect 20720 19728 20772 19780
rect 22192 19796 22244 19848
rect 24400 19796 24452 19848
rect 25688 19796 25740 19848
rect 28816 19796 28868 19848
rect 29552 19796 29604 19848
rect 31944 19796 31996 19848
rect 32864 19839 32916 19848
rect 32864 19805 32873 19839
rect 32873 19805 32907 19839
rect 32907 19805 32916 19839
rect 32864 19796 32916 19805
rect 37188 19796 37240 19848
rect 22376 19728 22428 19780
rect 27436 19771 27488 19780
rect 27436 19737 27445 19771
rect 27445 19737 27479 19771
rect 27479 19737 27488 19771
rect 27436 19728 27488 19737
rect 37096 19728 37148 19780
rect 38752 19796 38804 19848
rect 40040 19796 40092 19848
rect 40776 19864 40828 19916
rect 40684 19839 40736 19848
rect 40684 19805 40693 19839
rect 40693 19805 40727 19839
rect 40727 19805 40736 19839
rect 40684 19796 40736 19805
rect 41144 19796 41196 19848
rect 58164 19839 58216 19848
rect 58164 19805 58173 19839
rect 58173 19805 58207 19839
rect 58207 19805 58216 19839
rect 58164 19796 58216 19805
rect 41696 19728 41748 19780
rect 2412 19703 2464 19712
rect 2412 19669 2421 19703
rect 2421 19669 2455 19703
rect 2455 19669 2464 19703
rect 2412 19660 2464 19669
rect 5632 19703 5684 19712
rect 5632 19669 5641 19703
rect 5641 19669 5675 19703
rect 5675 19669 5684 19703
rect 5632 19660 5684 19669
rect 5908 19660 5960 19712
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 8392 19660 8444 19669
rect 10508 19660 10560 19712
rect 11336 19660 11388 19712
rect 13912 19660 13964 19712
rect 20352 19703 20404 19712
rect 20352 19669 20361 19703
rect 20361 19669 20395 19703
rect 20395 19669 20404 19703
rect 20352 19660 20404 19669
rect 26608 19660 26660 19712
rect 27252 19660 27304 19712
rect 27896 19703 27948 19712
rect 27896 19669 27905 19703
rect 27905 19669 27939 19703
rect 27939 19669 27948 19703
rect 27896 19660 27948 19669
rect 32220 19660 32272 19712
rect 40040 19660 40092 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 5632 19456 5684 19508
rect 5908 19388 5960 19440
rect 7564 19456 7616 19508
rect 7932 19388 7984 19440
rect 4620 19320 4672 19372
rect 5264 19363 5316 19372
rect 5264 19329 5273 19363
rect 5273 19329 5307 19363
rect 5307 19329 5316 19363
rect 5264 19320 5316 19329
rect 8576 19388 8628 19440
rect 4896 19252 4948 19304
rect 11336 19456 11388 19508
rect 11704 19456 11756 19508
rect 14188 19499 14240 19508
rect 14188 19465 14197 19499
rect 14197 19465 14231 19499
rect 14231 19465 14240 19499
rect 14188 19456 14240 19465
rect 14372 19456 14424 19508
rect 14924 19456 14976 19508
rect 13636 19388 13688 19440
rect 21180 19456 21232 19508
rect 26884 19456 26936 19508
rect 10508 19320 10560 19372
rect 12532 19320 12584 19372
rect 13360 19320 13412 19372
rect 14280 19320 14332 19372
rect 20076 19388 20128 19440
rect 21916 19388 21968 19440
rect 30380 19456 30432 19508
rect 16488 19320 16540 19372
rect 16764 19320 16816 19372
rect 22192 19363 22244 19372
rect 8116 19295 8168 19304
rect 8116 19261 8125 19295
rect 8125 19261 8159 19295
rect 8159 19261 8168 19295
rect 8116 19252 8168 19261
rect 8392 19252 8444 19304
rect 2872 19227 2924 19236
rect 2872 19193 2881 19227
rect 2881 19193 2915 19227
rect 2915 19193 2924 19227
rect 2872 19184 2924 19193
rect 7656 19184 7708 19236
rect 4804 19159 4856 19168
rect 4804 19125 4813 19159
rect 4813 19125 4847 19159
rect 4847 19125 4856 19159
rect 4804 19116 4856 19125
rect 7472 19116 7524 19168
rect 11704 19184 11756 19236
rect 21456 19252 21508 19304
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 27528 19388 27580 19440
rect 32404 19388 32456 19440
rect 33784 19456 33836 19508
rect 36268 19456 36320 19508
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 27344 19320 27396 19372
rect 24676 19252 24728 19304
rect 26700 19252 26752 19304
rect 28356 19252 28408 19304
rect 28816 19363 28868 19372
rect 28816 19329 28825 19363
rect 28825 19329 28859 19363
rect 28859 19329 28868 19363
rect 28816 19320 28868 19329
rect 29368 19252 29420 19304
rect 30840 19320 30892 19372
rect 29736 19295 29788 19304
rect 29736 19261 29745 19295
rect 29745 19261 29779 19295
rect 29779 19261 29788 19295
rect 29736 19252 29788 19261
rect 30748 19252 30800 19304
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 8852 19116 8904 19125
rect 11244 19116 11296 19168
rect 12716 19116 12768 19168
rect 15016 19159 15068 19168
rect 15016 19125 15025 19159
rect 15025 19125 15059 19159
rect 15059 19125 15068 19159
rect 15016 19116 15068 19125
rect 15844 19116 15896 19168
rect 26240 19184 26292 19236
rect 27436 19184 27488 19236
rect 29552 19184 29604 19236
rect 31300 19363 31352 19372
rect 31300 19329 31309 19363
rect 31309 19329 31343 19363
rect 31343 19329 31352 19363
rect 31300 19320 31352 19329
rect 32128 19320 32180 19372
rect 33232 19320 33284 19372
rect 34244 19320 34296 19372
rect 35992 19320 36044 19372
rect 39672 19456 39724 19508
rect 41696 19499 41748 19508
rect 41696 19465 41705 19499
rect 41705 19465 41739 19499
rect 41739 19465 41748 19499
rect 41696 19456 41748 19465
rect 37280 19320 37332 19372
rect 18052 19159 18104 19168
rect 18052 19125 18061 19159
rect 18061 19125 18095 19159
rect 18095 19125 18104 19159
rect 21824 19159 21876 19168
rect 18052 19116 18104 19125
rect 21824 19125 21833 19159
rect 21833 19125 21867 19159
rect 21867 19125 21876 19159
rect 21824 19116 21876 19125
rect 25780 19116 25832 19168
rect 30748 19159 30800 19168
rect 30748 19125 30757 19159
rect 30757 19125 30791 19159
rect 30791 19125 30800 19159
rect 30748 19116 30800 19125
rect 30840 19116 30892 19168
rect 36912 19252 36964 19304
rect 40408 19320 40460 19372
rect 39948 19252 40000 19304
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 5264 18912 5316 18964
rect 6644 18912 6696 18964
rect 3792 18844 3844 18896
rect 12164 18912 12216 18964
rect 14372 18912 14424 18964
rect 16764 18912 16816 18964
rect 4896 18776 4948 18828
rect 2872 18708 2924 18760
rect 4712 18708 4764 18760
rect 12716 18844 12768 18896
rect 8300 18776 8352 18828
rect 8668 18776 8720 18828
rect 9588 18776 9640 18828
rect 11244 18708 11296 18760
rect 12532 18708 12584 18760
rect 2412 18640 2464 18692
rect 5356 18640 5408 18692
rect 6000 18640 6052 18692
rect 6184 18683 6236 18692
rect 6184 18649 6193 18683
rect 6193 18649 6227 18683
rect 6227 18649 6236 18683
rect 6184 18640 6236 18649
rect 6920 18640 6972 18692
rect 11520 18640 11572 18692
rect 13820 18708 13872 18760
rect 17776 18776 17828 18828
rect 25780 18955 25832 18964
rect 25780 18921 25789 18955
rect 25789 18921 25823 18955
rect 25823 18921 25832 18955
rect 25780 18912 25832 18921
rect 26148 18912 26200 18964
rect 28356 18912 28408 18964
rect 33232 18912 33284 18964
rect 40408 18955 40460 18964
rect 40408 18921 40417 18955
rect 40417 18921 40451 18955
rect 40451 18921 40460 18955
rect 40408 18912 40460 18921
rect 16764 18751 16816 18760
rect 16764 18717 16773 18751
rect 16773 18717 16807 18751
rect 16807 18717 16816 18751
rect 16764 18708 16816 18717
rect 17040 18708 17092 18760
rect 17868 18751 17920 18760
rect 17868 18717 17877 18751
rect 17877 18717 17911 18751
rect 17911 18717 17920 18751
rect 17868 18708 17920 18717
rect 18144 18708 18196 18760
rect 19248 18751 19300 18760
rect 19248 18717 19257 18751
rect 19257 18717 19291 18751
rect 19291 18717 19300 18751
rect 19248 18708 19300 18717
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 4528 18572 4580 18624
rect 6736 18572 6788 18624
rect 11612 18615 11664 18624
rect 11612 18581 11621 18615
rect 11621 18581 11655 18615
rect 11655 18581 11664 18615
rect 11612 18572 11664 18581
rect 11980 18572 12032 18624
rect 18788 18572 18840 18624
rect 31300 18844 31352 18896
rect 36084 18887 36136 18896
rect 22100 18776 22152 18828
rect 22192 18776 22244 18828
rect 23848 18776 23900 18828
rect 23940 18776 23992 18828
rect 26240 18776 26292 18828
rect 24584 18708 24636 18760
rect 25412 18751 25464 18760
rect 25412 18717 25421 18751
rect 25421 18717 25455 18751
rect 25455 18717 25464 18751
rect 25412 18708 25464 18717
rect 25596 18751 25648 18760
rect 25596 18717 25605 18751
rect 25605 18717 25639 18751
rect 25639 18717 25648 18751
rect 25596 18708 25648 18717
rect 26332 18708 26384 18760
rect 29736 18751 29788 18760
rect 29736 18717 29745 18751
rect 29745 18717 29779 18751
rect 29779 18717 29788 18751
rect 29736 18708 29788 18717
rect 29920 18751 29972 18760
rect 29920 18717 29929 18751
rect 29929 18717 29963 18751
rect 29963 18717 29972 18751
rect 29920 18708 29972 18717
rect 30932 18776 30984 18828
rect 30840 18751 30892 18760
rect 30840 18717 30849 18751
rect 30849 18717 30883 18751
rect 30883 18717 30892 18751
rect 31024 18751 31076 18760
rect 30840 18708 30892 18717
rect 31024 18717 31033 18751
rect 31033 18717 31067 18751
rect 31067 18717 31076 18751
rect 31024 18708 31076 18717
rect 25504 18683 25556 18692
rect 25504 18649 25513 18683
rect 25513 18649 25547 18683
rect 25547 18649 25556 18683
rect 25504 18640 25556 18649
rect 26792 18640 26844 18692
rect 27436 18640 27488 18692
rect 29828 18683 29880 18692
rect 29828 18649 29837 18683
rect 29837 18649 29871 18683
rect 29871 18649 29880 18683
rect 36084 18853 36093 18887
rect 36093 18853 36127 18887
rect 36127 18853 36136 18887
rect 36084 18844 36136 18853
rect 32312 18751 32364 18760
rect 32312 18717 32321 18751
rect 32321 18717 32355 18751
rect 32355 18717 32364 18751
rect 32312 18708 32364 18717
rect 35992 18708 36044 18760
rect 36452 18751 36504 18760
rect 36452 18717 36461 18751
rect 36461 18717 36495 18751
rect 36495 18717 36504 18751
rect 36452 18708 36504 18717
rect 36636 18751 36688 18760
rect 36636 18717 36645 18751
rect 36645 18717 36679 18751
rect 36679 18717 36688 18751
rect 36636 18708 36688 18717
rect 40500 18708 40552 18760
rect 40776 18751 40828 18760
rect 40776 18717 40785 18751
rect 40785 18717 40819 18751
rect 40819 18717 40828 18751
rect 40776 18708 40828 18717
rect 41144 18708 41196 18760
rect 41696 18751 41748 18760
rect 41696 18717 41705 18751
rect 41705 18717 41739 18751
rect 41739 18717 41748 18751
rect 41696 18708 41748 18717
rect 58164 18751 58216 18760
rect 58164 18717 58173 18751
rect 58173 18717 58207 18751
rect 58207 18717 58216 18751
rect 58164 18708 58216 18717
rect 29828 18640 29880 18649
rect 25412 18572 25464 18624
rect 26148 18572 26200 18624
rect 27068 18572 27120 18624
rect 29276 18572 29328 18624
rect 30564 18615 30616 18624
rect 30564 18581 30573 18615
rect 30573 18581 30607 18615
rect 30607 18581 30616 18615
rect 30564 18572 30616 18581
rect 36360 18683 36412 18692
rect 36360 18649 36369 18683
rect 36369 18649 36403 18683
rect 36403 18649 36412 18683
rect 36360 18640 36412 18649
rect 39764 18640 39816 18692
rect 32588 18572 32640 18624
rect 32680 18572 32732 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 2596 18368 2648 18420
rect 4620 18368 4672 18420
rect 9036 18368 9088 18420
rect 3792 18300 3844 18352
rect 6920 18343 6972 18352
rect 6920 18309 6929 18343
rect 6929 18309 6963 18343
rect 6963 18309 6972 18343
rect 6920 18300 6972 18309
rect 8484 18300 8536 18352
rect 9588 18368 9640 18420
rect 11060 18368 11112 18420
rect 11520 18411 11572 18420
rect 11520 18377 11529 18411
rect 11529 18377 11563 18411
rect 11563 18377 11572 18411
rect 11520 18368 11572 18377
rect 11704 18368 11756 18420
rect 5908 18232 5960 18284
rect 6736 18232 6788 18284
rect 7196 18232 7248 18284
rect 7481 18273 7533 18284
rect 7481 18239 7493 18273
rect 7493 18239 7527 18273
rect 7527 18239 7533 18273
rect 7481 18232 7533 18239
rect 7932 18232 7984 18284
rect 4804 18164 4856 18216
rect 5448 18164 5500 18216
rect 7748 18164 7800 18216
rect 2228 18096 2280 18148
rect 5080 18096 5132 18148
rect 11520 18232 11572 18284
rect 12072 18300 12124 18352
rect 12440 18300 12492 18352
rect 11980 18275 12032 18284
rect 11980 18241 11989 18275
rect 11989 18241 12023 18275
rect 12023 18241 12032 18275
rect 12164 18275 12216 18284
rect 11980 18232 12032 18241
rect 12164 18241 12173 18275
rect 12173 18241 12207 18275
rect 12207 18241 12216 18275
rect 12164 18232 12216 18241
rect 8484 18164 8536 18216
rect 16764 18300 16816 18352
rect 17868 18300 17920 18352
rect 18788 18343 18840 18352
rect 18788 18309 18797 18343
rect 18797 18309 18831 18343
rect 18831 18309 18840 18343
rect 18788 18300 18840 18309
rect 19248 18300 19300 18352
rect 23940 18343 23992 18352
rect 13452 18275 13504 18284
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 13636 18275 13688 18284
rect 13636 18241 13645 18275
rect 13645 18241 13679 18275
rect 13679 18241 13688 18275
rect 13636 18232 13688 18241
rect 3700 18071 3752 18080
rect 3700 18037 3709 18071
rect 3709 18037 3743 18071
rect 3743 18037 3752 18071
rect 3700 18028 3752 18037
rect 5356 18028 5408 18080
rect 6184 18028 6236 18080
rect 10968 18096 11020 18148
rect 11244 18096 11296 18148
rect 12532 18096 12584 18148
rect 13820 18275 13872 18284
rect 13820 18241 13829 18275
rect 13829 18241 13863 18275
rect 13863 18241 13872 18275
rect 13820 18232 13872 18241
rect 19340 18232 19392 18284
rect 17960 18164 18012 18216
rect 18144 18164 18196 18216
rect 17868 18096 17920 18148
rect 22376 18232 22428 18284
rect 21272 18207 21324 18216
rect 21272 18173 21281 18207
rect 21281 18173 21315 18207
rect 21315 18173 21324 18207
rect 21272 18164 21324 18173
rect 23940 18309 23949 18343
rect 23949 18309 23983 18343
rect 23983 18309 23992 18343
rect 23940 18300 23992 18309
rect 25504 18368 25556 18420
rect 25964 18368 26016 18420
rect 26332 18368 26384 18420
rect 28540 18368 28592 18420
rect 32588 18411 32640 18420
rect 32588 18377 32597 18411
rect 32597 18377 32631 18411
rect 32631 18377 32640 18411
rect 32588 18368 32640 18377
rect 30196 18300 30248 18352
rect 31944 18300 31996 18352
rect 32404 18343 32456 18352
rect 25688 18232 25740 18284
rect 32404 18309 32413 18343
rect 32413 18309 32447 18343
rect 32447 18309 32456 18343
rect 32404 18300 32456 18309
rect 33876 18368 33928 18420
rect 38752 18411 38804 18420
rect 38752 18377 38761 18411
rect 38761 18377 38795 18411
rect 38795 18377 38804 18411
rect 38752 18368 38804 18377
rect 34152 18300 34204 18352
rect 23204 18164 23256 18216
rect 28540 18164 28592 18216
rect 38476 18232 38528 18284
rect 38936 18232 38988 18284
rect 33784 18164 33836 18216
rect 37648 18164 37700 18216
rect 40500 18232 40552 18284
rect 40960 18275 41012 18284
rect 40960 18241 40969 18275
rect 40969 18241 41003 18275
rect 41003 18241 41012 18275
rect 40960 18232 41012 18241
rect 41052 18275 41104 18284
rect 41052 18241 41061 18275
rect 41061 18241 41095 18275
rect 41095 18241 41104 18275
rect 41052 18232 41104 18241
rect 32956 18096 33008 18148
rect 15200 18028 15252 18080
rect 15844 18028 15896 18080
rect 20444 18028 20496 18080
rect 20904 18028 20956 18080
rect 24676 18028 24728 18080
rect 30748 18028 30800 18080
rect 33048 18071 33100 18080
rect 33048 18037 33057 18071
rect 33057 18037 33091 18071
rect 33091 18037 33100 18071
rect 33048 18028 33100 18037
rect 35624 18028 35676 18080
rect 38936 18028 38988 18080
rect 39948 18028 40000 18080
rect 40868 18096 40920 18148
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4068 17824 4120 17876
rect 4712 17756 4764 17808
rect 4988 17756 5040 17808
rect 5264 17756 5316 17808
rect 5448 17867 5500 17876
rect 5448 17833 5457 17867
rect 5457 17833 5491 17867
rect 5491 17833 5500 17867
rect 9036 17867 9088 17876
rect 5448 17824 5500 17833
rect 9036 17833 9045 17867
rect 9045 17833 9079 17867
rect 9079 17833 9088 17867
rect 9036 17824 9088 17833
rect 9404 17824 9456 17876
rect 5632 17620 5684 17672
rect 10876 17824 10928 17876
rect 11152 17824 11204 17876
rect 13636 17824 13688 17876
rect 21916 17824 21968 17876
rect 25688 17867 25740 17876
rect 25688 17833 25697 17867
rect 25697 17833 25731 17867
rect 25731 17833 25740 17867
rect 25688 17824 25740 17833
rect 31944 17824 31996 17876
rect 36728 17867 36780 17876
rect 25136 17756 25188 17808
rect 26976 17756 27028 17808
rect 34612 17756 34664 17808
rect 35808 17756 35860 17808
rect 36728 17833 36737 17867
rect 36737 17833 36771 17867
rect 36771 17833 36780 17867
rect 36728 17824 36780 17833
rect 41052 17824 41104 17876
rect 37372 17756 37424 17808
rect 40960 17756 41012 17808
rect 16488 17688 16540 17740
rect 20904 17688 20956 17740
rect 12164 17663 12216 17672
rect 12164 17629 12173 17663
rect 12173 17629 12207 17663
rect 12207 17629 12216 17663
rect 12164 17620 12216 17629
rect 4712 17484 4764 17536
rect 5908 17527 5960 17536
rect 5908 17493 5917 17527
rect 5917 17493 5951 17527
rect 5951 17493 5960 17527
rect 5908 17484 5960 17493
rect 7932 17527 7984 17536
rect 7932 17493 7941 17527
rect 7941 17493 7975 17527
rect 7975 17493 7984 17527
rect 7932 17484 7984 17493
rect 11520 17484 11572 17536
rect 11888 17527 11940 17536
rect 11888 17493 11897 17527
rect 11897 17493 11931 17527
rect 11931 17493 11940 17527
rect 11888 17484 11940 17493
rect 12072 17552 12124 17604
rect 12348 17663 12400 17672
rect 12348 17629 12357 17663
rect 12357 17629 12391 17663
rect 12391 17629 12400 17663
rect 12348 17620 12400 17629
rect 12624 17620 12676 17672
rect 13452 17620 13504 17672
rect 15200 17663 15252 17672
rect 15200 17629 15218 17663
rect 15218 17629 15252 17663
rect 15200 17620 15252 17629
rect 21824 17688 21876 17740
rect 23204 17731 23256 17740
rect 23204 17697 23213 17731
rect 23213 17697 23247 17731
rect 23247 17697 23256 17731
rect 23204 17688 23256 17697
rect 13084 17484 13136 17536
rect 20812 17552 20864 17604
rect 14280 17484 14332 17536
rect 21364 17663 21416 17672
rect 21364 17629 21373 17663
rect 21373 17629 21407 17663
rect 21407 17629 21416 17663
rect 21364 17620 21416 17629
rect 22928 17663 22980 17672
rect 22928 17629 22946 17663
rect 22946 17629 22980 17663
rect 24400 17663 24452 17672
rect 22928 17620 22980 17629
rect 24400 17629 24409 17663
rect 24409 17629 24443 17663
rect 24443 17629 24452 17663
rect 24400 17620 24452 17629
rect 23296 17552 23348 17604
rect 25412 17688 25464 17740
rect 24768 17663 24820 17672
rect 24768 17629 24777 17663
rect 24777 17629 24811 17663
rect 24811 17629 24820 17663
rect 24768 17620 24820 17629
rect 25596 17620 25648 17672
rect 25872 17552 25924 17604
rect 21088 17484 21140 17536
rect 26148 17663 26200 17672
rect 26148 17629 26157 17663
rect 26157 17629 26191 17663
rect 26191 17629 26200 17663
rect 26148 17620 26200 17629
rect 26608 17620 26660 17672
rect 28356 17620 28408 17672
rect 31392 17620 31444 17672
rect 32496 17663 32548 17672
rect 32496 17629 32505 17663
rect 32505 17629 32539 17663
rect 32539 17629 32548 17663
rect 32496 17620 32548 17629
rect 33048 17688 33100 17740
rect 40500 17688 40552 17740
rect 27068 17552 27120 17604
rect 28264 17552 28316 17604
rect 32588 17552 32640 17604
rect 32772 17629 32781 17648
rect 32781 17629 32815 17648
rect 32815 17629 32824 17648
rect 32772 17596 32824 17629
rect 35624 17663 35676 17672
rect 26884 17527 26936 17536
rect 26884 17493 26893 17527
rect 26893 17493 26927 17527
rect 26927 17493 26936 17527
rect 26884 17484 26936 17493
rect 31944 17527 31996 17536
rect 31944 17493 31953 17527
rect 31953 17493 31987 17527
rect 31987 17493 31996 17527
rect 35624 17629 35633 17663
rect 35633 17629 35667 17663
rect 35667 17629 35676 17663
rect 35624 17620 35676 17629
rect 35808 17663 35860 17672
rect 35808 17629 35817 17663
rect 35817 17629 35851 17663
rect 35851 17629 35860 17663
rect 35808 17620 35860 17629
rect 35992 17663 36044 17672
rect 35992 17629 36001 17663
rect 36001 17629 36035 17663
rect 36035 17629 36044 17663
rect 35992 17620 36044 17629
rect 37188 17620 37240 17672
rect 37464 17620 37516 17672
rect 38752 17620 38804 17672
rect 33140 17527 33192 17536
rect 31944 17484 31996 17493
rect 33140 17493 33149 17527
rect 33149 17493 33183 17527
rect 33183 17493 33192 17527
rect 33140 17484 33192 17493
rect 35072 17527 35124 17536
rect 35072 17493 35081 17527
rect 35081 17493 35115 17527
rect 35115 17493 35124 17527
rect 35072 17484 35124 17493
rect 35532 17484 35584 17536
rect 35992 17484 36044 17536
rect 36268 17527 36320 17536
rect 36268 17493 36277 17527
rect 36277 17493 36311 17527
rect 36311 17493 36320 17527
rect 36268 17484 36320 17493
rect 36544 17552 36596 17604
rect 37096 17595 37148 17604
rect 37096 17561 37105 17595
rect 37105 17561 37139 17595
rect 37139 17561 37148 17595
rect 37832 17595 37884 17604
rect 37096 17552 37148 17561
rect 37832 17561 37841 17595
rect 37841 17561 37875 17595
rect 37875 17561 37884 17595
rect 37832 17552 37884 17561
rect 38476 17552 38528 17604
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 4620 17280 4672 17332
rect 12348 17280 12400 17332
rect 13912 17280 13964 17332
rect 3700 17212 3752 17264
rect 2872 17144 2924 17196
rect 12624 17212 12676 17264
rect 13084 17212 13136 17264
rect 14188 17255 14240 17264
rect 14188 17221 14197 17255
rect 14197 17221 14231 17255
rect 14231 17221 14240 17255
rect 14188 17212 14240 17221
rect 14556 17212 14608 17264
rect 8024 17144 8076 17196
rect 8668 17187 8720 17196
rect 8668 17153 8677 17187
rect 8677 17153 8711 17187
rect 8711 17153 8720 17187
rect 8668 17144 8720 17153
rect 9128 17144 9180 17196
rect 12440 17144 12492 17196
rect 13820 17144 13872 17196
rect 4712 17119 4764 17128
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4712 17076 4764 17085
rect 5632 17076 5684 17128
rect 14280 17187 14332 17196
rect 14280 17153 14325 17187
rect 14325 17153 14332 17187
rect 14464 17187 14516 17196
rect 14280 17144 14332 17153
rect 14464 17153 14473 17187
rect 14473 17153 14507 17187
rect 14507 17153 14516 17187
rect 14464 17144 14516 17153
rect 17040 17212 17092 17264
rect 17960 17255 18012 17264
rect 17960 17221 17969 17255
rect 17969 17221 18003 17255
rect 18003 17221 18012 17255
rect 17960 17212 18012 17221
rect 25688 17280 25740 17332
rect 26148 17280 26200 17332
rect 26884 17280 26936 17332
rect 15752 17144 15804 17196
rect 16672 17144 16724 17196
rect 25964 17212 26016 17264
rect 18880 17187 18932 17196
rect 18880 17153 18889 17187
rect 18889 17153 18923 17187
rect 18923 17153 18932 17187
rect 18880 17144 18932 17153
rect 20352 17144 20404 17196
rect 22560 17144 22612 17196
rect 24768 17144 24820 17196
rect 24952 17187 25004 17196
rect 24952 17153 24978 17187
rect 24978 17153 25004 17187
rect 24952 17144 25004 17153
rect 31576 17212 31628 17264
rect 32772 17280 32824 17332
rect 33508 17280 33560 17332
rect 34152 17280 34204 17332
rect 35808 17280 35860 17332
rect 33140 17255 33192 17264
rect 26976 17187 27028 17196
rect 26976 17153 26985 17187
rect 26985 17153 27019 17187
rect 27019 17153 27028 17187
rect 26976 17144 27028 17153
rect 14648 17076 14700 17128
rect 15936 17076 15988 17128
rect 6644 16940 6696 16992
rect 7196 16940 7248 16992
rect 11520 16940 11572 16992
rect 16948 17008 17000 17060
rect 17960 17008 18012 17060
rect 18880 17008 18932 17060
rect 23296 17076 23348 17128
rect 23480 17119 23532 17128
rect 23480 17085 23489 17119
rect 23489 17085 23523 17119
rect 23523 17085 23532 17119
rect 23480 17076 23532 17085
rect 25872 17076 25924 17128
rect 30932 17144 30984 17196
rect 33140 17221 33174 17255
rect 33174 17221 33192 17255
rect 33140 17212 33192 17221
rect 35072 17212 35124 17264
rect 34520 17144 34572 17196
rect 39948 17212 40000 17264
rect 37464 17187 37516 17196
rect 37464 17153 37473 17187
rect 37473 17153 37507 17187
rect 37507 17153 37516 17187
rect 37464 17144 37516 17153
rect 37648 17187 37700 17196
rect 37648 17153 37657 17187
rect 37657 17153 37691 17187
rect 37691 17153 37700 17187
rect 37648 17144 37700 17153
rect 39764 17144 39816 17196
rect 21364 16940 21416 16992
rect 21824 16940 21876 16992
rect 23388 16940 23440 16992
rect 25688 17008 25740 17060
rect 29460 17076 29512 17128
rect 30380 17076 30432 17128
rect 32680 17076 32732 17128
rect 39856 17076 39908 17128
rect 28172 17008 28224 17060
rect 33876 17008 33928 17060
rect 58164 17051 58216 17060
rect 58164 17017 58173 17051
rect 58173 17017 58207 17051
rect 58207 17017 58216 17051
rect 58164 17008 58216 17017
rect 25136 16983 25188 16992
rect 25136 16949 25145 16983
rect 25145 16949 25179 16983
rect 25179 16949 25188 16983
rect 25136 16940 25188 16949
rect 27804 16940 27856 16992
rect 28632 16940 28684 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 7288 16736 7340 16788
rect 7748 16736 7800 16788
rect 8024 16779 8076 16788
rect 8024 16745 8033 16779
rect 8033 16745 8067 16779
rect 8067 16745 8076 16779
rect 8024 16736 8076 16745
rect 12164 16736 12216 16788
rect 15752 16736 15804 16788
rect 16304 16736 16356 16788
rect 25872 16779 25924 16788
rect 5632 16668 5684 16720
rect 7380 16668 7432 16720
rect 16764 16668 16816 16720
rect 25872 16745 25881 16779
rect 25881 16745 25915 16779
rect 25915 16745 25924 16779
rect 25872 16736 25924 16745
rect 28356 16736 28408 16788
rect 32312 16736 32364 16788
rect 2504 16532 2556 16584
rect 4344 16532 4396 16584
rect 7288 16575 7340 16584
rect 7288 16541 7297 16575
rect 7297 16541 7331 16575
rect 7331 16541 7340 16575
rect 7288 16532 7340 16541
rect 7472 16575 7524 16584
rect 7472 16541 7481 16575
rect 7481 16541 7515 16575
rect 7515 16541 7524 16575
rect 7472 16532 7524 16541
rect 12624 16600 12676 16652
rect 16304 16600 16356 16652
rect 15752 16575 15804 16584
rect 3976 16464 4028 16516
rect 7196 16464 7248 16516
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 15752 16532 15804 16541
rect 2320 16396 2372 16448
rect 4712 16396 4764 16448
rect 5264 16396 5316 16448
rect 8484 16396 8536 16448
rect 10324 16396 10376 16448
rect 14188 16464 14240 16516
rect 15936 16575 15988 16584
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 15936 16532 15988 16541
rect 16120 16575 16172 16584
rect 16120 16541 16129 16575
rect 16129 16541 16163 16575
rect 16163 16541 16172 16575
rect 17960 16600 18012 16652
rect 21180 16668 21232 16720
rect 20996 16600 21048 16652
rect 22376 16600 22428 16652
rect 22652 16600 22704 16652
rect 27252 16643 27304 16652
rect 27252 16609 27261 16643
rect 27261 16609 27295 16643
rect 27295 16609 27304 16643
rect 27252 16600 27304 16609
rect 27344 16600 27396 16652
rect 27804 16600 27856 16652
rect 16120 16532 16172 16541
rect 16764 16575 16816 16584
rect 16764 16541 16773 16575
rect 16773 16541 16807 16575
rect 16807 16541 16816 16575
rect 16764 16532 16816 16541
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 18236 16575 18288 16584
rect 18236 16541 18245 16575
rect 18245 16541 18279 16575
rect 18279 16541 18288 16575
rect 18236 16532 18288 16541
rect 22560 16575 22612 16584
rect 17776 16464 17828 16516
rect 11152 16439 11204 16448
rect 11152 16405 11161 16439
rect 11161 16405 11195 16439
rect 11195 16405 11204 16439
rect 11152 16396 11204 16405
rect 12808 16396 12860 16448
rect 15384 16396 15436 16448
rect 17224 16439 17276 16448
rect 17224 16405 17233 16439
rect 17233 16405 17267 16439
rect 17267 16405 17276 16439
rect 17224 16396 17276 16405
rect 18052 16396 18104 16448
rect 22560 16541 22569 16575
rect 22569 16541 22603 16575
rect 22603 16541 22612 16575
rect 22560 16532 22612 16541
rect 28172 16575 28224 16584
rect 28172 16541 28181 16575
rect 28181 16541 28215 16575
rect 28215 16541 28224 16575
rect 28172 16532 28224 16541
rect 28356 16575 28408 16584
rect 28356 16541 28365 16575
rect 28365 16541 28399 16575
rect 28399 16541 28408 16575
rect 28356 16532 28408 16541
rect 18696 16439 18748 16448
rect 18696 16405 18705 16439
rect 18705 16405 18739 16439
rect 18739 16405 18748 16439
rect 18696 16396 18748 16405
rect 19432 16439 19484 16448
rect 19432 16405 19441 16439
rect 19441 16405 19475 16439
rect 19475 16405 19484 16439
rect 19432 16396 19484 16405
rect 22100 16439 22152 16448
rect 22100 16405 22109 16439
rect 22109 16405 22143 16439
rect 22143 16405 22152 16439
rect 22100 16396 22152 16405
rect 27160 16396 27212 16448
rect 32680 16600 32732 16652
rect 38108 16736 38160 16788
rect 38200 16736 38252 16788
rect 38936 16779 38988 16788
rect 38936 16745 38945 16779
rect 38945 16745 38979 16779
rect 38979 16745 38988 16779
rect 38936 16736 38988 16745
rect 40776 16736 40828 16788
rect 37464 16668 37516 16720
rect 28632 16532 28684 16584
rect 30380 16464 30432 16516
rect 30564 16464 30616 16516
rect 30932 16532 30984 16584
rect 32036 16532 32088 16584
rect 32496 16532 32548 16584
rect 32956 16575 33008 16584
rect 32956 16541 32965 16575
rect 32965 16541 32999 16575
rect 32999 16541 33008 16575
rect 32956 16532 33008 16541
rect 31484 16464 31536 16516
rect 32312 16507 32364 16516
rect 32312 16473 32321 16507
rect 32321 16473 32355 16507
rect 32355 16473 32364 16507
rect 33968 16532 34020 16584
rect 36268 16575 36320 16584
rect 36268 16541 36302 16575
rect 36302 16541 36320 16575
rect 36268 16532 36320 16541
rect 32312 16464 32364 16473
rect 34520 16464 34572 16516
rect 40500 16464 40552 16516
rect 29828 16396 29880 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 4344 16235 4396 16244
rect 4344 16201 4353 16235
rect 4353 16201 4387 16235
rect 4387 16201 4396 16235
rect 4344 16192 4396 16201
rect 2872 16124 2924 16176
rect 6184 16192 6236 16244
rect 10876 16235 10928 16244
rect 10876 16201 10885 16235
rect 10885 16201 10919 16235
rect 10919 16201 10928 16235
rect 10876 16192 10928 16201
rect 13728 16192 13780 16244
rect 15936 16192 15988 16244
rect 16764 16192 16816 16244
rect 18236 16192 18288 16244
rect 26332 16192 26384 16244
rect 26976 16192 27028 16244
rect 31392 16192 31444 16244
rect 31484 16192 31536 16244
rect 15016 16124 15068 16176
rect 16120 16167 16172 16176
rect 16120 16133 16129 16167
rect 16129 16133 16163 16167
rect 16163 16133 16172 16167
rect 16120 16124 16172 16133
rect 19340 16124 19392 16176
rect 19892 16124 19944 16176
rect 2320 16099 2372 16108
rect 2320 16065 2354 16099
rect 2354 16065 2372 16099
rect 2320 16056 2372 16065
rect 10324 16099 10376 16108
rect 4712 15988 4764 16040
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 11428 16056 11480 16108
rect 11612 16099 11664 16108
rect 11612 16065 11622 16099
rect 11622 16065 11656 16099
rect 11656 16065 11664 16099
rect 11612 16056 11664 16065
rect 11796 16099 11848 16108
rect 11796 16065 11805 16099
rect 11805 16065 11839 16099
rect 11839 16065 11848 16099
rect 11796 16056 11848 16065
rect 11980 16056 12032 16108
rect 12624 16099 12676 16108
rect 10784 15920 10836 15972
rect 11152 15988 11204 16040
rect 11704 15988 11756 16040
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 13820 16056 13872 16108
rect 14280 16099 14332 16108
rect 14280 16065 14289 16099
rect 14289 16065 14323 16099
rect 14323 16065 14332 16099
rect 14280 16056 14332 16065
rect 14648 16056 14700 16108
rect 16948 16056 17000 16108
rect 18236 16056 18288 16108
rect 14556 16031 14608 16040
rect 14556 15997 14565 16031
rect 14565 15997 14599 16031
rect 14599 15997 14608 16031
rect 14556 15988 14608 15997
rect 19432 15988 19484 16040
rect 19892 16031 19944 16040
rect 19892 15997 19901 16031
rect 19901 15997 19935 16031
rect 19935 15997 19944 16031
rect 19892 15988 19944 15997
rect 20076 16099 20128 16108
rect 20076 16065 20085 16099
rect 20085 16065 20119 16099
rect 20119 16065 20128 16099
rect 20076 16056 20128 16065
rect 20628 15988 20680 16040
rect 20996 16056 21048 16108
rect 23480 16056 23532 16108
rect 26240 16124 26292 16176
rect 21180 15988 21232 16040
rect 27160 16056 27212 16108
rect 27528 16031 27580 16040
rect 3884 15895 3936 15904
rect 3884 15861 3893 15895
rect 3893 15861 3927 15895
rect 3927 15861 3936 15895
rect 3884 15852 3936 15861
rect 7104 15895 7156 15904
rect 7104 15861 7113 15895
rect 7113 15861 7147 15895
rect 7147 15861 7156 15895
rect 7104 15852 7156 15861
rect 9680 15852 9732 15904
rect 14188 15920 14240 15972
rect 22100 15920 22152 15972
rect 23204 15920 23256 15972
rect 27528 15997 27537 16031
rect 27537 15997 27571 16031
rect 27571 15997 27580 16031
rect 27528 15988 27580 15997
rect 27160 15920 27212 15972
rect 29828 16056 29880 16108
rect 30380 16056 30432 16108
rect 31392 16099 31444 16108
rect 31392 16065 31401 16099
rect 31401 16065 31435 16099
rect 31435 16065 31444 16099
rect 31392 16056 31444 16065
rect 29920 15988 29972 16040
rect 30656 15988 30708 16040
rect 30932 15988 30984 16040
rect 29828 15920 29880 15972
rect 12808 15852 12860 15904
rect 21456 15852 21508 15904
rect 22192 15852 22244 15904
rect 30380 15852 30432 15904
rect 32588 15852 32640 15904
rect 37372 16192 37424 16244
rect 39948 16192 40000 16244
rect 35348 15988 35400 16040
rect 37096 16124 37148 16176
rect 37188 16056 37240 16108
rect 38660 16056 38712 16108
rect 40132 16056 40184 16108
rect 38752 15920 38804 15972
rect 36912 15852 36964 15904
rect 38936 15852 38988 15904
rect 58164 15895 58216 15904
rect 58164 15861 58173 15895
rect 58173 15861 58207 15895
rect 58207 15861 58216 15895
rect 58164 15852 58216 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2504 15691 2556 15700
rect 2504 15657 2513 15691
rect 2513 15657 2547 15691
rect 2547 15657 2556 15691
rect 2504 15648 2556 15657
rect 6828 15691 6880 15700
rect 6828 15657 6837 15691
rect 6837 15657 6871 15691
rect 6871 15657 6880 15691
rect 6828 15648 6880 15657
rect 7840 15648 7892 15700
rect 9312 15691 9364 15700
rect 9312 15657 9321 15691
rect 9321 15657 9355 15691
rect 9355 15657 9364 15691
rect 9312 15648 9364 15657
rect 6460 15580 6512 15632
rect 7104 15512 7156 15564
rect 7564 15512 7616 15564
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 3884 15444 3936 15496
rect 7656 15487 7708 15496
rect 5080 15376 5132 15428
rect 6736 15376 6788 15428
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 9404 15487 9456 15496
rect 9404 15453 9413 15487
rect 9413 15453 9447 15487
rect 9447 15453 9456 15487
rect 9404 15444 9456 15453
rect 9680 15444 9732 15496
rect 11980 15648 12032 15700
rect 12440 15691 12492 15700
rect 12440 15657 12449 15691
rect 12449 15657 12483 15691
rect 12483 15657 12492 15691
rect 14280 15691 14332 15700
rect 12440 15648 12492 15657
rect 14280 15657 14289 15691
rect 14289 15657 14323 15691
rect 14323 15657 14332 15691
rect 14280 15648 14332 15657
rect 21548 15648 21600 15700
rect 22560 15648 22612 15700
rect 23480 15648 23532 15700
rect 27068 15691 27120 15700
rect 27068 15657 27077 15691
rect 27077 15657 27111 15691
rect 27111 15657 27120 15691
rect 27068 15648 27120 15657
rect 29552 15691 29604 15700
rect 29552 15657 29561 15691
rect 29561 15657 29595 15691
rect 29595 15657 29604 15691
rect 29552 15648 29604 15657
rect 30656 15648 30708 15700
rect 32588 15691 32640 15700
rect 10876 15512 10928 15564
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 30932 15580 30984 15632
rect 10508 15487 10560 15496
rect 10508 15453 10516 15487
rect 10516 15453 10550 15487
rect 10550 15453 10560 15487
rect 10508 15444 10560 15453
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 11888 15444 11940 15496
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 14556 15512 14608 15564
rect 19248 15555 19300 15564
rect 19248 15521 19257 15555
rect 19257 15521 19291 15555
rect 19291 15521 19300 15555
rect 19248 15512 19300 15521
rect 20996 15512 21048 15564
rect 6552 15351 6604 15360
rect 6552 15317 6561 15351
rect 6561 15317 6595 15351
rect 6595 15317 6604 15351
rect 6552 15308 6604 15317
rect 8392 15308 8444 15360
rect 11796 15376 11848 15428
rect 13820 15444 13872 15496
rect 13268 15419 13320 15428
rect 13268 15385 13277 15419
rect 13277 15385 13311 15419
rect 13311 15385 13320 15419
rect 14188 15444 14240 15496
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 15384 15487 15436 15496
rect 15384 15453 15418 15487
rect 15418 15453 15436 15487
rect 15384 15444 15436 15453
rect 18696 15444 18748 15496
rect 21272 15487 21324 15496
rect 13268 15376 13320 15385
rect 14372 15376 14424 15428
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 22100 15444 22152 15496
rect 23296 15487 23348 15496
rect 21180 15376 21232 15428
rect 22192 15376 22244 15428
rect 23296 15453 23305 15487
rect 23305 15453 23339 15487
rect 23339 15453 23348 15487
rect 23296 15444 23348 15453
rect 26976 15487 27028 15496
rect 26976 15453 26985 15487
rect 26985 15453 27019 15487
rect 27019 15453 27028 15487
rect 26976 15444 27028 15453
rect 27160 15487 27212 15496
rect 27160 15453 27169 15487
rect 27169 15453 27203 15487
rect 27203 15453 27212 15487
rect 27160 15444 27212 15453
rect 32588 15657 32597 15691
rect 32597 15657 32631 15691
rect 32631 15657 32640 15691
rect 32588 15648 32640 15657
rect 36912 15691 36964 15700
rect 36912 15657 36921 15691
rect 36921 15657 36955 15691
rect 36955 15657 36964 15691
rect 36912 15648 36964 15657
rect 40132 15648 40184 15700
rect 39580 15580 39632 15632
rect 40500 15580 40552 15632
rect 31024 15444 31076 15496
rect 37188 15512 37240 15564
rect 37832 15512 37884 15564
rect 32036 15487 32088 15496
rect 31484 15376 31536 15428
rect 32036 15453 32045 15487
rect 32045 15453 32079 15487
rect 32079 15453 32088 15487
rect 32036 15444 32088 15453
rect 33232 15444 33284 15496
rect 33600 15487 33652 15496
rect 33600 15453 33609 15487
rect 33609 15453 33643 15487
rect 33643 15453 33652 15487
rect 33600 15444 33652 15453
rect 34704 15444 34756 15496
rect 37648 15444 37700 15496
rect 38200 15487 38252 15496
rect 38200 15453 38209 15487
rect 38209 15453 38243 15487
rect 38243 15453 38252 15487
rect 38200 15444 38252 15453
rect 38752 15444 38804 15496
rect 40684 15487 40736 15496
rect 40684 15453 40693 15487
rect 40693 15453 40727 15487
rect 40727 15453 40736 15487
rect 40684 15444 40736 15453
rect 41144 15487 41196 15496
rect 41144 15453 41153 15487
rect 41153 15453 41187 15487
rect 41187 15453 41196 15487
rect 41144 15444 41196 15453
rect 41328 15487 41380 15496
rect 41328 15453 41337 15487
rect 41337 15453 41371 15487
rect 41371 15453 41380 15487
rect 41328 15444 41380 15453
rect 41512 15487 41564 15496
rect 41512 15453 41521 15487
rect 41521 15453 41555 15487
rect 41555 15453 41564 15487
rect 41512 15444 41564 15453
rect 16948 15308 17000 15360
rect 18788 15308 18840 15360
rect 20628 15351 20680 15360
rect 20628 15317 20637 15351
rect 20637 15317 20671 15351
rect 20671 15317 20680 15351
rect 20628 15308 20680 15317
rect 21916 15351 21968 15360
rect 21916 15317 21925 15351
rect 21925 15317 21959 15351
rect 21959 15317 21968 15351
rect 21916 15308 21968 15317
rect 22744 15308 22796 15360
rect 38660 15308 38712 15360
rect 38844 15351 38896 15360
rect 38844 15317 38853 15351
rect 38853 15317 38887 15351
rect 38887 15317 38896 15351
rect 38844 15308 38896 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 6736 15036 6788 15088
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 2872 14968 2924 15020
rect 5632 15011 5684 15020
rect 5632 14977 5641 15011
rect 5641 14977 5675 15011
rect 5675 14977 5684 15011
rect 5632 14968 5684 14977
rect 6368 15011 6420 15020
rect 6368 14977 6377 15011
rect 6377 14977 6411 15011
rect 6411 14977 6420 15011
rect 6368 14968 6420 14977
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 6644 15011 6696 15020
rect 6644 14977 6653 15011
rect 6653 14977 6687 15011
rect 6687 14977 6696 15011
rect 6644 14968 6696 14977
rect 9128 15011 9180 15020
rect 9128 14977 9137 15011
rect 9137 14977 9171 15011
rect 9171 14977 9180 15011
rect 9128 14968 9180 14977
rect 12808 15104 12860 15156
rect 13084 15104 13136 15156
rect 16672 15036 16724 15088
rect 17224 15036 17276 15088
rect 18512 15104 18564 15156
rect 24216 15147 24268 15156
rect 24216 15113 24225 15147
rect 24225 15113 24259 15147
rect 24259 15113 24268 15147
rect 24216 15104 24268 15113
rect 25044 15147 25096 15156
rect 25044 15113 25053 15147
rect 25053 15113 25087 15147
rect 25087 15113 25096 15147
rect 25044 15104 25096 15113
rect 25596 15104 25648 15156
rect 27620 15104 27672 15156
rect 28264 15147 28316 15156
rect 28264 15113 28273 15147
rect 28273 15113 28307 15147
rect 28307 15113 28316 15147
rect 28264 15104 28316 15113
rect 30564 15104 30616 15156
rect 37832 15104 37884 15156
rect 38568 15104 38620 15156
rect 38660 15104 38712 15156
rect 10140 15011 10192 15020
rect 10140 14977 10149 15011
rect 10149 14977 10183 15011
rect 10183 14977 10192 15011
rect 10140 14968 10192 14977
rect 11060 14968 11112 15020
rect 11980 14968 12032 15020
rect 22100 15036 22152 15088
rect 18788 14968 18840 15020
rect 20076 14968 20128 15020
rect 22744 15011 22796 15020
rect 22744 14977 22753 15011
rect 22753 14977 22787 15011
rect 22787 14977 22796 15011
rect 22744 14968 22796 14977
rect 2228 14900 2280 14952
rect 2688 14900 2740 14952
rect 2596 14764 2648 14816
rect 5264 14900 5316 14952
rect 3792 14764 3844 14816
rect 4988 14764 5040 14816
rect 7380 14900 7432 14952
rect 9772 14832 9824 14884
rect 10048 14943 10100 14952
rect 10048 14909 10057 14943
rect 10057 14909 10091 14943
rect 10091 14909 10100 14943
rect 10048 14900 10100 14909
rect 15108 14900 15160 14952
rect 16856 14943 16908 14952
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 20168 14943 20220 14952
rect 20168 14909 20177 14943
rect 20177 14909 20211 14943
rect 20211 14909 20220 14943
rect 20168 14900 20220 14909
rect 22192 14900 22244 14952
rect 23296 14968 23348 15020
rect 24124 14968 24176 15020
rect 27620 14968 27672 15020
rect 29644 14968 29696 15020
rect 29828 14900 29880 14952
rect 29920 14900 29972 14952
rect 30380 15011 30432 15020
rect 30380 14977 30389 15011
rect 30389 14977 30423 15011
rect 30423 14977 30432 15011
rect 30380 14968 30432 14977
rect 30564 15011 30616 15020
rect 30564 14977 30573 15011
rect 30573 14977 30607 15011
rect 30607 14977 30616 15011
rect 30564 14968 30616 14977
rect 32036 14968 32088 15020
rect 38844 15036 38896 15088
rect 35348 15011 35400 15020
rect 35348 14977 35357 15011
rect 35357 14977 35391 15011
rect 35391 14977 35400 15011
rect 35348 14968 35400 14977
rect 35716 14968 35768 15020
rect 35624 14900 35676 14952
rect 35808 14943 35860 14952
rect 35808 14909 35817 14943
rect 35817 14909 35851 14943
rect 35851 14909 35860 14943
rect 35808 14900 35860 14909
rect 13820 14832 13872 14884
rect 18236 14875 18288 14884
rect 5816 14807 5868 14816
rect 5816 14773 5825 14807
rect 5825 14773 5859 14807
rect 5859 14773 5868 14807
rect 5816 14764 5868 14773
rect 7104 14807 7156 14816
rect 7104 14773 7113 14807
rect 7113 14773 7147 14807
rect 7147 14773 7156 14807
rect 7104 14764 7156 14773
rect 14372 14764 14424 14816
rect 18236 14841 18245 14875
rect 18245 14841 18279 14875
rect 18279 14841 18288 14875
rect 18236 14832 18288 14841
rect 22836 14832 22888 14884
rect 34704 14832 34756 14884
rect 37464 15011 37516 15020
rect 37464 14977 37473 15011
rect 37473 14977 37507 15011
rect 37507 14977 37516 15011
rect 37464 14968 37516 14977
rect 38752 14968 38804 15020
rect 41512 14968 41564 15020
rect 38108 14900 38160 14952
rect 20352 14764 20404 14816
rect 20812 14764 20864 14816
rect 20996 14764 21048 14816
rect 22192 14764 22244 14816
rect 23480 14764 23532 14816
rect 26976 14764 27028 14816
rect 27712 14764 27764 14816
rect 29644 14764 29696 14816
rect 31024 14764 31076 14816
rect 33232 14807 33284 14816
rect 33232 14773 33241 14807
rect 33241 14773 33275 14807
rect 33275 14773 33284 14807
rect 33232 14764 33284 14773
rect 36728 14764 36780 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 2872 14560 2924 14612
rect 5816 14560 5868 14612
rect 10048 14560 10100 14612
rect 10232 14560 10284 14612
rect 16580 14560 16632 14612
rect 2136 14492 2188 14544
rect 4896 14492 4948 14544
rect 6736 14492 6788 14544
rect 18788 14560 18840 14612
rect 19616 14560 19668 14612
rect 20812 14560 20864 14612
rect 20996 14560 21048 14612
rect 31484 14560 31536 14612
rect 41328 14560 41380 14612
rect 4988 14467 5040 14476
rect 4988 14433 4997 14467
rect 4997 14433 5031 14467
rect 5031 14433 5040 14467
rect 4988 14424 5040 14433
rect 6000 14424 6052 14476
rect 9680 14424 9732 14476
rect 16948 14492 17000 14544
rect 2596 14399 2648 14408
rect 2596 14365 2605 14399
rect 2605 14365 2639 14399
rect 2639 14365 2648 14399
rect 2596 14356 2648 14365
rect 7104 14356 7156 14408
rect 7748 14399 7800 14408
rect 7748 14365 7757 14399
rect 7757 14365 7791 14399
rect 7791 14365 7800 14399
rect 7748 14356 7800 14365
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 14372 14356 14424 14408
rect 19340 14356 19392 14408
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 20168 14399 20220 14408
rect 20168 14365 20177 14399
rect 20177 14365 20211 14399
rect 20211 14365 20220 14399
rect 20168 14356 20220 14365
rect 20352 14399 20404 14408
rect 20352 14365 20361 14399
rect 20361 14365 20395 14399
rect 20395 14365 20404 14399
rect 20352 14356 20404 14365
rect 21364 14356 21416 14408
rect 24952 14492 25004 14544
rect 26976 14492 27028 14544
rect 22560 14424 22612 14476
rect 22652 14356 22704 14408
rect 22836 14399 22888 14408
rect 22836 14365 22845 14399
rect 22845 14365 22879 14399
rect 22879 14365 22888 14399
rect 22836 14356 22888 14365
rect 24124 14424 24176 14476
rect 24400 14424 24452 14476
rect 23204 14399 23256 14408
rect 23204 14365 23213 14399
rect 23213 14365 23247 14399
rect 23247 14365 23256 14399
rect 23204 14356 23256 14365
rect 24768 14356 24820 14408
rect 25044 14356 25096 14408
rect 26976 14356 27028 14408
rect 27528 14399 27580 14408
rect 27528 14365 27537 14399
rect 27537 14365 27571 14399
rect 27571 14365 27580 14399
rect 27528 14356 27580 14365
rect 5816 14263 5868 14272
rect 5816 14229 5825 14263
rect 5825 14229 5859 14263
rect 5859 14229 5868 14263
rect 5816 14220 5868 14229
rect 9680 14263 9732 14272
rect 9680 14229 9689 14263
rect 9689 14229 9723 14263
rect 9723 14229 9732 14263
rect 9680 14220 9732 14229
rect 10784 14220 10836 14272
rect 12072 14263 12124 14272
rect 12072 14229 12081 14263
rect 12081 14229 12115 14263
rect 12115 14229 12124 14263
rect 12072 14220 12124 14229
rect 13636 14220 13688 14272
rect 21732 14288 21784 14340
rect 21916 14288 21968 14340
rect 23296 14288 23348 14340
rect 23940 14220 23992 14272
rect 24308 14220 24360 14272
rect 28264 14356 28316 14408
rect 29368 14356 29420 14408
rect 29828 14399 29880 14408
rect 29828 14365 29837 14399
rect 29837 14365 29871 14399
rect 29871 14365 29880 14399
rect 29828 14356 29880 14365
rect 40868 14492 40920 14544
rect 32036 14424 32088 14476
rect 33600 14424 33652 14476
rect 34704 14467 34756 14476
rect 34704 14433 34713 14467
rect 34713 14433 34747 14467
rect 34747 14433 34756 14467
rect 34704 14424 34756 14433
rect 35808 14424 35860 14476
rect 33416 14356 33468 14408
rect 34796 14356 34848 14408
rect 35716 14356 35768 14408
rect 27804 14288 27856 14340
rect 29552 14288 29604 14340
rect 36912 14356 36964 14408
rect 37188 14399 37240 14408
rect 37188 14365 37197 14399
rect 37197 14365 37231 14399
rect 37231 14365 37240 14399
rect 37188 14356 37240 14365
rect 38936 14356 38988 14408
rect 40684 14356 40736 14408
rect 58164 14399 58216 14408
rect 58164 14365 58173 14399
rect 58173 14365 58207 14399
rect 58207 14365 58216 14399
rect 58164 14356 58216 14365
rect 39488 14288 39540 14340
rect 39856 14331 39908 14340
rect 39856 14297 39865 14331
rect 39865 14297 39899 14331
rect 39899 14297 39908 14331
rect 39856 14288 39908 14297
rect 35716 14220 35768 14272
rect 37648 14220 37700 14272
rect 38108 14220 38160 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 2688 14016 2740 14068
rect 19340 14059 19392 14068
rect 19340 14025 19349 14059
rect 19349 14025 19383 14059
rect 19383 14025 19392 14059
rect 19340 14016 19392 14025
rect 21272 14016 21324 14068
rect 22100 14059 22152 14068
rect 22100 14025 22109 14059
rect 22109 14025 22143 14059
rect 22143 14025 22152 14059
rect 22100 14016 22152 14025
rect 22560 14016 22612 14068
rect 23664 14059 23716 14068
rect 10784 13948 10836 14000
rect 22192 13948 22244 14000
rect 23664 14025 23673 14059
rect 23673 14025 23707 14059
rect 23707 14025 23716 14059
rect 23664 14016 23716 14025
rect 23940 14016 23992 14068
rect 24584 14059 24636 14068
rect 23296 13948 23348 14000
rect 24216 13948 24268 14000
rect 24584 14025 24593 14059
rect 24593 14025 24627 14059
rect 24627 14025 24636 14059
rect 24584 14016 24636 14025
rect 25596 14059 25648 14068
rect 25596 14025 25605 14059
rect 25605 14025 25639 14059
rect 25639 14025 25648 14059
rect 25596 14016 25648 14025
rect 26608 14016 26660 14068
rect 27528 14016 27580 14068
rect 27620 14016 27672 14068
rect 4620 13880 4672 13932
rect 6368 13880 6420 13932
rect 12072 13880 12124 13932
rect 14280 13923 14332 13932
rect 14280 13889 14298 13923
rect 14298 13889 14332 13923
rect 14280 13880 14332 13889
rect 15108 13880 15160 13932
rect 20628 13880 20680 13932
rect 22652 13880 22704 13932
rect 23204 13880 23256 13932
rect 24492 13880 24544 13932
rect 3792 13812 3844 13864
rect 7748 13812 7800 13864
rect 21364 13812 21416 13864
rect 23480 13812 23532 13864
rect 23572 13812 23624 13864
rect 25596 13880 25648 13932
rect 26148 13880 26200 13932
rect 26976 13923 27028 13932
rect 26976 13889 26985 13923
rect 26985 13889 27019 13923
rect 27019 13889 27028 13923
rect 26976 13880 27028 13889
rect 27252 13923 27304 13932
rect 27252 13889 27286 13923
rect 27286 13889 27304 13923
rect 27252 13880 27304 13889
rect 24860 13855 24912 13864
rect 24860 13821 24869 13855
rect 24869 13821 24903 13855
rect 24903 13821 24912 13855
rect 24860 13812 24912 13821
rect 30380 13880 30432 13932
rect 30932 13923 30984 13932
rect 30932 13889 30941 13923
rect 30941 13889 30975 13923
rect 30975 13889 30984 13923
rect 30932 13880 30984 13889
rect 33416 13880 33468 13932
rect 37464 14016 37516 14068
rect 36544 13991 36596 14000
rect 36544 13957 36553 13991
rect 36553 13957 36587 13991
rect 36587 13957 36596 13991
rect 36544 13948 36596 13957
rect 34796 13880 34848 13932
rect 33600 13812 33652 13864
rect 40684 13948 40736 14000
rect 36728 13923 36780 13932
rect 36728 13889 36737 13923
rect 36737 13889 36771 13923
rect 36771 13889 36780 13923
rect 38568 13923 38620 13932
rect 36728 13880 36780 13889
rect 35624 13855 35676 13864
rect 35624 13821 35633 13855
rect 35633 13821 35667 13855
rect 35667 13821 35676 13855
rect 35624 13812 35676 13821
rect 7656 13676 7708 13728
rect 13176 13719 13228 13728
rect 13176 13685 13185 13719
rect 13185 13685 13219 13719
rect 13219 13685 13228 13719
rect 13176 13676 13228 13685
rect 18696 13719 18748 13728
rect 18696 13685 18705 13719
rect 18705 13685 18739 13719
rect 18739 13685 18748 13719
rect 18696 13676 18748 13685
rect 20076 13676 20128 13728
rect 25872 13744 25924 13796
rect 29552 13787 29604 13796
rect 29552 13753 29561 13787
rect 29561 13753 29595 13787
rect 29595 13753 29604 13787
rect 29552 13744 29604 13753
rect 35992 13744 36044 13796
rect 38568 13889 38577 13923
rect 38577 13889 38611 13923
rect 38611 13889 38620 13923
rect 38568 13880 38620 13889
rect 38384 13812 38436 13864
rect 39488 13812 39540 13864
rect 40408 13812 40460 13864
rect 24952 13719 25004 13728
rect 24952 13685 24961 13719
rect 24961 13685 24995 13719
rect 24995 13685 25004 13719
rect 24952 13676 25004 13685
rect 35900 13676 35952 13728
rect 39304 13719 39356 13728
rect 39304 13685 39313 13719
rect 39313 13685 39347 13719
rect 39347 13685 39356 13719
rect 39304 13676 39356 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 14280 13515 14332 13524
rect 14280 13481 14289 13515
rect 14289 13481 14323 13515
rect 14323 13481 14332 13515
rect 14280 13472 14332 13481
rect 18788 13472 18840 13524
rect 22008 13472 22060 13524
rect 23664 13472 23716 13524
rect 27252 13515 27304 13524
rect 27252 13481 27261 13515
rect 27261 13481 27295 13515
rect 27295 13481 27304 13515
rect 27252 13472 27304 13481
rect 29092 13472 29144 13524
rect 30012 13472 30064 13524
rect 30380 13472 30432 13524
rect 35808 13472 35860 13524
rect 36544 13472 36596 13524
rect 17684 13404 17736 13456
rect 12532 13336 12584 13388
rect 19064 13336 19116 13388
rect 7748 13268 7800 13320
rect 8760 13268 8812 13320
rect 14280 13268 14332 13320
rect 9772 13200 9824 13252
rect 8300 13132 8352 13184
rect 9036 13132 9088 13184
rect 10508 13132 10560 13184
rect 14556 13132 14608 13184
rect 14832 13268 14884 13320
rect 15016 13268 15068 13320
rect 16396 13268 16448 13320
rect 21732 13404 21784 13456
rect 24768 13404 24820 13456
rect 24584 13336 24636 13388
rect 23756 13268 23808 13320
rect 27804 13336 27856 13388
rect 16672 13200 16724 13252
rect 22192 13200 22244 13252
rect 22376 13200 22428 13252
rect 25504 13243 25556 13252
rect 25504 13209 25513 13243
rect 25513 13209 25547 13243
rect 25547 13209 25556 13243
rect 25504 13200 25556 13209
rect 14740 13132 14792 13184
rect 15108 13132 15160 13184
rect 18512 13132 18564 13184
rect 18972 13132 19024 13184
rect 21364 13132 21416 13184
rect 26792 13175 26844 13184
rect 26792 13141 26801 13175
rect 26801 13141 26835 13175
rect 26835 13141 26844 13175
rect 26792 13132 26844 13141
rect 27712 13311 27764 13320
rect 27712 13277 27721 13311
rect 27721 13277 27755 13311
rect 27755 13277 27764 13311
rect 28264 13336 28316 13388
rect 30564 13336 30616 13388
rect 27712 13268 27764 13277
rect 29736 13268 29788 13320
rect 30012 13311 30064 13320
rect 30012 13277 30021 13311
rect 30021 13277 30055 13311
rect 30055 13277 30064 13311
rect 30012 13268 30064 13277
rect 30656 13268 30708 13320
rect 31208 13268 31260 13320
rect 38384 13404 38436 13456
rect 34428 13268 34480 13320
rect 38108 13268 38160 13320
rect 32312 13200 32364 13252
rect 33324 13200 33376 13252
rect 35440 13200 35492 13252
rect 37096 13200 37148 13252
rect 38568 13311 38620 13320
rect 38568 13277 38577 13311
rect 38577 13277 38611 13311
rect 38611 13277 38620 13311
rect 38568 13268 38620 13277
rect 58164 13311 58216 13320
rect 58164 13277 58173 13311
rect 58173 13277 58207 13311
rect 58207 13277 58216 13311
rect 58164 13268 58216 13277
rect 29920 13132 29972 13184
rect 32588 13132 32640 13184
rect 37280 13132 37332 13184
rect 39304 13200 39356 13252
rect 38844 13175 38896 13184
rect 38844 13141 38853 13175
rect 38853 13141 38887 13175
rect 38887 13141 38896 13175
rect 38844 13132 38896 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 7656 12928 7708 12980
rect 11060 12860 11112 12912
rect 14832 12928 14884 12980
rect 15752 12928 15804 12980
rect 16028 12928 16080 12980
rect 18788 12928 18840 12980
rect 21088 12928 21140 12980
rect 23480 12928 23532 12980
rect 23756 12928 23808 12980
rect 29736 12971 29788 12980
rect 29736 12937 29745 12971
rect 29745 12937 29779 12971
rect 29779 12937 29788 12971
rect 29736 12928 29788 12937
rect 30656 12971 30708 12980
rect 30656 12937 30665 12971
rect 30665 12937 30699 12971
rect 30699 12937 30708 12971
rect 30656 12928 30708 12937
rect 30840 12928 30892 12980
rect 32312 12928 32364 12980
rect 33324 12971 33376 12980
rect 33324 12937 33333 12971
rect 33333 12937 33367 12971
rect 33367 12937 33376 12971
rect 33324 12928 33376 12937
rect 35440 12971 35492 12980
rect 35440 12937 35449 12971
rect 35449 12937 35483 12971
rect 35483 12937 35492 12971
rect 35440 12928 35492 12937
rect 35532 12928 35584 12980
rect 37280 12928 37332 12980
rect 5356 12835 5408 12844
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 7840 12792 7892 12844
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 16856 12860 16908 12912
rect 2688 12767 2740 12776
rect 2688 12733 2697 12767
rect 2697 12733 2731 12767
rect 2731 12733 2740 12767
rect 2688 12724 2740 12733
rect 2872 12724 2924 12776
rect 4620 12724 4672 12776
rect 5448 12767 5500 12776
rect 5448 12733 5457 12767
rect 5457 12733 5491 12767
rect 5491 12733 5500 12767
rect 5448 12724 5500 12733
rect 6828 12767 6880 12776
rect 4712 12656 4764 12708
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 6000 12656 6052 12708
rect 9680 12724 9732 12776
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 13176 12792 13228 12844
rect 15108 12835 15160 12844
rect 15108 12801 15117 12835
rect 15117 12801 15151 12835
rect 15151 12801 15160 12835
rect 15108 12792 15160 12801
rect 18052 12835 18104 12844
rect 18972 12860 19024 12912
rect 18052 12801 18070 12835
rect 18070 12801 18104 12835
rect 18052 12792 18104 12801
rect 18696 12792 18748 12844
rect 11980 12724 12032 12733
rect 16672 12724 16724 12776
rect 18788 12724 18840 12776
rect 19248 12835 19300 12844
rect 19248 12801 19257 12835
rect 19257 12801 19291 12835
rect 19291 12801 19300 12835
rect 20628 12860 20680 12912
rect 20812 12860 20864 12912
rect 26148 12903 26200 12912
rect 26148 12869 26157 12903
rect 26157 12869 26191 12903
rect 26191 12869 26200 12903
rect 26148 12860 26200 12869
rect 29368 12903 29420 12912
rect 29368 12869 29377 12903
rect 29377 12869 29411 12903
rect 29411 12869 29420 12903
rect 29368 12860 29420 12869
rect 29552 12903 29604 12912
rect 29552 12869 29561 12903
rect 29561 12869 29595 12903
rect 29595 12869 29604 12903
rect 29552 12860 29604 12869
rect 19248 12792 19300 12801
rect 20076 12792 20128 12844
rect 21180 12792 21232 12844
rect 21456 12792 21508 12844
rect 26240 12792 26292 12844
rect 27068 12792 27120 12844
rect 32680 12835 32732 12844
rect 32680 12801 32689 12835
rect 32689 12801 32723 12835
rect 32723 12801 32732 12835
rect 32680 12792 32732 12801
rect 32864 12835 32916 12844
rect 32864 12801 32873 12835
rect 32873 12801 32907 12835
rect 32907 12801 32916 12835
rect 32864 12792 32916 12801
rect 32956 12835 33008 12844
rect 32956 12801 32965 12835
rect 32965 12801 32999 12835
rect 32999 12801 33008 12835
rect 32956 12792 33008 12801
rect 35624 12860 35676 12912
rect 2136 12588 2188 12640
rect 6368 12631 6420 12640
rect 6368 12597 6377 12631
rect 6377 12597 6411 12631
rect 6411 12597 6420 12631
rect 6368 12588 6420 12597
rect 8300 12631 8352 12640
rect 8300 12597 8309 12631
rect 8309 12597 8343 12631
rect 8343 12597 8352 12631
rect 8300 12588 8352 12597
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 15108 12588 15160 12640
rect 16396 12656 16448 12708
rect 21640 12724 21692 12776
rect 22192 12724 22244 12776
rect 27344 12724 27396 12776
rect 34336 12767 34388 12776
rect 18420 12588 18472 12640
rect 21916 12588 21968 12640
rect 25504 12588 25556 12640
rect 33232 12588 33284 12640
rect 33876 12588 33928 12640
rect 34336 12733 34345 12767
rect 34345 12733 34379 12767
rect 34379 12733 34388 12767
rect 34336 12724 34388 12733
rect 35624 12724 35676 12776
rect 35900 12835 35952 12844
rect 35900 12801 35909 12835
rect 35909 12801 35943 12835
rect 35943 12801 35952 12835
rect 38844 12860 38896 12912
rect 35900 12792 35952 12801
rect 37648 12835 37700 12844
rect 37648 12801 37657 12835
rect 37657 12801 37691 12835
rect 37691 12801 37700 12835
rect 37648 12792 37700 12801
rect 38108 12792 38160 12844
rect 35992 12724 36044 12776
rect 39580 12792 39632 12844
rect 36452 12588 36504 12640
rect 37096 12588 37148 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 6368 12384 6420 12436
rect 9772 12384 9824 12436
rect 6276 12316 6328 12368
rect 12532 12384 12584 12436
rect 14096 12384 14148 12436
rect 22376 12384 22428 12436
rect 3792 12291 3844 12300
rect 3792 12257 3801 12291
rect 3801 12257 3835 12291
rect 3835 12257 3844 12291
rect 3792 12248 3844 12257
rect 5356 12248 5408 12300
rect 7380 12248 7432 12300
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 6184 12180 6236 12232
rect 6460 12180 6512 12232
rect 7012 12180 7064 12232
rect 13820 12316 13872 12368
rect 15016 12316 15068 12368
rect 4620 12112 4672 12164
rect 5540 12044 5592 12096
rect 6552 12044 6604 12096
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 7656 12112 7708 12164
rect 10692 12180 10744 12232
rect 11520 12180 11572 12232
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 15200 12248 15252 12300
rect 16672 12316 16724 12368
rect 20168 12316 20220 12368
rect 9772 12112 9824 12164
rect 12072 12112 12124 12164
rect 12348 12112 12400 12164
rect 14556 12112 14608 12164
rect 15108 12223 15160 12232
rect 15108 12189 15117 12223
rect 15117 12189 15151 12223
rect 15151 12189 15160 12223
rect 16120 12248 16172 12300
rect 17132 12248 17184 12300
rect 20996 12291 21048 12300
rect 15108 12180 15160 12189
rect 10600 12044 10652 12096
rect 11704 12044 11756 12096
rect 13268 12044 13320 12096
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 14648 12087 14700 12096
rect 14648 12053 14657 12087
rect 14657 12053 14691 12087
rect 14691 12053 14700 12087
rect 14648 12044 14700 12053
rect 15200 12112 15252 12164
rect 16028 12180 16080 12232
rect 18144 12180 18196 12232
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 19064 12180 19116 12232
rect 19340 12180 19392 12232
rect 20996 12257 21005 12291
rect 21005 12257 21039 12291
rect 21039 12257 21048 12291
rect 20996 12248 21048 12257
rect 21456 12291 21508 12300
rect 21456 12257 21465 12291
rect 21465 12257 21499 12291
rect 21499 12257 21508 12291
rect 21456 12248 21508 12257
rect 15752 12112 15804 12164
rect 16580 12112 16632 12164
rect 18052 12155 18104 12164
rect 16856 12044 16908 12096
rect 18052 12121 18061 12155
rect 18061 12121 18095 12155
rect 18095 12121 18104 12155
rect 18052 12112 18104 12121
rect 18788 12112 18840 12164
rect 22008 12316 22060 12368
rect 22560 12316 22612 12368
rect 20168 12112 20220 12164
rect 21916 12223 21968 12232
rect 21916 12189 21930 12223
rect 21930 12189 21964 12223
rect 21964 12189 21968 12223
rect 21916 12180 21968 12189
rect 22100 12223 22152 12232
rect 22100 12189 22109 12223
rect 22109 12189 22143 12223
rect 22143 12189 22152 12223
rect 27896 12384 27948 12436
rect 32864 12427 32916 12436
rect 32864 12393 32873 12427
rect 32873 12393 32907 12427
rect 32907 12393 32916 12427
rect 32864 12384 32916 12393
rect 33876 12427 33928 12436
rect 33876 12393 33885 12427
rect 33885 12393 33919 12427
rect 33919 12393 33928 12427
rect 33876 12384 33928 12393
rect 35624 12384 35676 12436
rect 37004 12316 37056 12368
rect 38568 12316 38620 12368
rect 30104 12291 30156 12300
rect 30104 12257 30113 12291
rect 30113 12257 30147 12291
rect 30147 12257 30156 12291
rect 30104 12248 30156 12257
rect 25044 12223 25096 12232
rect 22100 12180 22152 12189
rect 25044 12189 25053 12223
rect 25053 12189 25087 12223
rect 25087 12189 25096 12223
rect 25044 12180 25096 12189
rect 26148 12180 26200 12232
rect 22192 12112 22244 12164
rect 25136 12112 25188 12164
rect 28080 12180 28132 12232
rect 30564 12223 30616 12232
rect 30564 12189 30573 12223
rect 30573 12189 30607 12223
rect 30607 12189 30616 12223
rect 30564 12180 30616 12189
rect 30748 12223 30800 12232
rect 30748 12189 30757 12223
rect 30757 12189 30791 12223
rect 30791 12189 30800 12223
rect 30748 12180 30800 12189
rect 31024 12248 31076 12300
rect 39028 12248 39080 12300
rect 19064 12044 19116 12096
rect 28172 12155 28224 12164
rect 28172 12121 28181 12155
rect 28181 12121 28215 12155
rect 28215 12121 28224 12155
rect 28172 12112 28224 12121
rect 31208 12180 31260 12232
rect 32956 12180 33008 12232
rect 34336 12180 34388 12232
rect 38292 12223 38344 12232
rect 38292 12189 38301 12223
rect 38301 12189 38335 12223
rect 38335 12189 38344 12223
rect 38292 12180 38344 12189
rect 39488 12180 39540 12232
rect 39764 12180 39816 12232
rect 26056 12044 26108 12096
rect 27436 12087 27488 12096
rect 27436 12053 27445 12087
rect 27445 12053 27479 12087
rect 27479 12053 27488 12087
rect 27436 12044 27488 12053
rect 30196 12044 30248 12096
rect 32588 12112 32640 12164
rect 31392 12044 31444 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 7656 11840 7708 11892
rect 14740 11840 14792 11892
rect 17132 11883 17184 11892
rect 17132 11849 17141 11883
rect 17141 11849 17175 11883
rect 17175 11849 17184 11883
rect 17132 11840 17184 11849
rect 17316 11840 17368 11892
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 3792 11772 3844 11824
rect 6184 11772 6236 11824
rect 5540 11747 5592 11756
rect 5540 11713 5549 11747
rect 5549 11713 5583 11747
rect 5583 11713 5592 11747
rect 5540 11704 5592 11713
rect 5264 11636 5316 11688
rect 6460 11636 6512 11688
rect 7104 11772 7156 11824
rect 12532 11772 12584 11824
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 13268 11747 13320 11756
rect 13268 11713 13277 11747
rect 13277 11713 13311 11747
rect 13311 11713 13320 11747
rect 13268 11704 13320 11713
rect 7104 11636 7156 11688
rect 12348 11679 12400 11688
rect 12348 11645 12357 11679
rect 12357 11645 12391 11679
rect 12391 11645 12400 11679
rect 12348 11636 12400 11645
rect 13452 11747 13504 11756
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 13820 11704 13872 11756
rect 14648 11704 14700 11756
rect 16856 11772 16908 11824
rect 20812 11840 20864 11892
rect 23848 11840 23900 11892
rect 24492 11840 24544 11892
rect 25136 11883 25188 11892
rect 18420 11704 18472 11756
rect 21456 11772 21508 11824
rect 23480 11772 23532 11824
rect 25136 11849 25145 11883
rect 25145 11849 25179 11883
rect 25179 11849 25188 11883
rect 25136 11840 25188 11849
rect 27896 11840 27948 11892
rect 30748 11840 30800 11892
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 14464 11636 14516 11688
rect 6736 11568 6788 11620
rect 7012 11568 7064 11620
rect 10876 11568 10928 11620
rect 22008 11704 22060 11756
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 21640 11636 21692 11688
rect 22376 11747 22428 11756
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 26148 11772 26200 11824
rect 22560 11704 22612 11713
rect 25596 11747 25648 11756
rect 25596 11713 25605 11747
rect 25605 11713 25639 11747
rect 25639 11713 25648 11747
rect 25596 11704 25648 11713
rect 27436 11704 27488 11756
rect 28172 11772 28224 11824
rect 30288 11747 30340 11756
rect 30288 11713 30297 11747
rect 30297 11713 30331 11747
rect 30331 11713 30340 11747
rect 30288 11704 30340 11713
rect 30564 11704 30616 11756
rect 31116 11747 31168 11756
rect 30196 11636 30248 11688
rect 31116 11713 31125 11747
rect 31125 11713 31159 11747
rect 31159 11713 31168 11747
rect 31116 11704 31168 11713
rect 31208 11747 31260 11756
rect 31208 11713 31217 11747
rect 31217 11713 31251 11747
rect 31251 11713 31260 11747
rect 31208 11704 31260 11713
rect 31484 11704 31536 11756
rect 31944 11704 31996 11756
rect 34428 11840 34480 11892
rect 39856 11840 39908 11892
rect 36636 11772 36688 11824
rect 38292 11772 38344 11824
rect 34336 11704 34388 11756
rect 34796 11704 34848 11756
rect 35808 11747 35860 11756
rect 32128 11636 32180 11688
rect 32680 11679 32732 11688
rect 32680 11645 32689 11679
rect 32689 11645 32723 11679
rect 32723 11645 32732 11679
rect 32680 11636 32732 11645
rect 35808 11713 35817 11747
rect 35817 11713 35851 11747
rect 35851 11713 35860 11747
rect 35808 11704 35860 11713
rect 38660 11704 38712 11756
rect 35716 11636 35768 11688
rect 38568 11679 38620 11688
rect 38568 11645 38577 11679
rect 38577 11645 38611 11679
rect 38611 11645 38620 11679
rect 38568 11636 38620 11645
rect 4896 11500 4948 11552
rect 5448 11500 5500 11552
rect 12992 11543 13044 11552
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 12992 11500 13044 11509
rect 15476 11500 15528 11552
rect 16028 11543 16080 11552
rect 16028 11509 16037 11543
rect 16037 11509 16071 11543
rect 16071 11509 16080 11543
rect 16028 11500 16080 11509
rect 16120 11500 16172 11552
rect 18696 11500 18748 11552
rect 21916 11543 21968 11552
rect 21916 11509 21925 11543
rect 21925 11509 21959 11543
rect 21959 11509 21968 11543
rect 21916 11500 21968 11509
rect 24492 11568 24544 11620
rect 27896 11568 27948 11620
rect 31668 11568 31720 11620
rect 35440 11568 35492 11620
rect 58164 11611 58216 11620
rect 58164 11577 58173 11611
rect 58173 11577 58207 11611
rect 58207 11577 58216 11611
rect 58164 11568 58216 11577
rect 24124 11543 24176 11552
rect 24124 11509 24133 11543
rect 24133 11509 24167 11543
rect 24167 11509 24176 11543
rect 24124 11500 24176 11509
rect 33048 11500 33100 11552
rect 40776 11543 40828 11552
rect 40776 11509 40785 11543
rect 40785 11509 40819 11543
rect 40819 11509 40828 11543
rect 40776 11500 40828 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 13452 11296 13504 11348
rect 18144 11296 18196 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 19064 11296 19116 11348
rect 20168 11339 20220 11348
rect 20168 11305 20177 11339
rect 20177 11305 20211 11339
rect 20211 11305 20220 11339
rect 20168 11296 20220 11305
rect 21640 11296 21692 11348
rect 25044 11296 25096 11348
rect 25596 11296 25648 11348
rect 30288 11296 30340 11348
rect 33416 11296 33468 11348
rect 37004 11296 37056 11348
rect 38108 11339 38160 11348
rect 38108 11305 38117 11339
rect 38117 11305 38151 11339
rect 38151 11305 38160 11339
rect 38108 11296 38160 11305
rect 38660 11339 38712 11348
rect 38660 11305 38669 11339
rect 38669 11305 38703 11339
rect 38703 11305 38712 11339
rect 38660 11296 38712 11305
rect 15476 11271 15528 11280
rect 15476 11237 15485 11271
rect 15485 11237 15519 11271
rect 15519 11237 15528 11271
rect 15476 11228 15528 11237
rect 21364 11228 21416 11280
rect 29092 11228 29144 11280
rect 29368 11228 29420 11280
rect 5632 11160 5684 11212
rect 6552 11160 6604 11212
rect 12532 11160 12584 11212
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 9772 11092 9824 11144
rect 12992 11092 13044 11144
rect 21640 11203 21692 11212
rect 21640 11169 21649 11203
rect 21649 11169 21683 11203
rect 21683 11169 21692 11203
rect 21640 11160 21692 11169
rect 23848 11203 23900 11212
rect 23848 11169 23857 11203
rect 23857 11169 23891 11203
rect 23891 11169 23900 11203
rect 23848 11160 23900 11169
rect 24124 11160 24176 11212
rect 16672 11092 16724 11144
rect 21088 11092 21140 11144
rect 21916 11135 21968 11144
rect 21916 11101 21950 11135
rect 21950 11101 21968 11135
rect 21916 11092 21968 11101
rect 23020 11092 23072 11144
rect 24584 11092 24636 11144
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 31024 11160 31076 11212
rect 26056 11135 26108 11144
rect 10140 11067 10192 11076
rect 10140 11033 10149 11067
rect 10149 11033 10183 11067
rect 10183 11033 10192 11067
rect 10140 11024 10192 11033
rect 11336 11024 11388 11076
rect 12716 11024 12768 11076
rect 14188 11024 14240 11076
rect 14924 11024 14976 11076
rect 20996 11067 21048 11076
rect 20996 11033 21005 11067
rect 21005 11033 21039 11067
rect 21039 11033 21048 11067
rect 20996 11024 21048 11033
rect 24860 11024 24912 11076
rect 26056 11101 26065 11135
rect 26065 11101 26099 11135
rect 26099 11101 26108 11135
rect 26056 11092 26108 11101
rect 26148 11092 26200 11144
rect 28448 11092 28500 11144
rect 29092 11092 29144 11144
rect 30932 11092 30984 11144
rect 35624 11135 35676 11144
rect 35624 11101 35633 11135
rect 35633 11101 35667 11135
rect 35667 11101 35676 11135
rect 35624 11092 35676 11101
rect 39028 11228 39080 11280
rect 36636 11135 36688 11144
rect 26240 11067 26292 11076
rect 26240 11033 26249 11067
rect 26249 11033 26283 11067
rect 26283 11033 26292 11067
rect 26240 11024 26292 11033
rect 28632 11024 28684 11076
rect 31392 11067 31444 11076
rect 31392 11033 31426 11067
rect 31426 11033 31444 11067
rect 31392 11024 31444 11033
rect 9680 10956 9732 11008
rect 11888 10956 11940 11008
rect 15016 10956 15068 11008
rect 15660 10956 15712 11008
rect 16488 10956 16540 11008
rect 19432 10956 19484 11008
rect 22468 10956 22520 11008
rect 23480 10999 23532 11008
rect 23480 10965 23489 10999
rect 23489 10965 23523 10999
rect 23523 10965 23532 10999
rect 23480 10956 23532 10965
rect 24676 10956 24728 11008
rect 25412 10999 25464 11008
rect 25412 10965 25421 10999
rect 25421 10965 25455 10999
rect 25455 10965 25464 10999
rect 25412 10956 25464 10965
rect 31484 10956 31536 11008
rect 31668 10956 31720 11008
rect 36636 11101 36645 11135
rect 36645 11101 36679 11135
rect 36679 11101 36688 11135
rect 36636 11092 36688 11101
rect 38476 11092 38528 11144
rect 40776 11160 40828 11212
rect 37556 11024 37608 11076
rect 38292 11024 38344 11076
rect 35348 10999 35400 11008
rect 35348 10965 35357 10999
rect 35357 10965 35391 10999
rect 35391 10965 35400 10999
rect 35348 10956 35400 10965
rect 38108 10956 38160 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 6276 10752 6328 10804
rect 11980 10752 12032 10804
rect 15016 10752 15068 10804
rect 17592 10752 17644 10804
rect 22376 10752 22428 10804
rect 23664 10752 23716 10804
rect 4620 10616 4672 10668
rect 9220 10684 9272 10736
rect 12624 10684 12676 10736
rect 17316 10727 17368 10736
rect 17316 10693 17325 10727
rect 17325 10693 17359 10727
rect 17359 10693 17368 10727
rect 17316 10684 17368 10693
rect 23480 10684 23532 10736
rect 6552 10659 6604 10668
rect 6552 10625 6561 10659
rect 6561 10625 6595 10659
rect 6595 10625 6604 10659
rect 6552 10616 6604 10625
rect 7288 10616 7340 10668
rect 9956 10616 10008 10668
rect 10140 10616 10192 10668
rect 10416 10616 10468 10668
rect 17132 10659 17184 10668
rect 17132 10625 17141 10659
rect 17141 10625 17175 10659
rect 17175 10625 17184 10659
rect 17132 10616 17184 10625
rect 22468 10616 22520 10668
rect 23020 10659 23072 10668
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 4896 10548 4948 10600
rect 5632 10523 5684 10532
rect 5632 10489 5641 10523
rect 5641 10489 5675 10523
rect 5675 10489 5684 10523
rect 5632 10480 5684 10489
rect 6000 10480 6052 10532
rect 9680 10548 9732 10600
rect 10876 10548 10928 10600
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 11980 10591 12032 10600
rect 11980 10557 11989 10591
rect 11989 10557 12023 10591
rect 12023 10557 12032 10591
rect 11980 10548 12032 10557
rect 21364 10548 21416 10600
rect 22836 10548 22888 10600
rect 23296 10616 23348 10668
rect 24768 10684 24820 10736
rect 25412 10684 25464 10736
rect 31116 10752 31168 10804
rect 36636 10795 36688 10804
rect 36636 10761 36645 10795
rect 36645 10761 36679 10795
rect 36679 10761 36688 10795
rect 36636 10752 36688 10761
rect 38108 10752 38160 10804
rect 33048 10684 33100 10736
rect 24216 10616 24268 10668
rect 24860 10616 24912 10668
rect 25044 10659 25096 10668
rect 25044 10625 25053 10659
rect 25053 10625 25087 10659
rect 25087 10625 25096 10659
rect 25044 10616 25096 10625
rect 24492 10548 24544 10600
rect 24676 10548 24728 10600
rect 26240 10616 26292 10668
rect 30288 10616 30340 10668
rect 31944 10616 31996 10668
rect 34704 10548 34756 10600
rect 38568 10684 38620 10736
rect 35348 10616 35400 10668
rect 37740 10616 37792 10668
rect 39028 10548 39080 10600
rect 39396 10659 39448 10668
rect 39396 10625 39405 10659
rect 39405 10625 39439 10659
rect 39439 10625 39448 10659
rect 39396 10616 39448 10625
rect 14096 10480 14148 10532
rect 27068 10480 27120 10532
rect 30380 10480 30432 10532
rect 9220 10455 9272 10464
rect 9220 10421 9229 10455
rect 9229 10421 9263 10455
rect 9263 10421 9272 10455
rect 9220 10412 9272 10421
rect 18144 10412 18196 10464
rect 19248 10412 19300 10464
rect 20996 10412 21048 10464
rect 21640 10412 21692 10464
rect 25412 10412 25464 10464
rect 27988 10412 28040 10464
rect 29552 10412 29604 10464
rect 29920 10455 29972 10464
rect 29920 10421 29929 10455
rect 29929 10421 29963 10455
rect 29963 10421 29972 10455
rect 29920 10412 29972 10421
rect 31944 10412 31996 10464
rect 32404 10412 32456 10464
rect 34520 10412 34572 10464
rect 35624 10412 35676 10464
rect 38936 10455 38988 10464
rect 38936 10421 38945 10455
rect 38945 10421 38979 10455
rect 38979 10421 38988 10455
rect 38936 10412 38988 10421
rect 58164 10455 58216 10464
rect 58164 10421 58173 10455
rect 58173 10421 58207 10455
rect 58207 10421 58216 10455
rect 58164 10412 58216 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 16488 10251 16540 10260
rect 16488 10217 16497 10251
rect 16497 10217 16531 10251
rect 16531 10217 16540 10251
rect 16488 10208 16540 10217
rect 22836 10251 22888 10260
rect 22836 10217 22845 10251
rect 22845 10217 22879 10251
rect 22879 10217 22888 10251
rect 22836 10208 22888 10217
rect 24952 10208 25004 10260
rect 28540 10208 28592 10260
rect 29276 10208 29328 10260
rect 38568 10251 38620 10260
rect 38568 10217 38577 10251
rect 38577 10217 38611 10251
rect 38611 10217 38620 10251
rect 38568 10208 38620 10217
rect 8208 10140 8260 10192
rect 24308 10140 24360 10192
rect 30380 10140 30432 10192
rect 5632 10115 5684 10124
rect 5632 10081 5641 10115
rect 5641 10081 5675 10115
rect 5675 10081 5684 10115
rect 10416 10115 10468 10124
rect 5632 10072 5684 10081
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 6184 10004 6236 10056
rect 8944 10047 8996 10056
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 10416 10081 10425 10115
rect 10425 10081 10459 10115
rect 10459 10081 10468 10115
rect 10416 10072 10468 10081
rect 13544 10072 13596 10124
rect 24492 10072 24544 10124
rect 26608 10072 26660 10124
rect 28632 10072 28684 10124
rect 24676 10004 24728 10056
rect 25412 10047 25464 10056
rect 25412 10013 25421 10047
rect 25421 10013 25455 10047
rect 25455 10013 25464 10047
rect 25412 10004 25464 10013
rect 27712 10047 27764 10056
rect 27712 10013 27721 10047
rect 27721 10013 27755 10047
rect 27755 10013 27764 10047
rect 27712 10004 27764 10013
rect 27988 10047 28040 10056
rect 27988 10013 27997 10047
rect 27997 10013 28031 10047
rect 28031 10013 28040 10047
rect 27988 10004 28040 10013
rect 28540 10004 28592 10056
rect 29276 10004 29328 10056
rect 31208 10072 31260 10124
rect 30012 10047 30064 10056
rect 30012 10013 30021 10047
rect 30021 10013 30055 10047
rect 30055 10013 30064 10047
rect 30012 10004 30064 10013
rect 32128 10004 32180 10056
rect 37188 10004 37240 10056
rect 6460 9979 6512 9988
rect 1676 9868 1728 9920
rect 5448 9911 5500 9920
rect 5448 9877 5457 9911
rect 5457 9877 5491 9911
rect 5491 9877 5500 9911
rect 6460 9945 6469 9979
rect 6469 9945 6503 9979
rect 6503 9945 6512 9979
rect 6460 9936 6512 9945
rect 11980 9936 12032 9988
rect 14096 9936 14148 9988
rect 17132 9936 17184 9988
rect 5448 9868 5500 9877
rect 6368 9868 6420 9920
rect 6828 9868 6880 9920
rect 8392 9868 8444 9920
rect 9128 9911 9180 9920
rect 9128 9877 9137 9911
rect 9137 9877 9171 9911
rect 9171 9877 9180 9911
rect 9128 9868 9180 9877
rect 10324 9911 10376 9920
rect 10324 9877 10333 9911
rect 10333 9877 10367 9911
rect 10367 9877 10376 9911
rect 10324 9868 10376 9877
rect 24676 9868 24728 9920
rect 28448 9936 28500 9988
rect 30656 9868 30708 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 8944 9664 8996 9716
rect 10416 9664 10468 9716
rect 19984 9664 20036 9716
rect 21364 9664 21416 9716
rect 22468 9664 22520 9716
rect 5540 9596 5592 9648
rect 7288 9639 7340 9648
rect 7288 9605 7297 9639
rect 7297 9605 7331 9639
rect 7331 9605 7340 9639
rect 7288 9596 7340 9605
rect 9128 9639 9180 9648
rect 9128 9605 9162 9639
rect 9162 9605 9180 9639
rect 9128 9596 9180 9605
rect 9588 9596 9640 9648
rect 16764 9596 16816 9648
rect 20720 9639 20772 9648
rect 20720 9605 20729 9639
rect 20729 9605 20763 9639
rect 20763 9605 20772 9639
rect 20720 9596 20772 9605
rect 26056 9596 26108 9648
rect 30012 9664 30064 9716
rect 28172 9596 28224 9648
rect 29552 9639 29604 9648
rect 29552 9605 29561 9639
rect 29561 9605 29595 9639
rect 29595 9605 29604 9639
rect 29552 9596 29604 9605
rect 30288 9596 30340 9648
rect 35808 9596 35860 9648
rect 36360 9596 36412 9648
rect 37556 9639 37608 9648
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 1860 9460 1912 9512
rect 5448 9528 5500 9580
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 12532 9528 12584 9580
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 14280 9528 14332 9580
rect 14464 9528 14516 9580
rect 17868 9528 17920 9580
rect 18696 9528 18748 9580
rect 22652 9571 22704 9580
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 5632 9460 5684 9512
rect 6460 9460 6512 9512
rect 8852 9503 8904 9512
rect 8852 9469 8861 9503
rect 8861 9469 8895 9503
rect 8895 9469 8904 9503
rect 8852 9460 8904 9469
rect 13544 9503 13596 9512
rect 13544 9469 13553 9503
rect 13553 9469 13587 9503
rect 13587 9469 13596 9503
rect 13544 9460 13596 9469
rect 22192 9460 22244 9512
rect 22928 9528 22980 9580
rect 25412 9571 25464 9580
rect 25412 9537 25421 9571
rect 25421 9537 25455 9571
rect 25455 9537 25464 9571
rect 25412 9528 25464 9537
rect 29736 9571 29788 9580
rect 29736 9537 29745 9571
rect 29745 9537 29779 9571
rect 29779 9537 29788 9571
rect 29736 9528 29788 9537
rect 32128 9571 32180 9580
rect 32128 9537 32137 9571
rect 32137 9537 32171 9571
rect 32171 9537 32180 9571
rect 32128 9528 32180 9537
rect 32312 9571 32364 9580
rect 32312 9537 32321 9571
rect 32321 9537 32355 9571
rect 32355 9537 32364 9571
rect 32312 9528 32364 9537
rect 28540 9503 28592 9512
rect 3976 9324 4028 9376
rect 6276 9324 6328 9376
rect 6368 9324 6420 9376
rect 6920 9324 6972 9376
rect 7380 9367 7432 9376
rect 7380 9333 7389 9367
rect 7389 9333 7423 9367
rect 7423 9333 7432 9367
rect 7380 9324 7432 9333
rect 13912 9392 13964 9444
rect 23388 9392 23440 9444
rect 26700 9392 26752 9444
rect 28540 9469 28549 9503
rect 28549 9469 28583 9503
rect 28583 9469 28592 9503
rect 28540 9460 28592 9469
rect 29920 9460 29972 9512
rect 32496 9571 32548 9580
rect 32496 9537 32505 9571
rect 32505 9537 32539 9571
rect 32539 9537 32548 9571
rect 32496 9528 32548 9537
rect 36452 9528 36504 9580
rect 37556 9605 37565 9639
rect 37565 9605 37599 9639
rect 37599 9605 37608 9639
rect 37556 9596 37608 9605
rect 39396 9664 39448 9716
rect 38936 9596 38988 9648
rect 32956 9460 33008 9512
rect 37924 9460 37976 9512
rect 28724 9392 28776 9444
rect 10324 9324 10376 9376
rect 10416 9324 10468 9376
rect 12532 9367 12584 9376
rect 12532 9333 12541 9367
rect 12541 9333 12575 9367
rect 12575 9333 12584 9367
rect 12532 9324 12584 9333
rect 13176 9324 13228 9376
rect 14372 9367 14424 9376
rect 14372 9333 14381 9367
rect 14381 9333 14415 9367
rect 14415 9333 14424 9367
rect 14372 9324 14424 9333
rect 15568 9324 15620 9376
rect 15936 9324 15988 9376
rect 17224 9324 17276 9376
rect 17868 9367 17920 9376
rect 17868 9333 17877 9367
rect 17877 9333 17911 9367
rect 17911 9333 17920 9367
rect 17868 9324 17920 9333
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 33600 9324 33652 9376
rect 35348 9324 35400 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 6644 9120 6696 9172
rect 10232 9163 10284 9172
rect 4712 9095 4764 9104
rect 4712 9061 4721 9095
rect 4721 9061 4755 9095
rect 4755 9061 4764 9095
rect 4712 9052 4764 9061
rect 2872 8984 2924 9036
rect 3976 8984 4028 9036
rect 5264 8984 5316 9036
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 4988 8916 5040 8968
rect 7012 8916 7064 8968
rect 9864 9052 9916 9104
rect 4620 8848 4672 8900
rect 6276 8848 6328 8900
rect 9772 8984 9824 9036
rect 10232 9129 10241 9163
rect 10241 9129 10275 9163
rect 10275 9129 10284 9163
rect 20628 9163 20680 9172
rect 10232 9120 10284 9129
rect 10324 9052 10376 9104
rect 11244 8984 11296 9036
rect 9496 8959 9548 8968
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 9496 8916 9548 8925
rect 9864 8916 9916 8968
rect 11888 8984 11940 9036
rect 14188 9052 14240 9104
rect 16120 9095 16172 9104
rect 16120 9061 16129 9095
rect 16129 9061 16163 9095
rect 16163 9061 16172 9095
rect 16120 9052 16172 9061
rect 17040 9052 17092 9104
rect 18696 9095 18748 9104
rect 18696 9061 18705 9095
rect 18705 9061 18739 9095
rect 18739 9061 18748 9095
rect 18696 9052 18748 9061
rect 20628 9129 20637 9163
rect 20637 9129 20671 9163
rect 20671 9129 20680 9163
rect 20628 9120 20680 9129
rect 25412 9120 25464 9172
rect 30472 9120 30524 9172
rect 31852 9120 31904 9172
rect 33692 9163 33744 9172
rect 33692 9129 33701 9163
rect 33701 9129 33735 9163
rect 33735 9129 33744 9163
rect 33692 9120 33744 9129
rect 35808 9120 35860 9172
rect 22560 9052 22612 9104
rect 28540 9052 28592 9104
rect 16856 8984 16908 9036
rect 21824 8984 21876 9036
rect 22192 9027 22244 9036
rect 22192 8993 22201 9027
rect 22201 8993 22235 9027
rect 22235 8993 22244 9027
rect 22192 8984 22244 8993
rect 34704 9027 34756 9036
rect 13176 8959 13228 8968
rect 10232 8848 10284 8900
rect 11244 8848 11296 8900
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 1676 8780 1728 8832
rect 2780 8780 2832 8832
rect 3884 8823 3936 8832
rect 3884 8789 3893 8823
rect 3893 8789 3927 8823
rect 3927 8789 3936 8823
rect 3884 8780 3936 8789
rect 6552 8780 6604 8832
rect 8116 8780 8168 8832
rect 9680 8823 9732 8832
rect 9680 8789 9689 8823
rect 9689 8789 9723 8823
rect 9723 8789 9732 8823
rect 9680 8780 9732 8789
rect 9772 8780 9824 8832
rect 13176 8925 13185 8959
rect 13185 8925 13219 8959
rect 13219 8925 13228 8959
rect 13176 8916 13228 8925
rect 14372 8916 14424 8968
rect 15936 8959 15988 8968
rect 15936 8925 15945 8959
rect 15945 8925 15979 8959
rect 15979 8925 15988 8959
rect 15936 8916 15988 8925
rect 13452 8848 13504 8900
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 13912 8780 13964 8832
rect 14188 8780 14240 8832
rect 14464 8780 14516 8832
rect 18972 8916 19024 8968
rect 19064 8916 19116 8968
rect 20720 8916 20772 8968
rect 28356 8959 28408 8968
rect 28356 8925 28365 8959
rect 28365 8925 28399 8959
rect 28399 8925 28408 8959
rect 28356 8916 28408 8925
rect 28724 8959 28776 8968
rect 28724 8925 28733 8959
rect 28733 8925 28767 8959
rect 28767 8925 28776 8959
rect 28724 8916 28776 8925
rect 31300 8916 31352 8968
rect 32404 8959 32456 8968
rect 32404 8925 32413 8959
rect 32413 8925 32447 8959
rect 32447 8925 32456 8959
rect 32404 8916 32456 8925
rect 32680 8916 32732 8968
rect 33140 8959 33192 8968
rect 33140 8925 33149 8959
rect 33149 8925 33183 8959
rect 33183 8925 33192 8959
rect 33140 8916 33192 8925
rect 33416 8959 33468 8968
rect 33416 8925 33425 8959
rect 33425 8925 33459 8959
rect 33459 8925 33468 8959
rect 33416 8916 33468 8925
rect 34704 8993 34713 9027
rect 34713 8993 34747 9027
rect 34747 8993 34756 9027
rect 34704 8984 34756 8993
rect 37924 8959 37976 8968
rect 37924 8925 37933 8959
rect 37933 8925 37967 8959
rect 37967 8925 37976 8959
rect 37924 8916 37976 8925
rect 58164 8959 58216 8968
rect 58164 8925 58173 8959
rect 58173 8925 58207 8959
rect 58207 8925 58216 8959
rect 58164 8916 58216 8925
rect 17316 8848 17368 8900
rect 19156 8848 19208 8900
rect 21180 8848 21232 8900
rect 28172 8848 28224 8900
rect 29736 8848 29788 8900
rect 29920 8891 29972 8900
rect 29920 8857 29929 8891
rect 29929 8857 29963 8891
rect 29963 8857 29972 8891
rect 29920 8848 29972 8857
rect 16672 8823 16724 8832
rect 16672 8789 16681 8823
rect 16681 8789 16715 8823
rect 16715 8789 16724 8823
rect 16672 8780 16724 8789
rect 17040 8780 17092 8832
rect 23388 8823 23440 8832
rect 23388 8789 23397 8823
rect 23397 8789 23431 8823
rect 23431 8789 23440 8823
rect 23388 8780 23440 8789
rect 28448 8780 28500 8832
rect 34980 8891 35032 8900
rect 34980 8857 35014 8891
rect 35014 8857 35032 8891
rect 30932 8780 30984 8832
rect 34980 8848 35032 8857
rect 36452 8848 36504 8900
rect 32496 8780 32548 8832
rect 36728 8780 36780 8832
rect 37556 8780 37608 8832
rect 38016 8848 38068 8900
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 7564 8576 7616 8628
rect 4620 8508 4672 8560
rect 9680 8551 9732 8560
rect 1676 8440 1728 8492
rect 5172 8440 5224 8492
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 1860 8372 1912 8424
rect 4988 8415 5040 8424
rect 4988 8381 4997 8415
rect 4997 8381 5031 8415
rect 5031 8381 5040 8415
rect 4988 8372 5040 8381
rect 2872 8236 2924 8288
rect 3976 8279 4028 8288
rect 3976 8245 3985 8279
rect 3985 8245 4019 8279
rect 4019 8245 4028 8279
rect 3976 8236 4028 8245
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 9680 8517 9714 8551
rect 9714 8517 9732 8551
rect 9680 8508 9732 8517
rect 11244 8576 11296 8628
rect 13728 8576 13780 8628
rect 16856 8576 16908 8628
rect 17316 8619 17368 8628
rect 17316 8585 17325 8619
rect 17325 8585 17359 8619
rect 17359 8585 17368 8619
rect 17316 8576 17368 8585
rect 11520 8551 11572 8560
rect 11520 8517 11529 8551
rect 11529 8517 11563 8551
rect 11563 8517 11572 8551
rect 11520 8508 11572 8517
rect 13820 8508 13872 8560
rect 16764 8551 16816 8560
rect 16764 8517 16773 8551
rect 16773 8517 16807 8551
rect 16807 8517 16816 8551
rect 16764 8508 16816 8517
rect 8852 8440 8904 8492
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 9496 8440 9548 8492
rect 13912 8440 13964 8492
rect 14740 8483 14792 8492
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 17500 8440 17552 8492
rect 17960 8483 18012 8492
rect 5540 8236 5592 8288
rect 7564 8236 7616 8288
rect 11704 8304 11756 8356
rect 13544 8347 13596 8356
rect 13544 8313 13553 8347
rect 13553 8313 13587 8347
rect 13587 8313 13596 8347
rect 13544 8304 13596 8313
rect 17960 8449 17969 8483
rect 17969 8449 18003 8483
rect 18003 8449 18012 8483
rect 17960 8440 18012 8449
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 19156 8576 19208 8628
rect 18328 8372 18380 8424
rect 18880 8372 18932 8424
rect 19156 8440 19208 8492
rect 20628 8508 20680 8560
rect 19432 8440 19484 8492
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 22836 8440 22888 8492
rect 23020 8440 23072 8492
rect 23388 8440 23440 8492
rect 24216 8508 24268 8560
rect 29736 8576 29788 8628
rect 32772 8576 32824 8628
rect 34980 8576 35032 8628
rect 38016 8619 38068 8628
rect 38016 8585 38025 8619
rect 38025 8585 38059 8619
rect 38059 8585 38068 8619
rect 38016 8576 38068 8585
rect 30564 8508 30616 8560
rect 30656 8551 30708 8560
rect 30656 8517 30674 8551
rect 30674 8517 30708 8551
rect 32588 8551 32640 8560
rect 30656 8508 30708 8517
rect 32588 8517 32597 8551
rect 32597 8517 32631 8551
rect 32631 8517 32640 8551
rect 32588 8508 32640 8517
rect 20076 8372 20128 8424
rect 21088 8372 21140 8424
rect 9588 8236 9640 8288
rect 9772 8236 9824 8288
rect 15016 8304 15068 8356
rect 18972 8304 19024 8356
rect 23388 8304 23440 8356
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 24584 8440 24636 8492
rect 26332 8440 26384 8492
rect 27436 8483 27488 8492
rect 27436 8449 27445 8483
rect 27445 8449 27479 8483
rect 27479 8449 27488 8483
rect 27436 8440 27488 8449
rect 28448 8483 28500 8492
rect 28172 8415 28224 8424
rect 28172 8381 28181 8415
rect 28181 8381 28215 8415
rect 28215 8381 28224 8415
rect 28172 8372 28224 8381
rect 28448 8449 28457 8483
rect 28457 8449 28491 8483
rect 28491 8449 28500 8483
rect 28448 8440 28500 8449
rect 28540 8372 28592 8424
rect 26792 8304 26844 8356
rect 30932 8415 30984 8424
rect 30932 8381 30941 8415
rect 30941 8381 30975 8415
rect 30975 8381 30984 8415
rect 30932 8372 30984 8381
rect 32404 8440 32456 8492
rect 32496 8483 32548 8492
rect 32496 8449 32505 8483
rect 32505 8449 32539 8483
rect 32539 8449 32548 8483
rect 32496 8440 32548 8449
rect 32680 8483 32732 8492
rect 32680 8449 32689 8483
rect 32689 8449 32723 8483
rect 32723 8449 32732 8483
rect 35808 8508 35860 8560
rect 32680 8440 32732 8449
rect 35348 8483 35400 8492
rect 35348 8449 35357 8483
rect 35357 8449 35391 8483
rect 35391 8449 35400 8483
rect 35348 8440 35400 8449
rect 35532 8483 35584 8492
rect 35532 8449 35541 8483
rect 35541 8449 35575 8483
rect 35575 8449 35584 8483
rect 35532 8440 35584 8449
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 38384 8508 38436 8560
rect 37740 8483 37792 8492
rect 37740 8449 37749 8483
rect 37749 8449 37783 8483
rect 37783 8449 37792 8483
rect 37740 8440 37792 8449
rect 35624 8372 35676 8424
rect 14188 8279 14240 8288
rect 14188 8245 14197 8279
rect 14197 8245 14231 8279
rect 14231 8245 14240 8279
rect 14188 8236 14240 8245
rect 14924 8279 14976 8288
rect 14924 8245 14933 8279
rect 14933 8245 14967 8279
rect 14967 8245 14976 8279
rect 14924 8236 14976 8245
rect 18236 8236 18288 8288
rect 18604 8236 18656 8288
rect 19156 8236 19208 8288
rect 23572 8236 23624 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 2320 8032 2372 8084
rect 5356 8075 5408 8084
rect 5356 8041 5365 8075
rect 5365 8041 5399 8075
rect 5399 8041 5408 8075
rect 5356 8032 5408 8041
rect 7288 8032 7340 8084
rect 7932 8032 7984 8084
rect 8300 8032 8352 8084
rect 9496 8032 9548 8084
rect 16580 8032 16632 8084
rect 18328 8075 18380 8084
rect 18328 8041 18337 8075
rect 18337 8041 18371 8075
rect 18371 8041 18380 8075
rect 18328 8032 18380 8041
rect 23940 8032 23992 8084
rect 26240 8032 26292 8084
rect 27436 8032 27488 8084
rect 29000 8075 29052 8084
rect 29000 8041 29009 8075
rect 29009 8041 29043 8075
rect 29043 8041 29052 8075
rect 29000 8032 29052 8041
rect 32312 8032 32364 8084
rect 2872 7939 2924 7948
rect 2872 7905 2881 7939
rect 2881 7905 2915 7939
rect 2915 7905 2924 7939
rect 2872 7896 2924 7905
rect 9404 7964 9456 8016
rect 12072 7964 12124 8016
rect 2964 7828 3016 7880
rect 5540 7896 5592 7948
rect 18052 7896 18104 7948
rect 5632 7828 5684 7880
rect 6276 7871 6328 7880
rect 6276 7837 6285 7871
rect 6285 7837 6319 7871
rect 6319 7837 6328 7871
rect 6276 7828 6328 7837
rect 6552 7871 6604 7880
rect 6552 7837 6586 7871
rect 6586 7837 6604 7871
rect 6552 7828 6604 7837
rect 7104 7828 7156 7880
rect 4620 7760 4672 7812
rect 4988 7760 5040 7812
rect 1768 7692 1820 7744
rect 3976 7692 4028 7744
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 9496 7692 9548 7744
rect 15108 7828 15160 7880
rect 19064 7828 19116 7880
rect 23572 7871 23624 7880
rect 23572 7837 23590 7871
rect 23590 7837 23624 7871
rect 23572 7828 23624 7837
rect 25136 7828 25188 7880
rect 25872 7828 25924 7880
rect 28724 7896 28776 7948
rect 29644 7964 29696 8016
rect 37740 8032 37792 8084
rect 28448 7871 28500 7880
rect 28448 7837 28457 7871
rect 28457 7837 28491 7871
rect 28491 7837 28500 7871
rect 28448 7828 28500 7837
rect 31392 7871 31444 7880
rect 10876 7692 10928 7744
rect 12716 7692 12768 7744
rect 13728 7692 13780 7744
rect 14740 7692 14792 7744
rect 15660 7803 15712 7812
rect 15660 7769 15694 7803
rect 15694 7769 15712 7803
rect 15660 7760 15712 7769
rect 17960 7760 18012 7812
rect 18604 7760 18656 7812
rect 16764 7735 16816 7744
rect 16764 7701 16773 7735
rect 16773 7701 16807 7735
rect 16807 7701 16816 7735
rect 16764 7692 16816 7701
rect 20536 7760 20588 7812
rect 19432 7692 19484 7744
rect 20352 7735 20404 7744
rect 20352 7701 20361 7735
rect 20361 7701 20395 7735
rect 20395 7701 20404 7735
rect 20352 7692 20404 7701
rect 21640 7735 21692 7744
rect 21640 7701 21649 7735
rect 21649 7701 21683 7735
rect 21683 7701 21692 7735
rect 21640 7692 21692 7701
rect 22744 7692 22796 7744
rect 24676 7760 24728 7812
rect 25596 7803 25648 7812
rect 25596 7769 25630 7803
rect 25630 7769 25648 7803
rect 25596 7760 25648 7769
rect 28172 7760 28224 7812
rect 31392 7837 31401 7871
rect 31401 7837 31435 7871
rect 31435 7837 31444 7871
rect 31392 7828 31444 7837
rect 34796 7828 34848 7880
rect 35256 7871 35308 7880
rect 35256 7837 35265 7871
rect 35265 7837 35299 7871
rect 35299 7837 35308 7871
rect 35256 7828 35308 7837
rect 36268 7828 36320 7880
rect 58164 7871 58216 7880
rect 58164 7837 58173 7871
rect 58173 7837 58207 7871
rect 58207 7837 58216 7871
rect 58164 7828 58216 7837
rect 30288 7692 30340 7744
rect 35440 7803 35492 7812
rect 35440 7769 35449 7803
rect 35449 7769 35483 7803
rect 35483 7769 35492 7803
rect 35440 7760 35492 7769
rect 37096 7692 37148 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 6184 7488 6236 7540
rect 6552 7488 6604 7540
rect 3424 7420 3476 7472
rect 3700 7395 3752 7404
rect 3700 7361 3709 7395
rect 3709 7361 3743 7395
rect 3743 7361 3752 7395
rect 3700 7352 3752 7361
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 6368 7352 6420 7404
rect 7380 7420 7432 7472
rect 7564 7463 7616 7472
rect 7564 7429 7573 7463
rect 7573 7429 7607 7463
rect 7607 7429 7616 7463
rect 7564 7420 7616 7429
rect 12532 7488 12584 7540
rect 6920 7395 6972 7404
rect 6920 7361 6929 7395
rect 6929 7361 6963 7395
rect 6963 7361 6972 7395
rect 6920 7352 6972 7361
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 7932 7395 7984 7404
rect 7932 7361 7941 7395
rect 7941 7361 7975 7395
rect 7975 7361 7984 7395
rect 7932 7352 7984 7361
rect 11888 7420 11940 7472
rect 12072 7395 12124 7404
rect 12072 7361 12081 7395
rect 12081 7361 12115 7395
rect 12115 7361 12124 7395
rect 12072 7352 12124 7361
rect 5356 7284 5408 7336
rect 5908 7284 5960 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 2596 7148 2648 7200
rect 4896 7216 4948 7268
rect 5264 7216 5316 7268
rect 6644 7216 6696 7268
rect 10048 7216 10100 7268
rect 14188 7395 14240 7404
rect 14188 7361 14197 7395
rect 14197 7361 14231 7395
rect 14231 7361 14240 7395
rect 14924 7395 14976 7404
rect 14188 7352 14240 7361
rect 14924 7361 14933 7395
rect 14933 7361 14967 7395
rect 14967 7361 14976 7395
rect 14924 7352 14976 7361
rect 15660 7488 15712 7540
rect 17592 7488 17644 7540
rect 18144 7488 18196 7540
rect 18512 7488 18564 7540
rect 16764 7420 16816 7472
rect 17040 7395 17092 7404
rect 14556 7284 14608 7336
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 3148 7148 3200 7200
rect 3516 7191 3568 7200
rect 3516 7157 3525 7191
rect 3525 7157 3559 7191
rect 3559 7157 3568 7191
rect 3516 7148 3568 7157
rect 3976 7148 4028 7200
rect 4252 7148 4304 7200
rect 7748 7148 7800 7200
rect 8576 7148 8628 7200
rect 10324 7148 10376 7200
rect 10876 7148 10928 7200
rect 15936 7216 15988 7268
rect 13176 7148 13228 7200
rect 13452 7191 13504 7200
rect 13452 7157 13461 7191
rect 13461 7157 13495 7191
rect 13495 7157 13504 7191
rect 13452 7148 13504 7157
rect 14096 7191 14148 7200
rect 14096 7157 14105 7191
rect 14105 7157 14139 7191
rect 14139 7157 14148 7191
rect 14096 7148 14148 7157
rect 18144 7327 18196 7336
rect 18144 7293 18153 7327
rect 18153 7293 18187 7327
rect 18187 7293 18196 7327
rect 18144 7284 18196 7293
rect 19432 7352 19484 7404
rect 20168 7352 20220 7404
rect 20444 7352 20496 7404
rect 18880 7284 18932 7336
rect 21180 7352 21232 7404
rect 21640 7352 21692 7404
rect 22192 7420 22244 7472
rect 22744 7463 22796 7472
rect 22744 7429 22753 7463
rect 22753 7429 22787 7463
rect 22787 7429 22796 7463
rect 22744 7420 22796 7429
rect 24124 7488 24176 7540
rect 24676 7488 24728 7540
rect 25596 7531 25648 7540
rect 22836 7395 22888 7404
rect 22836 7361 22845 7395
rect 22845 7361 22879 7395
rect 22879 7361 22888 7395
rect 22836 7352 22888 7361
rect 22928 7352 22980 7404
rect 24216 7420 24268 7472
rect 25596 7497 25605 7531
rect 25605 7497 25639 7531
rect 25639 7497 25648 7531
rect 25596 7488 25648 7497
rect 28356 7488 28408 7540
rect 31392 7488 31444 7540
rect 34520 7488 34572 7540
rect 38108 7531 38160 7540
rect 38108 7497 38117 7531
rect 38117 7497 38151 7531
rect 38151 7497 38160 7531
rect 38108 7488 38160 7497
rect 24400 7352 24452 7404
rect 24584 7352 24636 7404
rect 26240 7463 26292 7472
rect 26240 7429 26249 7463
rect 26249 7429 26283 7463
rect 26283 7429 26292 7463
rect 26240 7420 26292 7429
rect 20444 7216 20496 7268
rect 24676 7284 24728 7336
rect 25320 7395 25372 7404
rect 25320 7361 25329 7395
rect 25329 7361 25363 7395
rect 25363 7361 25372 7395
rect 29644 7420 29696 7472
rect 31300 7420 31352 7472
rect 33600 7463 33652 7472
rect 33600 7429 33618 7463
rect 33618 7429 33652 7463
rect 35440 7463 35492 7472
rect 33600 7420 33652 7429
rect 35440 7429 35449 7463
rect 35449 7429 35483 7463
rect 35483 7429 35492 7463
rect 35440 7420 35492 7429
rect 37648 7420 37700 7472
rect 25320 7352 25372 7361
rect 27344 7352 27396 7404
rect 31116 7352 31168 7404
rect 35256 7395 35308 7404
rect 35256 7361 35265 7395
rect 35265 7361 35299 7395
rect 35299 7361 35308 7395
rect 35256 7352 35308 7361
rect 35624 7395 35676 7404
rect 27252 7327 27304 7336
rect 27252 7293 27261 7327
rect 27261 7293 27295 7327
rect 27295 7293 27304 7327
rect 27252 7284 27304 7293
rect 34796 7284 34848 7336
rect 35624 7361 35633 7395
rect 35633 7361 35667 7395
rect 35667 7361 35676 7395
rect 35624 7352 35676 7361
rect 39672 7284 39724 7336
rect 25320 7216 25372 7268
rect 19248 7148 19300 7200
rect 20168 7148 20220 7200
rect 21272 7191 21324 7200
rect 21272 7157 21281 7191
rect 21281 7157 21315 7191
rect 21315 7157 21324 7191
rect 21272 7148 21324 7157
rect 21916 7191 21968 7200
rect 21916 7157 21925 7191
rect 21925 7157 21959 7191
rect 21959 7157 21968 7191
rect 21916 7148 21968 7157
rect 23664 7148 23716 7200
rect 29644 7148 29696 7200
rect 38844 7148 38896 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 4068 6944 4120 6996
rect 14096 6944 14148 6996
rect 21180 6944 21232 6996
rect 21272 6944 21324 6996
rect 26976 6944 27028 6996
rect 3332 6740 3384 6792
rect 3976 6808 4028 6860
rect 4528 6740 4580 6792
rect 4620 6740 4672 6792
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 8668 6808 8720 6860
rect 9864 6876 9916 6928
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 8576 6740 8628 6792
rect 9956 6783 10008 6792
rect 3056 6672 3108 6724
rect 9496 6672 9548 6724
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 13360 6808 13412 6860
rect 15476 6851 15528 6860
rect 15476 6817 15485 6851
rect 15485 6817 15519 6851
rect 15519 6817 15528 6851
rect 19432 6876 19484 6928
rect 23940 6876 23992 6928
rect 24584 6876 24636 6928
rect 15476 6808 15528 6817
rect 20168 6808 20220 6860
rect 22652 6808 22704 6860
rect 10140 6740 10192 6749
rect 10508 6740 10560 6792
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 12348 6740 12400 6792
rect 12440 6740 12492 6792
rect 13544 6740 13596 6792
rect 14556 6783 14608 6792
rect 14556 6749 14565 6783
rect 14565 6749 14599 6783
rect 14599 6749 14608 6783
rect 14556 6740 14608 6749
rect 14648 6783 14700 6792
rect 14648 6749 14662 6783
rect 14662 6749 14696 6783
rect 14696 6749 14700 6783
rect 14648 6740 14700 6749
rect 14924 6740 14976 6792
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 11060 6672 11112 6724
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 4528 6604 4580 6656
rect 5172 6604 5224 6656
rect 7012 6604 7064 6656
rect 8208 6604 8260 6656
rect 8484 6604 8536 6656
rect 9128 6647 9180 6656
rect 9128 6613 9137 6647
rect 9137 6613 9171 6647
rect 9171 6613 9180 6647
rect 9128 6604 9180 6613
rect 9864 6604 9916 6656
rect 12900 6672 12952 6724
rect 14096 6672 14148 6724
rect 13912 6604 13964 6656
rect 14004 6604 14056 6656
rect 14924 6604 14976 6656
rect 17776 6740 17828 6792
rect 18236 6740 18288 6792
rect 21640 6783 21692 6792
rect 20168 6672 20220 6724
rect 21640 6749 21649 6783
rect 21649 6749 21683 6783
rect 21683 6749 21692 6783
rect 21640 6740 21692 6749
rect 23388 6740 23440 6792
rect 23664 6783 23716 6792
rect 23664 6749 23673 6783
rect 23673 6749 23707 6783
rect 23707 6749 23716 6783
rect 23664 6740 23716 6749
rect 23940 6740 23992 6792
rect 24952 6808 25004 6860
rect 24584 6740 24636 6792
rect 27252 6876 27304 6928
rect 30932 6944 30984 6996
rect 31300 6987 31352 6996
rect 31300 6953 31309 6987
rect 31309 6953 31343 6987
rect 31343 6953 31352 6987
rect 31300 6944 31352 6953
rect 25964 6851 26016 6860
rect 25964 6817 25973 6851
rect 25973 6817 26007 6851
rect 26007 6817 26016 6851
rect 25964 6808 26016 6817
rect 27068 6808 27120 6860
rect 27528 6783 27580 6792
rect 24216 6672 24268 6724
rect 17592 6647 17644 6656
rect 17592 6613 17601 6647
rect 17601 6613 17635 6647
rect 17635 6613 17644 6647
rect 17592 6604 17644 6613
rect 18328 6647 18380 6656
rect 18328 6613 18337 6647
rect 18337 6613 18371 6647
rect 18371 6613 18380 6647
rect 18328 6604 18380 6613
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 20720 6647 20772 6656
rect 20720 6613 20729 6647
rect 20729 6613 20763 6647
rect 20763 6613 20772 6647
rect 20720 6604 20772 6613
rect 23572 6604 23624 6656
rect 24768 6604 24820 6656
rect 27528 6749 27537 6783
rect 27537 6749 27571 6783
rect 27571 6749 27580 6783
rect 27528 6740 27580 6749
rect 38568 6944 38620 6996
rect 38752 6944 38804 6996
rect 27344 6672 27396 6724
rect 28172 6740 28224 6792
rect 31116 6740 31168 6792
rect 28356 6672 28408 6724
rect 30196 6715 30248 6724
rect 30196 6681 30230 6715
rect 30230 6681 30248 6715
rect 30196 6672 30248 6681
rect 27528 6604 27580 6656
rect 28724 6604 28776 6656
rect 35808 6876 35860 6928
rect 34152 6715 34204 6724
rect 34152 6681 34161 6715
rect 34161 6681 34195 6715
rect 34195 6681 34204 6715
rect 34152 6672 34204 6681
rect 35532 6783 35584 6792
rect 35532 6749 35541 6783
rect 35541 6749 35575 6783
rect 35575 6749 35584 6783
rect 35532 6740 35584 6749
rect 36820 6783 36872 6792
rect 36820 6749 36829 6783
rect 36829 6749 36863 6783
rect 36863 6749 36872 6783
rect 36820 6740 36872 6749
rect 39028 6876 39080 6928
rect 37004 6783 37056 6792
rect 37004 6749 37013 6783
rect 37013 6749 37047 6783
rect 37047 6749 37056 6783
rect 37004 6740 37056 6749
rect 38568 6740 38620 6792
rect 38108 6672 38160 6724
rect 38844 6783 38896 6792
rect 38844 6749 38858 6783
rect 38858 6749 38892 6783
rect 38892 6749 38896 6783
rect 38844 6740 38896 6749
rect 34520 6604 34572 6656
rect 35440 6604 35492 6656
rect 37556 6604 37608 6656
rect 38384 6647 38436 6656
rect 38384 6613 38393 6647
rect 38393 6613 38427 6647
rect 38427 6613 38436 6647
rect 38384 6604 38436 6613
rect 38936 6672 38988 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 6460 6400 6512 6452
rect 11520 6400 11572 6452
rect 11980 6400 12032 6452
rect 14648 6400 14700 6452
rect 16028 6400 16080 6452
rect 22008 6400 22060 6452
rect 23480 6400 23532 6452
rect 27436 6400 27488 6452
rect 29092 6400 29144 6452
rect 30012 6400 30064 6452
rect 30196 6443 30248 6452
rect 30196 6409 30205 6443
rect 30205 6409 30239 6443
rect 30239 6409 30248 6443
rect 30196 6400 30248 6409
rect 34152 6400 34204 6452
rect 36820 6400 36872 6452
rect 39672 6443 39724 6452
rect 39672 6409 39681 6443
rect 39681 6409 39715 6443
rect 39715 6409 39724 6443
rect 39672 6400 39724 6409
rect 3792 6332 3844 6384
rect 5540 6332 5592 6384
rect 6276 6332 6328 6384
rect 9864 6375 9916 6384
rect 9864 6341 9898 6375
rect 9898 6341 9916 6375
rect 9864 6332 9916 6341
rect 19064 6375 19116 6384
rect 2504 6307 2556 6316
rect 2504 6273 2513 6307
rect 2513 6273 2547 6307
rect 2547 6273 2556 6307
rect 2504 6264 2556 6273
rect 5356 6264 5408 6316
rect 7380 6264 7432 6316
rect 7656 6264 7708 6316
rect 8484 6264 8536 6316
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 9404 6264 9456 6316
rect 19064 6341 19073 6375
rect 19073 6341 19107 6375
rect 19107 6341 19116 6375
rect 19064 6332 19116 6341
rect 19340 6332 19392 6384
rect 19524 6375 19576 6384
rect 19524 6341 19533 6375
rect 19533 6341 19567 6375
rect 19567 6341 19576 6375
rect 19524 6332 19576 6341
rect 22192 6332 22244 6384
rect 23756 6332 23808 6384
rect 33140 6332 33192 6384
rect 34428 6375 34480 6384
rect 34428 6341 34437 6375
rect 34437 6341 34471 6375
rect 34471 6341 34480 6375
rect 34428 6332 34480 6341
rect 6828 6196 6880 6248
rect 6000 6128 6052 6180
rect 8024 6196 8076 6248
rect 8668 6128 8720 6180
rect 11060 6128 11112 6180
rect 11980 6128 12032 6180
rect 14004 6307 14056 6316
rect 14004 6273 14038 6307
rect 14038 6273 14056 6307
rect 14004 6264 14056 6273
rect 2044 6060 2096 6112
rect 2136 6060 2188 6112
rect 5632 6103 5684 6112
rect 5632 6069 5641 6103
rect 5641 6069 5675 6103
rect 5675 6069 5684 6103
rect 5632 6060 5684 6069
rect 7564 6060 7616 6112
rect 7840 6060 7892 6112
rect 8852 6103 8904 6112
rect 8852 6069 8861 6103
rect 8861 6069 8895 6103
rect 8895 6069 8904 6103
rect 8852 6060 8904 6069
rect 11612 6103 11664 6112
rect 11612 6069 11621 6103
rect 11621 6069 11655 6103
rect 11655 6069 11664 6103
rect 11612 6060 11664 6069
rect 12164 6060 12216 6112
rect 12992 6060 13044 6112
rect 15752 6128 15804 6180
rect 16580 6264 16632 6316
rect 20628 6264 20680 6316
rect 23112 6307 23164 6316
rect 23112 6273 23121 6307
rect 23121 6273 23155 6307
rect 23155 6273 23164 6307
rect 23112 6264 23164 6273
rect 17040 6196 17092 6248
rect 18604 6196 18656 6248
rect 21640 6196 21692 6248
rect 22192 6196 22244 6248
rect 22836 6196 22888 6248
rect 24860 6264 24912 6316
rect 26976 6307 27028 6316
rect 26976 6273 26985 6307
rect 26985 6273 27019 6307
rect 27019 6273 27028 6307
rect 26976 6264 27028 6273
rect 27528 6264 27580 6316
rect 29552 6307 29604 6316
rect 29552 6273 29561 6307
rect 29561 6273 29595 6307
rect 29595 6273 29604 6307
rect 29552 6264 29604 6273
rect 29644 6264 29696 6316
rect 24584 6196 24636 6248
rect 28724 6196 28776 6248
rect 28816 6196 28868 6248
rect 29092 6196 29144 6248
rect 30012 6264 30064 6316
rect 31116 6264 31168 6316
rect 35808 6332 35860 6384
rect 36268 6375 36320 6384
rect 36268 6341 36277 6375
rect 36277 6341 36311 6375
rect 36311 6341 36320 6375
rect 36268 6332 36320 6341
rect 36452 6375 36504 6384
rect 36452 6341 36461 6375
rect 36461 6341 36495 6375
rect 36495 6341 36504 6375
rect 36452 6332 36504 6341
rect 37648 6375 37700 6384
rect 37648 6341 37657 6375
rect 37657 6341 37691 6375
rect 37691 6341 37700 6375
rect 37648 6332 37700 6341
rect 38384 6332 38436 6384
rect 18512 6128 18564 6180
rect 18696 6060 18748 6112
rect 20076 6060 20128 6112
rect 20812 6060 20864 6112
rect 21180 6103 21232 6112
rect 21180 6069 21189 6103
rect 21189 6069 21223 6103
rect 21223 6069 21232 6103
rect 21180 6060 21232 6069
rect 22008 6128 22060 6180
rect 25596 6128 25648 6180
rect 23112 6060 23164 6112
rect 23388 6060 23440 6112
rect 26148 6103 26200 6112
rect 26148 6069 26157 6103
rect 26157 6069 26191 6103
rect 26191 6069 26200 6103
rect 26148 6060 26200 6069
rect 28172 6128 28224 6180
rect 29828 6128 29880 6180
rect 35532 6264 35584 6316
rect 37188 6264 37240 6316
rect 37924 6264 37976 6316
rect 37004 6128 37056 6180
rect 58164 6171 58216 6180
rect 58164 6137 58173 6171
rect 58173 6137 58207 6171
rect 58207 6137 58216 6171
rect 58164 6128 58216 6137
rect 29368 6060 29420 6112
rect 30196 6060 30248 6112
rect 34704 6060 34756 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 6920 5856 6972 5908
rect 4804 5788 4856 5840
rect 12440 5856 12492 5908
rect 18604 5856 18656 5908
rect 19432 5856 19484 5908
rect 20628 5899 20680 5908
rect 20628 5865 20637 5899
rect 20637 5865 20671 5899
rect 20671 5865 20680 5899
rect 20628 5856 20680 5865
rect 10784 5788 10836 5840
rect 11336 5831 11388 5840
rect 11336 5797 11345 5831
rect 11345 5797 11379 5831
rect 11379 5797 11388 5831
rect 11336 5788 11388 5797
rect 1860 5695 1912 5704
rect 1860 5661 1869 5695
rect 1869 5661 1903 5695
rect 1903 5661 1912 5695
rect 1860 5652 1912 5661
rect 2136 5695 2188 5704
rect 2136 5661 2170 5695
rect 2170 5661 2188 5695
rect 2136 5652 2188 5661
rect 3240 5652 3292 5704
rect 4712 5720 4764 5772
rect 6552 5720 6604 5772
rect 10232 5720 10284 5772
rect 2688 5584 2740 5636
rect 6368 5695 6420 5704
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 9956 5652 10008 5704
rect 11336 5652 11388 5704
rect 11520 5695 11572 5704
rect 11520 5661 11529 5695
rect 11529 5661 11563 5695
rect 11563 5661 11572 5695
rect 11520 5652 11572 5661
rect 6644 5584 6696 5636
rect 7012 5584 7064 5636
rect 8300 5584 8352 5636
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 13268 5652 13320 5704
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 14924 5652 14976 5704
rect 23296 5856 23348 5908
rect 24768 5899 24820 5908
rect 24768 5865 24777 5899
rect 24777 5865 24811 5899
rect 24811 5865 24820 5899
rect 24768 5856 24820 5865
rect 29184 5856 29236 5908
rect 30564 5856 30616 5908
rect 33140 5856 33192 5908
rect 34520 5856 34572 5908
rect 35532 5856 35584 5908
rect 36268 5856 36320 5908
rect 37188 5856 37240 5908
rect 27712 5788 27764 5840
rect 15752 5720 15804 5772
rect 17868 5720 17920 5772
rect 14556 5584 14608 5636
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 17776 5652 17828 5704
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 19064 5720 19116 5772
rect 23388 5720 23440 5772
rect 25596 5763 25648 5772
rect 25596 5729 25605 5763
rect 25605 5729 25639 5763
rect 25639 5729 25648 5763
rect 25596 5720 25648 5729
rect 30196 5720 30248 5772
rect 4988 5516 5040 5568
rect 5448 5516 5500 5568
rect 14832 5516 14884 5568
rect 16120 5516 16172 5568
rect 17040 5584 17092 5636
rect 17684 5584 17736 5636
rect 18144 5584 18196 5636
rect 18696 5652 18748 5704
rect 22192 5652 22244 5704
rect 22836 5652 22888 5704
rect 23756 5652 23808 5704
rect 27528 5652 27580 5704
rect 29552 5652 29604 5704
rect 19340 5584 19392 5636
rect 22928 5584 22980 5636
rect 24400 5627 24452 5636
rect 24400 5593 24409 5627
rect 24409 5593 24443 5627
rect 24443 5593 24452 5627
rect 24400 5584 24452 5593
rect 27068 5584 27120 5636
rect 29828 5584 29880 5636
rect 30564 5652 30616 5704
rect 31024 5652 31076 5704
rect 34796 5695 34848 5704
rect 34796 5661 34805 5695
rect 34805 5661 34839 5695
rect 34839 5661 34848 5695
rect 34796 5652 34848 5661
rect 37556 5652 37608 5704
rect 34704 5584 34756 5636
rect 18512 5516 18564 5568
rect 21640 5559 21692 5568
rect 21640 5525 21649 5559
rect 21649 5525 21683 5559
rect 21683 5525 21692 5559
rect 21640 5516 21692 5525
rect 23480 5516 23532 5568
rect 24860 5516 24912 5568
rect 29000 5516 29052 5568
rect 30288 5516 30340 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 2504 5355 2556 5364
rect 2504 5321 2513 5355
rect 2513 5321 2547 5355
rect 2547 5321 2556 5355
rect 2504 5312 2556 5321
rect 4988 5355 5040 5364
rect 4988 5321 4997 5355
rect 4997 5321 5031 5355
rect 5031 5321 5040 5355
rect 4988 5312 5040 5321
rect 5632 5312 5684 5364
rect 6368 5312 6420 5364
rect 6552 5355 6604 5364
rect 6552 5321 6561 5355
rect 6561 5321 6595 5355
rect 6595 5321 6604 5355
rect 6552 5312 6604 5321
rect 14280 5312 14332 5364
rect 17592 5312 17644 5364
rect 2688 5219 2740 5228
rect 2688 5185 2697 5219
rect 2697 5185 2731 5219
rect 2731 5185 2740 5219
rect 2688 5176 2740 5185
rect 3976 5176 4028 5228
rect 4804 5176 4856 5228
rect 4988 5176 5040 5228
rect 5356 5176 5408 5228
rect 6368 5219 6420 5228
rect 4528 5108 4580 5160
rect 4712 5108 4764 5160
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 6460 5176 6512 5228
rect 7840 5244 7892 5296
rect 18236 5312 18288 5364
rect 6920 5219 6972 5228
rect 6920 5185 6929 5219
rect 6929 5185 6963 5219
rect 6963 5185 6972 5219
rect 6920 5176 6972 5185
rect 7472 5176 7524 5228
rect 5356 4972 5408 5024
rect 6276 5040 6328 5092
rect 6460 4972 6512 5024
rect 8024 5176 8076 5228
rect 10968 5176 11020 5228
rect 11520 5176 11572 5228
rect 12072 5176 12124 5228
rect 14740 5176 14792 5228
rect 15016 5219 15068 5228
rect 15016 5185 15025 5219
rect 15025 5185 15059 5219
rect 15059 5185 15068 5219
rect 15016 5176 15068 5185
rect 17776 5219 17828 5228
rect 17776 5185 17785 5219
rect 17785 5185 17819 5219
rect 17819 5185 17828 5219
rect 17776 5176 17828 5185
rect 17868 5176 17920 5228
rect 20996 5312 21048 5364
rect 23756 5355 23808 5364
rect 23756 5321 23765 5355
rect 23765 5321 23799 5355
rect 23799 5321 23808 5355
rect 23756 5312 23808 5321
rect 25596 5355 25648 5364
rect 25596 5321 25605 5355
rect 25605 5321 25639 5355
rect 25639 5321 25648 5355
rect 25596 5312 25648 5321
rect 34796 5312 34848 5364
rect 19524 5244 19576 5296
rect 24952 5244 25004 5296
rect 27988 5287 28040 5296
rect 27988 5253 27997 5287
rect 27997 5253 28031 5287
rect 28031 5253 28040 5287
rect 27988 5244 28040 5253
rect 28448 5244 28500 5296
rect 29000 5244 29052 5296
rect 29920 5244 29972 5296
rect 25136 5219 25188 5228
rect 7104 5040 7156 5092
rect 8760 5108 8812 5160
rect 11244 5108 11296 5160
rect 12440 5108 12492 5160
rect 17684 5108 17736 5160
rect 25136 5185 25145 5219
rect 25145 5185 25179 5219
rect 25179 5185 25188 5219
rect 25136 5176 25188 5185
rect 26148 5176 26200 5228
rect 28172 5219 28224 5228
rect 28172 5185 28181 5219
rect 28181 5185 28215 5219
rect 28215 5185 28224 5219
rect 28172 5176 28224 5185
rect 8484 5083 8536 5092
rect 8484 5049 8493 5083
rect 8493 5049 8527 5083
rect 8527 5049 8536 5083
rect 8484 5040 8536 5049
rect 15844 5040 15896 5092
rect 7932 4972 7984 5024
rect 8852 4972 8904 5024
rect 11888 4972 11940 5024
rect 12256 5015 12308 5024
rect 12256 4981 12265 5015
rect 12265 4981 12299 5015
rect 12299 4981 12308 5015
rect 12256 4972 12308 4981
rect 13820 4972 13872 5024
rect 14188 5015 14240 5024
rect 14188 4981 14197 5015
rect 14197 4981 14231 5015
rect 14231 4981 14240 5015
rect 14188 4972 14240 4981
rect 14832 5015 14884 5024
rect 14832 4981 14841 5015
rect 14841 4981 14875 5015
rect 14875 4981 14884 5015
rect 14832 4972 14884 4981
rect 15660 4972 15712 5024
rect 17592 4972 17644 5024
rect 17868 4972 17920 5024
rect 20076 5108 20128 5160
rect 53748 5108 53800 5160
rect 19340 5040 19392 5092
rect 20076 4972 20128 5024
rect 20904 4972 20956 5024
rect 21732 4972 21784 5024
rect 22560 4972 22612 5024
rect 23020 4972 23072 5024
rect 31576 5040 31628 5092
rect 54116 5040 54168 5092
rect 27344 4972 27396 5024
rect 53656 4972 53708 5024
rect 58164 5015 58216 5024
rect 58164 4981 58173 5015
rect 58173 4981 58207 5015
rect 58207 4981 58216 5015
rect 58164 4972 58216 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4620 4768 4672 4820
rect 5356 4768 5408 4820
rect 5632 4768 5684 4820
rect 6920 4811 6972 4820
rect 6920 4777 6929 4811
rect 6929 4777 6963 4811
rect 6963 4777 6972 4811
rect 6920 4768 6972 4777
rect 7104 4768 7156 4820
rect 6276 4700 6328 4752
rect 5816 4632 5868 4684
rect 7104 4632 7156 4684
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 3332 4564 3384 4616
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 5172 4564 5224 4616
rect 6736 4564 6788 4616
rect 7472 4768 7524 4820
rect 7932 4811 7984 4820
rect 7932 4777 7941 4811
rect 7941 4777 7975 4811
rect 7975 4777 7984 4811
rect 7932 4768 7984 4777
rect 8392 4768 8444 4820
rect 8944 4811 8996 4820
rect 8944 4777 8953 4811
rect 8953 4777 8987 4811
rect 8987 4777 8996 4811
rect 8944 4768 8996 4777
rect 9312 4768 9364 4820
rect 10876 4768 10928 4820
rect 7288 4700 7340 4752
rect 11428 4768 11480 4820
rect 11520 4700 11572 4752
rect 11796 4768 11848 4820
rect 21088 4768 21140 4820
rect 22928 4768 22980 4820
rect 23204 4768 23256 4820
rect 42064 4768 42116 4820
rect 12256 4700 12308 4752
rect 18696 4700 18748 4752
rect 26424 4743 26476 4752
rect 26424 4709 26433 4743
rect 26433 4709 26467 4743
rect 26467 4709 26476 4743
rect 26424 4700 26476 4709
rect 52184 4700 52236 4752
rect 53932 4700 53984 4752
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 7840 4564 7892 4616
rect 8852 4564 8904 4616
rect 3976 4496 4028 4548
rect 7104 4496 7156 4548
rect 3240 4428 3292 4480
rect 4344 4428 4396 4480
rect 4528 4471 4580 4480
rect 4528 4437 4537 4471
rect 4537 4437 4571 4471
rect 4571 4437 4580 4471
rect 4528 4428 4580 4437
rect 5908 4428 5960 4480
rect 6552 4428 6604 4480
rect 8208 4428 8260 4480
rect 9404 4632 9456 4684
rect 12072 4632 12124 4684
rect 13544 4632 13596 4684
rect 17040 4632 17092 4684
rect 18972 4632 19024 4684
rect 25136 4632 25188 4684
rect 11244 4607 11296 4616
rect 11244 4573 11253 4607
rect 11253 4573 11287 4607
rect 11287 4573 11296 4607
rect 11244 4564 11296 4573
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 14280 4564 14332 4616
rect 15384 4564 15436 4616
rect 15936 4564 15988 4616
rect 11520 4496 11572 4548
rect 19248 4564 19300 4616
rect 19340 4564 19392 4616
rect 20628 4564 20680 4616
rect 21088 4564 21140 4616
rect 21916 4564 21968 4616
rect 22192 4564 22244 4616
rect 23572 4607 23624 4616
rect 23572 4573 23590 4607
rect 23590 4573 23624 4607
rect 23572 4564 23624 4573
rect 18052 4496 18104 4548
rect 23296 4496 23348 4548
rect 23756 4496 23808 4548
rect 13912 4428 13964 4480
rect 17868 4428 17920 4480
rect 22376 4428 22428 4480
rect 27068 4632 27120 4684
rect 27344 4607 27396 4616
rect 27344 4573 27353 4607
rect 27353 4573 27387 4607
rect 27387 4573 27396 4607
rect 27344 4564 27396 4573
rect 27528 4607 27580 4616
rect 27528 4573 27537 4607
rect 27537 4573 27571 4607
rect 27571 4573 27580 4607
rect 53196 4632 53248 4684
rect 54300 4632 54352 4684
rect 27528 4564 27580 4573
rect 30288 4607 30340 4616
rect 30288 4573 30297 4607
rect 30297 4573 30331 4607
rect 30331 4573 30340 4607
rect 30288 4564 30340 4573
rect 30840 4564 30892 4616
rect 31116 4607 31168 4616
rect 31116 4573 31125 4607
rect 31125 4573 31159 4607
rect 31159 4573 31168 4607
rect 31116 4564 31168 4573
rect 32404 4564 32456 4616
rect 52092 4564 52144 4616
rect 52644 4564 52696 4616
rect 23940 4496 23992 4548
rect 24400 4471 24452 4480
rect 24400 4437 24409 4471
rect 24409 4437 24443 4471
rect 24443 4437 24452 4471
rect 24400 4428 24452 4437
rect 26884 4471 26936 4480
rect 26884 4437 26893 4471
rect 26893 4437 26927 4471
rect 26927 4437 26936 4471
rect 26884 4428 26936 4437
rect 30656 4471 30708 4480
rect 30656 4437 30665 4471
rect 30665 4437 30699 4471
rect 30699 4437 30708 4471
rect 30656 4428 30708 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 4712 4224 4764 4276
rect 6092 4224 6144 4276
rect 7932 4224 7984 4276
rect 8760 4267 8812 4276
rect 8760 4233 8769 4267
rect 8769 4233 8803 4267
rect 8803 4233 8812 4267
rect 8760 4224 8812 4233
rect 8944 4224 8996 4276
rect 9772 4267 9824 4276
rect 4896 4199 4948 4208
rect 4896 4165 4905 4199
rect 4905 4165 4939 4199
rect 4939 4165 4948 4199
rect 4896 4156 4948 4165
rect 5356 4156 5408 4208
rect 6368 4199 6420 4208
rect 6368 4165 6377 4199
rect 6377 4165 6411 4199
rect 6411 4165 6420 4199
rect 6368 4156 6420 4165
rect 2780 4131 2832 4140
rect 2780 4097 2789 4131
rect 2789 4097 2823 4131
rect 2823 4097 2832 4131
rect 2780 4088 2832 4097
rect 3148 4088 3200 4140
rect 4068 4131 4120 4140
rect 4068 4097 4077 4131
rect 4077 4097 4111 4131
rect 4111 4097 4120 4131
rect 4068 4088 4120 4097
rect 4344 4088 4396 4140
rect 5816 4131 5868 4140
rect 4528 4020 4580 4072
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 7288 4088 7340 4140
rect 7472 4088 7524 4140
rect 8208 4088 8260 4140
rect 8852 4088 8904 4140
rect 9772 4233 9781 4267
rect 9781 4233 9815 4267
rect 9815 4233 9824 4267
rect 9772 4224 9824 4233
rect 16396 4224 16448 4276
rect 22468 4224 22520 4276
rect 25872 4224 25924 4276
rect 29920 4267 29972 4276
rect 29920 4233 29929 4267
rect 29929 4233 29963 4267
rect 29963 4233 29972 4267
rect 29920 4224 29972 4233
rect 30840 4224 30892 4276
rect 5908 3952 5960 4004
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 2136 3884 2188 3893
rect 3792 3884 3844 3936
rect 4896 3884 4948 3936
rect 5448 3884 5500 3936
rect 6000 3884 6052 3936
rect 7840 4020 7892 4072
rect 8024 3952 8076 4004
rect 8760 4020 8812 4072
rect 9220 4088 9272 4140
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 11520 4131 11572 4140
rect 11520 4097 11529 4131
rect 11529 4097 11563 4131
rect 11563 4097 11572 4131
rect 11520 4088 11572 4097
rect 12716 4088 12768 4140
rect 14096 4088 14148 4140
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 13084 4020 13136 4072
rect 16028 4020 16080 4072
rect 16120 4020 16172 4072
rect 26424 4156 26476 4208
rect 19064 4088 19116 4140
rect 19524 4088 19576 4140
rect 20996 4088 21048 4140
rect 34796 4088 34848 4140
rect 35440 4088 35492 4140
rect 53012 4088 53064 4140
rect 6736 3927 6788 3936
rect 6736 3893 6745 3927
rect 6745 3893 6779 3927
rect 6779 3893 6788 3927
rect 6736 3884 6788 3893
rect 7564 3884 7616 3936
rect 8300 3927 8352 3936
rect 8300 3893 8309 3927
rect 8309 3893 8343 3927
rect 8343 3893 8352 3927
rect 8300 3884 8352 3893
rect 9220 3952 9272 4004
rect 11428 3952 11480 4004
rect 12624 3952 12676 4004
rect 13636 3952 13688 4004
rect 15200 3952 15252 4004
rect 16672 3952 16724 4004
rect 11244 3884 11296 3936
rect 14648 3884 14700 3936
rect 18420 3952 18472 4004
rect 26332 4020 26384 4072
rect 51816 4020 51868 4072
rect 54024 4020 54076 4072
rect 21548 3952 21600 4004
rect 52828 3952 52880 4004
rect 18512 3884 18564 3936
rect 18880 3884 18932 3936
rect 19432 3884 19484 3936
rect 20352 3884 20404 3936
rect 22928 3884 22980 3936
rect 23112 3884 23164 3936
rect 23388 3884 23440 3936
rect 24216 3884 24268 3936
rect 25320 3884 25372 3936
rect 35624 3884 35676 3936
rect 51080 3884 51132 3936
rect 51356 3884 51408 3936
rect 52460 3884 52512 3936
rect 55312 3927 55364 3936
rect 55312 3893 55321 3927
rect 55321 3893 55355 3927
rect 55355 3893 55364 3927
rect 55312 3884 55364 3893
rect 58440 3884 58492 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4068 3680 4120 3732
rect 4896 3680 4948 3732
rect 5724 3680 5776 3732
rect 5908 3723 5960 3732
rect 5908 3689 5917 3723
rect 5917 3689 5951 3723
rect 5951 3689 5960 3723
rect 5908 3680 5960 3689
rect 6092 3723 6144 3732
rect 6092 3689 6101 3723
rect 6101 3689 6135 3723
rect 6135 3689 6144 3723
rect 6092 3680 6144 3689
rect 8300 3723 8352 3732
rect 8300 3689 8309 3723
rect 8309 3689 8343 3723
rect 8343 3689 8352 3723
rect 8300 3680 8352 3689
rect 9128 3680 9180 3732
rect 9496 3680 9548 3732
rect 9588 3680 9640 3732
rect 14372 3680 14424 3732
rect 16120 3723 16172 3732
rect 16120 3689 16129 3723
rect 16129 3689 16163 3723
rect 16163 3689 16172 3723
rect 16120 3680 16172 3689
rect 17132 3680 17184 3732
rect 17776 3723 17828 3732
rect 17776 3689 17785 3723
rect 17785 3689 17819 3723
rect 17819 3689 17828 3723
rect 17776 3680 17828 3689
rect 18604 3723 18656 3732
rect 18604 3689 18613 3723
rect 18613 3689 18647 3723
rect 18647 3689 18656 3723
rect 18604 3680 18656 3689
rect 18788 3680 18840 3732
rect 27988 3723 28040 3732
rect 27988 3689 27997 3723
rect 27997 3689 28031 3723
rect 28031 3689 28040 3723
rect 27988 3680 28040 3689
rect 32404 3723 32456 3732
rect 32404 3689 32413 3723
rect 32413 3689 32447 3723
rect 32447 3689 32456 3723
rect 32404 3680 32456 3689
rect 52736 3680 52788 3732
rect 3424 3612 3476 3664
rect 3792 3612 3844 3664
rect 7564 3612 7616 3664
rect 8760 3612 8812 3664
rect 9036 3612 9088 3664
rect 16856 3612 16908 3664
rect 17960 3612 18012 3664
rect 20352 3655 20404 3664
rect 20352 3621 20361 3655
rect 20361 3621 20395 3655
rect 20395 3621 20404 3655
rect 20352 3612 20404 3621
rect 21364 3612 21416 3664
rect 26148 3612 26200 3664
rect 1860 3519 1912 3528
rect 1860 3485 1869 3519
rect 1869 3485 1903 3519
rect 1903 3485 1912 3519
rect 1860 3476 1912 3485
rect 2412 3476 2464 3528
rect 5448 3544 5500 3596
rect 6460 3544 6512 3596
rect 6828 3587 6880 3596
rect 6828 3553 6837 3587
rect 6837 3553 6871 3587
rect 6871 3553 6880 3587
rect 6828 3544 6880 3553
rect 5356 3476 5408 3528
rect 7748 3476 7800 3528
rect 8208 3476 8260 3528
rect 8668 3544 8720 3596
rect 12624 3544 12676 3596
rect 9404 3476 9456 3528
rect 9588 3476 9640 3528
rect 10324 3519 10376 3528
rect 10324 3485 10333 3519
rect 10333 3485 10367 3519
rect 10367 3485 10376 3519
rect 10324 3476 10376 3485
rect 10692 3476 10744 3528
rect 12532 3476 12584 3528
rect 13176 3476 13228 3528
rect 13912 3544 13964 3596
rect 15844 3544 15896 3596
rect 17500 3544 17552 3596
rect 14464 3476 14516 3528
rect 15752 3476 15804 3528
rect 16580 3476 16632 3528
rect 16856 3519 16908 3528
rect 16856 3485 16865 3519
rect 16865 3485 16899 3519
rect 16899 3485 16908 3519
rect 16856 3476 16908 3485
rect 21456 3544 21508 3596
rect 46296 3612 46348 3664
rect 51448 3612 51500 3664
rect 31024 3587 31076 3596
rect 31024 3553 31033 3587
rect 31033 3553 31067 3587
rect 31067 3553 31076 3587
rect 31024 3544 31076 3553
rect 50804 3544 50856 3596
rect 51632 3544 51684 3596
rect 53840 3544 53892 3596
rect 18328 3476 18380 3528
rect 20812 3476 20864 3528
rect 21640 3476 21692 3528
rect 23664 3476 23716 3528
rect 23940 3476 23992 3528
rect 24768 3476 24820 3528
rect 25596 3476 25648 3528
rect 26148 3519 26200 3528
rect 26148 3485 26157 3519
rect 26157 3485 26191 3519
rect 26191 3485 26200 3519
rect 26148 3476 26200 3485
rect 26884 3519 26936 3528
rect 26884 3485 26918 3519
rect 26918 3485 26936 3519
rect 26884 3476 26936 3485
rect 28632 3476 28684 3528
rect 30656 3476 30708 3528
rect 34704 3476 34756 3528
rect 35348 3476 35400 3528
rect 35808 3476 35860 3528
rect 36636 3476 36688 3528
rect 37464 3476 37516 3528
rect 38568 3476 38620 3528
rect 39948 3476 40000 3528
rect 40500 3476 40552 3528
rect 41052 3476 41104 3528
rect 42432 3476 42484 3528
rect 42708 3476 42760 3528
rect 44364 3476 44416 3528
rect 45192 3476 45244 3528
rect 46020 3476 46072 3528
rect 47676 3476 47728 3528
rect 48228 3476 48280 3528
rect 50160 3476 50212 3528
rect 50620 3476 50672 3528
rect 51172 3476 51224 3528
rect 52276 3476 52328 3528
rect 2136 3451 2188 3460
rect 2136 3417 2170 3451
rect 2170 3417 2188 3451
rect 2136 3408 2188 3417
rect 5264 3408 5316 3460
rect 5632 3408 5684 3460
rect 6552 3408 6604 3460
rect 8300 3408 8352 3460
rect 2780 3340 2832 3392
rect 4896 3340 4948 3392
rect 5908 3383 5960 3392
rect 5908 3349 5933 3383
rect 5933 3349 5960 3383
rect 5908 3340 5960 3349
rect 8576 3340 8628 3392
rect 9220 3340 9272 3392
rect 14832 3451 14884 3460
rect 14832 3417 14841 3451
rect 14841 3417 14875 3451
rect 14875 3417 14884 3451
rect 14832 3408 14884 3417
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 16672 3340 16724 3392
rect 16948 3340 17000 3392
rect 17776 3340 17828 3392
rect 19432 3340 19484 3392
rect 53288 3408 53340 3460
rect 57520 3519 57572 3528
rect 57520 3485 57529 3519
rect 57529 3485 57563 3519
rect 57563 3485 57572 3519
rect 57520 3476 57572 3485
rect 58164 3519 58216 3528
rect 58164 3485 58173 3519
rect 58173 3485 58207 3519
rect 58207 3485 58216 3519
rect 58164 3476 58216 3485
rect 20260 3340 20312 3392
rect 22836 3340 22888 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 1676 3136 1728 3188
rect 3516 3068 3568 3120
rect 3700 3136 3752 3188
rect 4068 3136 4120 3188
rect 4804 3136 4856 3188
rect 5908 3136 5960 3188
rect 8944 3179 8996 3188
rect 8944 3145 8953 3179
rect 8953 3145 8987 3179
rect 8987 3145 8996 3179
rect 8944 3136 8996 3145
rect 9128 3136 9180 3188
rect 14556 3179 14608 3188
rect 14556 3145 14565 3179
rect 14565 3145 14599 3179
rect 14599 3145 14608 3179
rect 14556 3136 14608 3145
rect 15292 3179 15344 3188
rect 15292 3145 15301 3179
rect 15301 3145 15335 3179
rect 15335 3145 15344 3179
rect 15292 3136 15344 3145
rect 16120 3136 16172 3188
rect 17684 3136 17736 3188
rect 18144 3179 18196 3188
rect 18144 3145 18153 3179
rect 18153 3145 18187 3179
rect 18187 3145 18196 3179
rect 18144 3136 18196 3145
rect 19432 3136 19484 3188
rect 20352 3179 20404 3188
rect 20352 3145 20361 3179
rect 20361 3145 20395 3179
rect 20395 3145 20404 3179
rect 20352 3136 20404 3145
rect 22284 3179 22336 3188
rect 22284 3145 22293 3179
rect 22293 3145 22327 3179
rect 22327 3145 22336 3179
rect 22284 3136 22336 3145
rect 23204 3136 23256 3188
rect 8760 3068 8812 3120
rect 8852 3068 8904 3120
rect 9220 3068 9272 3120
rect 11244 3068 11296 3120
rect 1768 3043 1820 3052
rect 1768 3009 1777 3043
rect 1777 3009 1811 3043
rect 1811 3009 1820 3043
rect 1768 3000 1820 3009
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 5080 3043 5132 3052
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 6736 3000 6788 3052
rect 7932 3000 7984 3052
rect 8024 3000 8076 3052
rect 10048 3000 10100 3052
rect 10416 3000 10468 3052
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 13452 3068 13504 3120
rect 11980 3000 12032 3052
rect 14004 3000 14056 3052
rect 17868 3068 17920 3120
rect 18604 3068 18656 3120
rect 18788 3111 18840 3120
rect 18788 3077 18797 3111
rect 18797 3077 18831 3111
rect 18831 3077 18840 3111
rect 18788 3068 18840 3077
rect 19064 3068 19116 3120
rect 20168 3068 20220 3120
rect 20536 3068 20588 3120
rect 20720 3068 20772 3120
rect 20996 3111 21048 3120
rect 20996 3077 21005 3111
rect 21005 3077 21039 3111
rect 21039 3077 21048 3111
rect 20996 3068 21048 3077
rect 21180 3111 21232 3120
rect 21180 3077 21189 3111
rect 21189 3077 21223 3111
rect 21223 3077 21232 3111
rect 21180 3068 21232 3077
rect 22100 3068 22152 3120
rect 24400 3068 24452 3120
rect 51908 3068 51960 3120
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 15292 3000 15344 3052
rect 16672 3000 16724 3052
rect 17224 3000 17276 3052
rect 17776 3000 17828 3052
rect 18512 3000 18564 3052
rect 3424 2932 3476 2984
rect 6000 2932 6052 2984
rect 6276 2932 6328 2984
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 6828 2932 6880 2941
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 7656 2932 7708 2984
rect 8944 2932 8996 2984
rect 17316 2932 17368 2984
rect 5448 2864 5500 2916
rect 3608 2796 3660 2848
rect 7380 2864 7432 2916
rect 9036 2864 9088 2916
rect 16488 2864 16540 2916
rect 19432 2864 19484 2916
rect 19984 3000 20036 3052
rect 22836 3043 22888 3052
rect 22836 3009 22845 3043
rect 22845 3009 22879 3043
rect 22879 3009 22888 3043
rect 22836 3000 22888 3009
rect 51724 3000 51776 3052
rect 54760 3000 54812 3052
rect 20260 2932 20312 2984
rect 20444 2932 20496 2984
rect 24492 2932 24544 2984
rect 26424 2932 26476 2984
rect 32772 2932 32824 2984
rect 38292 2932 38344 2984
rect 42156 2932 42208 2984
rect 53104 2932 53156 2984
rect 56600 2975 56652 2984
rect 56600 2941 56609 2975
rect 56609 2941 56643 2975
rect 56643 2941 56652 2975
rect 56600 2932 56652 2941
rect 23296 2864 23348 2916
rect 33324 2864 33376 2916
rect 34428 2864 34480 2916
rect 37188 2864 37240 2916
rect 39120 2864 39172 2916
rect 40224 2864 40276 2916
rect 42984 2864 43036 2916
rect 44088 2864 44140 2916
rect 8024 2796 8076 2848
rect 9496 2796 9548 2848
rect 9772 2796 9824 2848
rect 13176 2796 13228 2848
rect 15016 2796 15068 2848
rect 15108 2796 15160 2848
rect 15568 2796 15620 2848
rect 18880 2796 18932 2848
rect 20444 2796 20496 2848
rect 21272 2796 21324 2848
rect 21824 2796 21876 2848
rect 23480 2796 23532 2848
rect 25044 2796 25096 2848
rect 25872 2796 25924 2848
rect 26976 2796 27028 2848
rect 27804 2796 27856 2848
rect 28080 2839 28132 2848
rect 28080 2805 28089 2839
rect 28089 2805 28123 2839
rect 28123 2805 28132 2839
rect 28080 2796 28132 2805
rect 29184 2796 29236 2848
rect 29736 2796 29788 2848
rect 30012 2839 30064 2848
rect 30012 2805 30021 2839
rect 30021 2805 30055 2839
rect 30055 2805 30064 2839
rect 30012 2796 30064 2805
rect 30564 2796 30616 2848
rect 31668 2796 31720 2848
rect 32220 2796 32272 2848
rect 33876 2796 33928 2848
rect 35440 2796 35492 2848
rect 36360 2796 36412 2848
rect 37740 2796 37792 2848
rect 39672 2796 39724 2848
rect 41604 2796 41656 2848
rect 43536 2796 43588 2848
rect 44916 2796 44968 2848
rect 47400 2864 47452 2916
rect 48780 2864 48832 2916
rect 49884 2864 49936 2916
rect 50988 2864 51040 2916
rect 54208 2864 54260 2916
rect 45468 2796 45520 2848
rect 46848 2796 46900 2848
rect 47952 2796 48004 2848
rect 49332 2796 49384 2848
rect 50712 2796 50764 2848
rect 51540 2796 51592 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3976 2592 4028 2644
rect 5632 2592 5684 2644
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 10600 2592 10652 2644
rect 13452 2635 13504 2644
rect 13452 2601 13461 2635
rect 13461 2601 13495 2635
rect 13495 2601 13504 2635
rect 13452 2592 13504 2601
rect 14556 2635 14608 2644
rect 14556 2601 14565 2635
rect 14565 2601 14599 2635
rect 14599 2601 14608 2635
rect 14556 2592 14608 2601
rect 2964 2524 3016 2576
rect 7012 2524 7064 2576
rect 1584 2431 1636 2440
rect 1584 2397 1593 2431
rect 1593 2397 1627 2431
rect 1627 2397 1636 2431
rect 1584 2388 1636 2397
rect 3792 2456 3844 2508
rect 4068 2456 4120 2508
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 3884 2388 3936 2440
rect 4988 2456 5040 2508
rect 9220 2456 9272 2508
rect 2596 2320 2648 2372
rect 6276 2388 6328 2440
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 9404 2524 9456 2576
rect 13728 2524 13780 2576
rect 15844 2592 15896 2644
rect 17408 2635 17460 2644
rect 17408 2601 17417 2635
rect 17417 2601 17451 2635
rect 17451 2601 17460 2635
rect 17408 2592 17460 2601
rect 25412 2592 25464 2644
rect 29276 2592 29328 2644
rect 52000 2592 52052 2644
rect 14924 2456 14976 2508
rect 16212 2524 16264 2576
rect 18052 2567 18104 2576
rect 18052 2533 18061 2567
rect 18061 2533 18095 2567
rect 18095 2533 18104 2567
rect 18052 2524 18104 2533
rect 19156 2524 19208 2576
rect 20168 2524 20220 2576
rect 22468 2524 22520 2576
rect 22928 2524 22980 2576
rect 27252 2524 27304 2576
rect 28356 2524 28408 2576
rect 34152 2524 34204 2576
rect 38016 2524 38068 2576
rect 41880 2524 41932 2576
rect 45744 2524 45796 2576
rect 49608 2524 49660 2576
rect 11704 2388 11756 2440
rect 1768 2295 1820 2304
rect 1768 2261 1777 2295
rect 1777 2261 1811 2295
rect 1811 2261 1820 2295
rect 1768 2252 1820 2261
rect 7748 2320 7800 2372
rect 8484 2320 8536 2372
rect 10324 2320 10376 2372
rect 14004 2388 14056 2440
rect 14556 2388 14608 2440
rect 15476 2388 15528 2440
rect 15844 2388 15896 2440
rect 17868 2388 17920 2440
rect 19524 2388 19576 2440
rect 21272 2431 21324 2440
rect 21272 2397 21281 2431
rect 21281 2397 21315 2431
rect 21315 2397 21324 2431
rect 21272 2388 21324 2397
rect 22376 2388 22428 2440
rect 23020 2388 23072 2440
rect 23296 2388 23348 2440
rect 26240 2456 26292 2508
rect 26516 2456 26568 2508
rect 31944 2456 31996 2508
rect 33048 2456 33100 2508
rect 35532 2456 35584 2508
rect 38844 2456 38896 2508
rect 40776 2456 40828 2508
rect 43260 2456 43312 2508
rect 46572 2456 46624 2508
rect 48504 2456 48556 2508
rect 6736 2252 6788 2304
rect 17224 2320 17276 2372
rect 16028 2252 16080 2304
rect 20260 2320 20312 2372
rect 21548 2320 21600 2372
rect 27528 2388 27580 2440
rect 28908 2388 28960 2440
rect 29460 2388 29512 2440
rect 30288 2388 30340 2440
rect 30840 2388 30892 2440
rect 31116 2388 31168 2440
rect 31392 2388 31444 2440
rect 32496 2388 32548 2440
rect 33600 2388 33652 2440
rect 36084 2388 36136 2440
rect 26700 2320 26752 2372
rect 36912 2320 36964 2372
rect 39396 2388 39448 2440
rect 41328 2388 41380 2440
rect 43812 2388 43864 2440
rect 44640 2320 44692 2372
rect 47124 2388 47176 2440
rect 49056 2388 49108 2440
rect 50896 2388 50948 2440
rect 57888 2499 57940 2508
rect 52552 2388 52604 2440
rect 18512 2252 18564 2304
rect 22008 2295 22060 2304
rect 22008 2261 22017 2295
rect 22017 2261 22051 2295
rect 22051 2261 22060 2295
rect 22008 2252 22060 2261
rect 23020 2252 23072 2304
rect 51264 2252 51316 2304
rect 57888 2465 57897 2499
rect 57897 2465 57931 2499
rect 57931 2465 57940 2499
rect 57888 2456 57940 2465
rect 55956 2431 56008 2440
rect 55956 2397 55965 2431
rect 55965 2397 55999 2431
rect 55999 2397 56008 2431
rect 55956 2388 56008 2397
rect 56600 2431 56652 2440
rect 56600 2397 56609 2431
rect 56609 2397 56643 2431
rect 56643 2397 56652 2431
rect 56600 2388 56652 2397
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 7196 2048 7248 2100
rect 10324 2048 10376 2100
rect 10692 2048 10744 2100
rect 14004 2048 14056 2100
rect 1768 1912 1820 1964
rect 9496 1980 9548 2032
rect 10416 1980 10468 2032
rect 25412 2048 25464 2100
rect 26240 2048 26292 2100
rect 34612 2048 34664 2100
rect 52368 2048 52420 2100
rect 55956 2048 56008 2100
rect 14556 1980 14608 2032
rect 16396 1980 16448 2032
rect 22008 1980 22060 2032
rect 45560 1980 45612 2032
rect 53564 1980 53616 2032
rect 57888 1980 57940 2032
rect 6736 1912 6788 1964
rect 28816 1912 28868 1964
rect 5448 1844 5500 1896
rect 10692 1844 10744 1896
rect 15844 1844 15896 1896
rect 18052 1844 18104 1896
rect 1584 1708 1636 1760
rect 7196 1708 7248 1760
rect 8116 1708 8168 1760
rect 18512 1708 18564 1760
rect 18880 1708 18932 1760
rect 21088 1640 21140 1692
rect 21548 1640 21600 1692
rect 8116 1572 8168 1624
rect 20260 1572 20312 1624
rect 6000 1504 6052 1556
rect 6368 1504 6420 1556
rect 20352 1504 20404 1556
rect 20260 1436 20312 1488
rect 2964 1368 3016 1420
rect 8852 1368 8904 1420
rect 10600 1368 10652 1420
rect 19340 1300 19392 1352
rect 19800 1300 19852 1352
rect 19984 1300 20036 1352
rect 52736 1368 52788 1420
rect 53012 1368 53064 1420
rect 19432 1232 19484 1284
rect 6276 1164 6328 1216
rect 52552 1096 52604 1148
rect 19524 892 19576 944
rect 50988 892 51040 944
rect 52552 892 52604 944
rect 52920 892 52972 944
rect 56600 1368 56652 1420
rect 54760 824 54812 876
<< metal2 >>
rect 1766 59200 1822 60000
rect 3330 59200 3386 60000
rect 4894 59200 4950 60000
rect 6458 59200 6514 60000
rect 8022 59200 8078 60000
rect 9586 59200 9642 60000
rect 11150 59200 11206 60000
rect 12714 59200 12770 60000
rect 14278 59200 14334 60000
rect 15842 59200 15898 60000
rect 17406 59200 17462 60000
rect 18970 59200 19026 60000
rect 19076 59214 19288 59242
rect 1780 57594 1808 59200
rect 3344 57594 3372 59200
rect 4908 57594 4936 59200
rect 5264 57792 5316 57798
rect 5264 57734 5316 57740
rect 1768 57588 1820 57594
rect 1768 57530 1820 57536
rect 3332 57588 3384 57594
rect 3332 57530 3384 57536
rect 4896 57588 4948 57594
rect 4896 57530 4948 57536
rect 5276 57458 5304 57734
rect 6472 57594 6500 59200
rect 8036 57594 8064 59200
rect 6460 57588 6512 57594
rect 6460 57530 6512 57536
rect 8024 57588 8076 57594
rect 9600 57576 9628 59200
rect 11164 57594 11192 59200
rect 12728 57594 12756 59200
rect 14292 57594 14320 59200
rect 15856 57594 15884 59200
rect 17420 57594 17448 59200
rect 18984 59106 19012 59200
rect 19076 59106 19104 59214
rect 18984 59078 19104 59106
rect 18328 57792 18380 57798
rect 18328 57734 18380 57740
rect 9680 57588 9732 57594
rect 9600 57548 9680 57576
rect 8024 57530 8076 57536
rect 9680 57530 9732 57536
rect 11152 57588 11204 57594
rect 11152 57530 11204 57536
rect 12716 57588 12768 57594
rect 12716 57530 12768 57536
rect 14280 57588 14332 57594
rect 14280 57530 14332 57536
rect 15844 57588 15896 57594
rect 15844 57530 15896 57536
rect 17408 57588 17460 57594
rect 17408 57530 17460 57536
rect 2688 57452 2740 57458
rect 2688 57394 2740 57400
rect 4068 57452 4120 57458
rect 4068 57394 4120 57400
rect 5264 57452 5316 57458
rect 5264 57394 5316 57400
rect 11796 57452 11848 57458
rect 11796 57394 11848 57400
rect 13084 57452 13136 57458
rect 13084 57394 13136 57400
rect 15936 57452 15988 57458
rect 15936 57394 15988 57400
rect 16948 57452 17000 57458
rect 16948 57394 17000 57400
rect 17500 57452 17552 57458
rect 17500 57394 17552 57400
rect 2700 57254 2728 57394
rect 2688 57248 2740 57254
rect 2688 57190 2740 57196
rect 2700 56302 2728 57190
rect 2688 56296 2740 56302
rect 2688 56238 2740 56244
rect 4080 56234 4108 57394
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 11808 56982 11836 57394
rect 11796 56976 11848 56982
rect 11796 56918 11848 56924
rect 13096 56506 13124 57394
rect 15948 56506 15976 57394
rect 13084 56500 13136 56506
rect 13084 56442 13136 56448
rect 15936 56500 15988 56506
rect 15936 56442 15988 56448
rect 13728 56364 13780 56370
rect 13728 56306 13780 56312
rect 16212 56364 16264 56370
rect 16212 56306 16264 56312
rect 4068 56228 4120 56234
rect 4068 56170 4120 56176
rect 13740 56166 13768 56306
rect 13728 56160 13780 56166
rect 13728 56102 13780 56108
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 16224 55622 16252 56306
rect 16960 55962 16988 57394
rect 17512 56506 17540 57394
rect 17868 57248 17920 57254
rect 17868 57190 17920 57196
rect 17880 56506 17908 57190
rect 18340 57050 18368 57734
rect 19260 57610 19288 59214
rect 20534 59200 20590 60000
rect 22098 59200 22154 60000
rect 23662 59200 23718 60000
rect 25226 59200 25282 60000
rect 26790 59200 26846 60000
rect 28354 59200 28410 60000
rect 29918 59200 29974 60000
rect 31482 59200 31538 60000
rect 33046 59200 33102 60000
rect 34610 59200 34666 60000
rect 36174 59200 36230 60000
rect 37738 59200 37794 60000
rect 39302 59200 39358 60000
rect 40866 59200 40922 60000
rect 42430 59200 42486 60000
rect 43994 59200 44050 60000
rect 45558 59200 45614 60000
rect 47122 59200 47178 60000
rect 48686 59200 48742 60000
rect 50250 59200 50306 60000
rect 51814 59200 51870 60000
rect 53378 59200 53434 60000
rect 54942 59200 54998 60000
rect 56506 59200 56562 60000
rect 58070 59200 58126 60000
rect 58438 59256 58494 59265
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 20548 57610 20576 59200
rect 19260 57594 19380 57610
rect 20548 57594 20760 57610
rect 22112 57594 22140 59200
rect 23676 57594 23704 59200
rect 25240 57594 25268 59200
rect 26804 57594 26832 59200
rect 28368 57594 28396 59200
rect 29932 57594 29960 59200
rect 31496 57594 31524 59200
rect 19260 57588 19392 57594
rect 19260 57582 19340 57588
rect 20548 57588 20772 57594
rect 20548 57582 20720 57588
rect 19340 57530 19392 57536
rect 20720 57530 20772 57536
rect 22100 57588 22152 57594
rect 22100 57530 22152 57536
rect 23664 57588 23716 57594
rect 23664 57530 23716 57536
rect 25228 57588 25280 57594
rect 25228 57530 25280 57536
rect 26792 57588 26844 57594
rect 26792 57530 26844 57536
rect 28356 57588 28408 57594
rect 28356 57530 28408 57536
rect 29920 57588 29972 57594
rect 29920 57530 29972 57536
rect 31484 57588 31536 57594
rect 33060 57576 33088 59200
rect 34624 57594 34652 59200
rect 36188 57594 36216 59200
rect 37752 57594 37780 59200
rect 39316 57594 39344 59200
rect 40880 57594 40908 59200
rect 42444 57594 42472 59200
rect 33140 57588 33192 57594
rect 33060 57548 33140 57576
rect 31484 57530 31536 57536
rect 33140 57530 33192 57536
rect 34612 57588 34664 57594
rect 34612 57530 34664 57536
rect 36176 57588 36228 57594
rect 36176 57530 36228 57536
rect 37740 57588 37792 57594
rect 37740 57530 37792 57536
rect 39304 57588 39356 57594
rect 39304 57530 39356 57536
rect 40868 57588 40920 57594
rect 40868 57530 40920 57536
rect 42432 57588 42484 57594
rect 44008 57576 44036 59200
rect 45572 57594 45600 59200
rect 47136 57594 47164 59200
rect 44180 57588 44232 57594
rect 44008 57548 44180 57576
rect 42432 57530 42484 57536
rect 44180 57530 44232 57536
rect 45560 57588 45612 57594
rect 45560 57530 45612 57536
rect 47124 57588 47176 57594
rect 47124 57530 47176 57536
rect 19156 57520 19208 57526
rect 19156 57462 19208 57468
rect 18420 57316 18472 57322
rect 18420 57258 18472 57264
rect 18328 57044 18380 57050
rect 18328 56986 18380 56992
rect 18052 56704 18104 56710
rect 18052 56646 18104 56652
rect 17500 56500 17552 56506
rect 17500 56442 17552 56448
rect 17868 56500 17920 56506
rect 17868 56442 17920 56448
rect 18064 56370 18092 56646
rect 18432 56506 18460 57258
rect 18512 57248 18564 57254
rect 18512 57190 18564 57196
rect 18524 56846 18552 57190
rect 19168 57050 19196 57462
rect 48700 57458 48728 59200
rect 50264 57882 50292 59200
rect 50172 57854 50292 57882
rect 50172 57458 50200 57854
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 51828 57458 51856 59200
rect 53392 57458 53420 59200
rect 19248 57452 19300 57458
rect 19248 57394 19300 57400
rect 19340 57452 19392 57458
rect 19340 57394 19392 57400
rect 22192 57452 22244 57458
rect 22192 57394 22244 57400
rect 24400 57452 24452 57458
rect 24400 57394 24452 57400
rect 25320 57452 25372 57458
rect 25320 57394 25372 57400
rect 26976 57452 27028 57458
rect 26976 57394 27028 57400
rect 28448 57452 28500 57458
rect 28448 57394 28500 57400
rect 30012 57452 30064 57458
rect 30012 57394 30064 57400
rect 33232 57452 33284 57458
rect 33232 57394 33284 57400
rect 34796 57452 34848 57458
rect 34796 57394 34848 57400
rect 37832 57452 37884 57458
rect 37832 57394 37884 57400
rect 37924 57452 37976 57458
rect 37924 57394 37976 57400
rect 40960 57452 41012 57458
rect 40960 57394 41012 57400
rect 42340 57452 42392 57458
rect 42340 57394 42392 57400
rect 44088 57452 44140 57458
rect 44088 57394 44140 57400
rect 45652 57452 45704 57458
rect 45652 57394 45704 57400
rect 47584 57452 47636 57458
rect 47584 57394 47636 57400
rect 48688 57452 48740 57458
rect 48688 57394 48740 57400
rect 50160 57452 50212 57458
rect 50160 57394 50212 57400
rect 51816 57452 51868 57458
rect 51816 57394 51868 57400
rect 53380 57452 53432 57458
rect 53380 57394 53432 57400
rect 19156 57044 19208 57050
rect 19156 56986 19208 56992
rect 18512 56840 18564 56846
rect 18510 56808 18512 56817
rect 18564 56808 18566 56817
rect 18510 56743 18566 56752
rect 18420 56500 18472 56506
rect 18420 56442 18472 56448
rect 18880 56432 18932 56438
rect 18880 56374 18932 56380
rect 17408 56364 17460 56370
rect 17408 56306 17460 56312
rect 18052 56364 18104 56370
rect 18052 56306 18104 56312
rect 18696 56364 18748 56370
rect 18696 56306 18748 56312
rect 16948 55956 17000 55962
rect 16948 55898 17000 55904
rect 17316 55820 17368 55826
rect 17316 55762 17368 55768
rect 17132 55752 17184 55758
rect 17132 55694 17184 55700
rect 16212 55616 16264 55622
rect 16210 55584 16212 55593
rect 16264 55584 16266 55593
rect 16210 55519 16266 55528
rect 17144 55350 17172 55694
rect 17132 55344 17184 55350
rect 17130 55312 17132 55321
rect 17184 55312 17186 55321
rect 17130 55247 17186 55256
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 15292 47592 15344 47598
rect 15292 47534 15344 47540
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 12808 42288 12860 42294
rect 12808 42230 12860 42236
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 12164 41540 12216 41546
rect 12164 41482 12216 41488
rect 10416 41268 10468 41274
rect 10416 41210 10468 41216
rect 11796 41268 11848 41274
rect 11796 41210 11848 41216
rect 9864 41132 9916 41138
rect 9864 41074 9916 41080
rect 9680 40996 9732 41002
rect 9680 40938 9732 40944
rect 8300 40928 8352 40934
rect 8300 40870 8352 40876
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 5264 40520 5316 40526
rect 5316 40468 5488 40474
rect 5264 40462 5488 40468
rect 5276 40446 5488 40462
rect 4988 40180 5040 40186
rect 4988 40122 5040 40128
rect 3792 40044 3844 40050
rect 3792 39986 3844 39992
rect 4804 40044 4856 40050
rect 4804 39986 4856 39992
rect 2504 39976 2556 39982
rect 2504 39918 2556 39924
rect 1952 38752 2004 38758
rect 1952 38694 2004 38700
rect 1964 38282 1992 38694
rect 1952 38276 2004 38282
rect 1952 38218 2004 38224
rect 1768 38208 1820 38214
rect 1768 38150 1820 38156
rect 1780 37942 1808 38150
rect 1768 37936 1820 37942
rect 1768 37878 1820 37884
rect 1964 29102 1992 38218
rect 2516 37874 2544 39918
rect 3804 39642 3832 39986
rect 4620 39840 4672 39846
rect 4620 39782 4672 39788
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4632 39642 4660 39782
rect 3792 39636 3844 39642
rect 3792 39578 3844 39584
rect 4620 39636 4672 39642
rect 4620 39578 4672 39584
rect 4160 38956 4212 38962
rect 4160 38898 4212 38904
rect 3976 38752 4028 38758
rect 4172 38740 4200 38898
rect 4620 38888 4672 38894
rect 4620 38830 4672 38836
rect 3976 38694 4028 38700
rect 4080 38712 4200 38740
rect 3988 38418 4016 38694
rect 4080 38434 4108 38712
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 3976 38412 4028 38418
rect 4080 38406 4200 38434
rect 3976 38354 4028 38360
rect 2872 38344 2924 38350
rect 2872 38286 2924 38292
rect 2688 38208 2740 38214
rect 2688 38150 2740 38156
rect 2700 37874 2728 38150
rect 2504 37868 2556 37874
rect 2504 37810 2556 37816
rect 2688 37868 2740 37874
rect 2688 37810 2740 37816
rect 2516 36174 2544 37810
rect 2504 36168 2556 36174
rect 2504 36110 2556 36116
rect 2516 34610 2544 36110
rect 2504 34604 2556 34610
rect 2504 34546 2556 34552
rect 2780 34604 2832 34610
rect 2780 34546 2832 34552
rect 2792 34202 2820 34546
rect 2780 34196 2832 34202
rect 2780 34138 2832 34144
rect 2884 33998 2912 38286
rect 4172 38010 4200 38406
rect 4436 38412 4488 38418
rect 4436 38354 4488 38360
rect 4448 38214 4476 38354
rect 4632 38214 4660 38830
rect 4816 38554 4844 39986
rect 5000 39438 5028 40122
rect 5264 39840 5316 39846
rect 5264 39782 5316 39788
rect 4988 39432 5040 39438
rect 4988 39374 5040 39380
rect 5000 38876 5028 39374
rect 5276 39302 5304 39782
rect 5356 39568 5408 39574
rect 5356 39510 5408 39516
rect 5264 39296 5316 39302
rect 5264 39238 5316 39244
rect 5080 38888 5132 38894
rect 5000 38848 5080 38876
rect 5080 38830 5132 38836
rect 4804 38548 4856 38554
rect 4804 38490 4856 38496
rect 4436 38208 4488 38214
rect 4436 38150 4488 38156
rect 4620 38208 4672 38214
rect 4620 38150 4672 38156
rect 4160 38004 4212 38010
rect 4160 37946 4212 37952
rect 4448 37806 4476 38150
rect 4436 37800 4488 37806
rect 4436 37742 4488 37748
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37262 4660 38150
rect 4816 37942 4844 38490
rect 5092 38350 5120 38830
rect 5080 38344 5132 38350
rect 5080 38286 5132 38292
rect 4804 37936 4856 37942
rect 4804 37878 4856 37884
rect 5092 37874 5120 38286
rect 5080 37868 5132 37874
rect 5080 37810 5132 37816
rect 4804 37800 4856 37806
rect 4724 37760 4804 37788
rect 4724 37670 4752 37760
rect 4804 37742 4856 37748
rect 4712 37664 4764 37670
rect 4712 37606 4764 37612
rect 4620 37256 4672 37262
rect 4620 37198 4672 37204
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36174 4660 37198
rect 4620 36168 4672 36174
rect 4620 36110 4672 36116
rect 4620 36032 4672 36038
rect 4620 35974 4672 35980
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 35290 4660 35974
rect 4620 35284 4672 35290
rect 4620 35226 4672 35232
rect 3240 35148 3292 35154
rect 3240 35090 3292 35096
rect 3148 34400 3200 34406
rect 3148 34342 3200 34348
rect 3160 33998 3188 34342
rect 2872 33992 2924 33998
rect 2872 33934 2924 33940
rect 3148 33992 3200 33998
rect 3148 33934 3200 33940
rect 2228 33448 2280 33454
rect 2228 33390 2280 33396
rect 2240 32434 2268 33390
rect 2228 32428 2280 32434
rect 2228 32370 2280 32376
rect 2320 32428 2372 32434
rect 2320 32370 2372 32376
rect 2240 30258 2268 32370
rect 2332 32026 2360 32370
rect 2320 32020 2372 32026
rect 2320 31962 2372 31968
rect 2688 31816 2740 31822
rect 2688 31758 2740 31764
rect 2596 30592 2648 30598
rect 2596 30534 2648 30540
rect 2228 30252 2280 30258
rect 2228 30194 2280 30200
rect 2504 30252 2556 30258
rect 2504 30194 2556 30200
rect 2516 29850 2544 30194
rect 2504 29844 2556 29850
rect 2504 29786 2556 29792
rect 2608 29782 2636 30534
rect 2596 29776 2648 29782
rect 2596 29718 2648 29724
rect 2320 29640 2372 29646
rect 2700 29628 2728 31758
rect 2884 31754 2912 33934
rect 3252 31958 3280 35090
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4068 33992 4120 33998
rect 4344 33992 4396 33998
rect 4120 33940 4200 33946
rect 4068 33934 4200 33940
rect 4344 33934 4396 33940
rect 4080 33918 4200 33934
rect 4172 33862 4200 33918
rect 3792 33856 3844 33862
rect 3792 33798 3844 33804
rect 4068 33856 4120 33862
rect 4068 33798 4120 33804
rect 4160 33856 4212 33862
rect 4160 33798 4212 33804
rect 3804 33522 3832 33798
rect 3792 33516 3844 33522
rect 3792 33458 3844 33464
rect 4080 32774 4108 33798
rect 4356 33658 4384 33934
rect 4344 33652 4396 33658
rect 4344 33594 4396 33600
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4068 32768 4120 32774
rect 4068 32710 4120 32716
rect 3608 32224 3660 32230
rect 3608 32166 3660 32172
rect 3240 31952 3292 31958
rect 3240 31894 3292 31900
rect 2780 31748 2832 31754
rect 2884 31726 3096 31754
rect 2780 31690 2832 31696
rect 2792 31482 2820 31690
rect 2780 31476 2832 31482
rect 2780 31418 2832 31424
rect 2780 31340 2832 31346
rect 2780 31282 2832 31288
rect 2792 30666 2820 31282
rect 2780 30660 2832 30666
rect 2780 30602 2832 30608
rect 2780 29640 2832 29646
rect 2700 29600 2780 29628
rect 2320 29582 2372 29588
rect 2780 29582 2832 29588
rect 1952 29096 2004 29102
rect 1952 29038 2004 29044
rect 2332 28762 2360 29582
rect 2964 29164 3016 29170
rect 2964 29106 3016 29112
rect 2780 28960 2832 28966
rect 2780 28902 2832 28908
rect 2320 28756 2372 28762
rect 2320 28698 2372 28704
rect 2792 28150 2820 28902
rect 2872 28756 2924 28762
rect 2872 28698 2924 28704
rect 2780 28144 2832 28150
rect 2780 28086 2832 28092
rect 2412 28008 2464 28014
rect 2412 27950 2464 27956
rect 2424 25838 2452 27950
rect 2504 27328 2556 27334
rect 2504 27270 2556 27276
rect 2516 26994 2544 27270
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 2412 25832 2464 25838
rect 2412 25774 2464 25780
rect 2424 25294 2452 25774
rect 2412 25288 2464 25294
rect 2412 25230 2464 25236
rect 2424 24750 2452 25230
rect 2412 24744 2464 24750
rect 2412 24686 2464 24692
rect 2228 23724 2280 23730
rect 2228 23666 2280 23672
rect 1584 23044 1636 23050
rect 1584 22986 1636 22992
rect 1596 22778 1624 22986
rect 1584 22772 1636 22778
rect 1584 22714 1636 22720
rect 2240 22574 2268 23666
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2332 22710 2360 22918
rect 2320 22704 2372 22710
rect 2320 22646 2372 22652
rect 2424 22642 2452 24686
rect 2412 22636 2464 22642
rect 2412 22578 2464 22584
rect 2228 22568 2280 22574
rect 2228 22510 2280 22516
rect 2136 21956 2188 21962
rect 2136 21898 2188 21904
rect 2148 21690 2176 21898
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 2516 21350 2544 26930
rect 2780 26784 2832 26790
rect 2780 26726 2832 26732
rect 2792 24818 2820 26726
rect 2884 26382 2912 28698
rect 2976 28422 3004 29106
rect 2964 28416 3016 28422
rect 2964 28358 3016 28364
rect 2872 26376 2924 26382
rect 2924 26324 3004 26330
rect 2872 26318 3004 26324
rect 2884 26302 3004 26318
rect 2872 26240 2924 26246
rect 2872 26182 2924 26188
rect 2884 25974 2912 26182
rect 2872 25968 2924 25974
rect 2872 25910 2924 25916
rect 2780 24812 2832 24818
rect 2780 24754 2832 24760
rect 2596 23520 2648 23526
rect 2596 23462 2648 23468
rect 2608 21554 2636 23462
rect 2976 23254 3004 26302
rect 2964 23248 3016 23254
rect 2964 23190 3016 23196
rect 2688 23112 2740 23118
rect 2688 23054 2740 23060
rect 2700 21570 2728 23054
rect 2872 22024 2924 22030
rect 2872 21966 2924 21972
rect 2780 21616 2832 21622
rect 2700 21564 2780 21570
rect 2700 21558 2832 21564
rect 2596 21548 2648 21554
rect 2700 21542 2820 21558
rect 2596 21490 2648 21496
rect 2504 21344 2556 21350
rect 2504 21286 2556 21292
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2412 19712 2464 19718
rect 2412 19654 2464 19660
rect 2424 18698 2452 19654
rect 2412 18692 2464 18698
rect 2412 18634 2464 18640
rect 2608 18426 2636 19790
rect 2884 19242 2912 21966
rect 3068 20534 3096 31726
rect 3252 29578 3280 31894
rect 3332 31680 3384 31686
rect 3332 31622 3384 31628
rect 3240 29572 3292 29578
rect 3240 29514 3292 29520
rect 3148 29164 3200 29170
rect 3252 29152 3280 29514
rect 3200 29124 3280 29152
rect 3148 29106 3200 29112
rect 3344 27334 3372 31622
rect 3620 31414 3648 32166
rect 4080 31414 4108 32710
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3608 31408 3660 31414
rect 3608 31350 3660 31356
rect 4068 31408 4120 31414
rect 4068 31350 4120 31356
rect 3516 30048 3568 30054
rect 3516 29990 3568 29996
rect 3424 29640 3476 29646
rect 3424 29582 3476 29588
rect 3436 29170 3464 29582
rect 3528 29238 3556 29990
rect 3620 29646 3648 31350
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3792 30728 3844 30734
rect 3792 30670 3844 30676
rect 3804 30122 3832 30670
rect 3792 30116 3844 30122
rect 3792 30058 3844 30064
rect 3608 29640 3660 29646
rect 3608 29582 3660 29588
rect 3516 29232 3568 29238
rect 3516 29174 3568 29180
rect 3804 29170 3832 30058
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4724 29714 4752 37606
rect 5172 36780 5224 36786
rect 5172 36722 5224 36728
rect 5184 36378 5212 36722
rect 5172 36372 5224 36378
rect 5172 36314 5224 36320
rect 5184 35766 5212 36314
rect 5172 35760 5224 35766
rect 5172 35702 5224 35708
rect 4896 35692 4948 35698
rect 4896 35634 4948 35640
rect 4804 35488 4856 35494
rect 4804 35430 4856 35436
rect 4816 35086 4844 35430
rect 4804 35080 4856 35086
rect 4804 35022 4856 35028
rect 4908 30666 4936 35634
rect 4988 35080 5040 35086
rect 4988 35022 5040 35028
rect 5000 34474 5028 35022
rect 5080 34672 5132 34678
rect 5080 34614 5132 34620
rect 4988 34468 5040 34474
rect 4988 34410 5040 34416
rect 5000 31822 5028 34410
rect 4988 31816 5040 31822
rect 4988 31758 5040 31764
rect 4896 30660 4948 30666
rect 4896 30602 4948 30608
rect 4908 30326 4936 30602
rect 4896 30320 4948 30326
rect 4896 30262 4948 30268
rect 4712 29708 4764 29714
rect 4712 29650 4764 29656
rect 4344 29572 4396 29578
rect 4344 29514 4396 29520
rect 4356 29238 4384 29514
rect 4896 29504 4948 29510
rect 4896 29446 4948 29452
rect 4344 29232 4396 29238
rect 4344 29174 4396 29180
rect 3424 29164 3476 29170
rect 3424 29106 3476 29112
rect 3792 29164 3844 29170
rect 3792 29106 3844 29112
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3976 27396 4028 27402
rect 3976 27338 4028 27344
rect 3332 27328 3384 27334
rect 3332 27270 3384 27276
rect 3148 27124 3200 27130
rect 3148 27066 3200 27072
rect 3160 26246 3188 27066
rect 3240 26988 3292 26994
rect 3240 26930 3292 26936
rect 3884 26988 3936 26994
rect 3884 26930 3936 26936
rect 3252 26382 3280 26930
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3148 26240 3200 26246
rect 3148 26182 3200 26188
rect 3608 26240 3660 26246
rect 3608 26182 3660 26188
rect 3620 25838 3648 26182
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3896 24954 3924 26930
rect 3988 26518 4016 27338
rect 4068 26988 4120 26994
rect 4068 26930 4120 26936
rect 3976 26512 4028 26518
rect 3976 26454 4028 26460
rect 3988 26042 4016 26454
rect 4080 26382 4108 26930
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4068 26376 4120 26382
rect 4632 26353 4660 28358
rect 4908 26994 4936 29446
rect 4988 29028 5040 29034
rect 4988 28970 5040 28976
rect 5000 27470 5028 28970
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 5092 27130 5120 34614
rect 5276 31482 5304 39238
rect 5368 38418 5396 39510
rect 5460 39506 5488 40446
rect 5632 40452 5684 40458
rect 5632 40394 5684 40400
rect 6460 40452 6512 40458
rect 6460 40394 6512 40400
rect 5540 40112 5592 40118
rect 5540 40054 5592 40060
rect 5448 39500 5500 39506
rect 5448 39442 5500 39448
rect 5460 39030 5488 39442
rect 5448 39024 5500 39030
rect 5448 38966 5500 38972
rect 5356 38412 5408 38418
rect 5356 38354 5408 38360
rect 5356 38276 5408 38282
rect 5356 38218 5408 38224
rect 5368 38010 5396 38218
rect 5356 38004 5408 38010
rect 5356 37946 5408 37952
rect 5356 33448 5408 33454
rect 5356 33390 5408 33396
rect 5264 31476 5316 31482
rect 5264 31418 5316 31424
rect 5276 31385 5304 31418
rect 5262 31376 5318 31385
rect 5262 31311 5318 31320
rect 5264 30252 5316 30258
rect 5264 30194 5316 30200
rect 5276 29170 5304 30194
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 5276 28218 5304 29106
rect 5264 28212 5316 28218
rect 5264 28154 5316 28160
rect 5368 27470 5396 33390
rect 5552 29238 5580 40054
rect 5644 39642 5672 40394
rect 6472 40050 6500 40394
rect 6552 40384 6604 40390
rect 6552 40326 6604 40332
rect 7564 40384 7616 40390
rect 7564 40326 7616 40332
rect 6460 40044 6512 40050
rect 6460 39986 6512 39992
rect 5816 39908 5868 39914
rect 5816 39850 5868 39856
rect 5632 39636 5684 39642
rect 5632 39578 5684 39584
rect 5828 39438 5856 39850
rect 6368 39840 6420 39846
rect 6368 39782 6420 39788
rect 6380 39438 6408 39782
rect 5816 39432 5868 39438
rect 5816 39374 5868 39380
rect 6368 39432 6420 39438
rect 6368 39374 6420 39380
rect 6276 39364 6328 39370
rect 6276 39306 6328 39312
rect 6288 38554 6316 39306
rect 6276 38548 6328 38554
rect 6276 38490 6328 38496
rect 6564 38350 6592 40326
rect 6828 40044 6880 40050
rect 6828 39986 6880 39992
rect 6644 39908 6696 39914
rect 6644 39850 6696 39856
rect 6736 39908 6788 39914
rect 6736 39850 6788 39856
rect 6552 38344 6604 38350
rect 6552 38286 6604 38292
rect 5908 38276 5960 38282
rect 5908 38218 5960 38224
rect 5920 37738 5948 38218
rect 5724 37732 5776 37738
rect 5724 37674 5776 37680
rect 5908 37732 5960 37738
rect 5908 37674 5960 37680
rect 5736 37330 5764 37674
rect 5724 37324 5776 37330
rect 5724 37266 5776 37272
rect 5632 35012 5684 35018
rect 5632 34954 5684 34960
rect 5644 34610 5672 34954
rect 5632 34604 5684 34610
rect 5632 34546 5684 34552
rect 5644 33522 5672 34546
rect 5736 33862 5764 37266
rect 6564 36854 6592 38286
rect 6656 37890 6684 39850
rect 6748 39642 6776 39850
rect 6736 39636 6788 39642
rect 6736 39578 6788 39584
rect 6840 39098 6868 39986
rect 7104 39296 7156 39302
rect 7104 39238 7156 39244
rect 6828 39092 6880 39098
rect 6828 39034 6880 39040
rect 7116 39030 7144 39238
rect 7104 39024 7156 39030
rect 7104 38966 7156 38972
rect 6828 38888 6880 38894
rect 6828 38830 6880 38836
rect 6840 38298 6868 38830
rect 6748 38282 6868 38298
rect 6736 38276 6868 38282
rect 6788 38270 6868 38276
rect 6736 38218 6788 38224
rect 6748 38010 6776 38218
rect 6736 38004 6788 38010
rect 6736 37946 6788 37952
rect 6656 37862 6776 37890
rect 6552 36848 6604 36854
rect 6552 36790 6604 36796
rect 6552 36032 6604 36038
rect 6552 35974 6604 35980
rect 6092 34944 6144 34950
rect 6092 34886 6144 34892
rect 5724 33856 5776 33862
rect 5724 33798 5776 33804
rect 5632 33516 5684 33522
rect 5632 33458 5684 33464
rect 5644 31754 5672 33458
rect 5632 31748 5684 31754
rect 5632 31690 5684 31696
rect 5644 31482 5672 31690
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 5644 30734 5672 31418
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 5632 29640 5684 29646
rect 5632 29582 5684 29588
rect 5540 29232 5592 29238
rect 5540 29174 5592 29180
rect 5644 29170 5672 29582
rect 5632 29164 5684 29170
rect 5632 29106 5684 29112
rect 5644 28694 5672 29106
rect 5632 28688 5684 28694
rect 5632 28630 5684 28636
rect 5356 27464 5408 27470
rect 5356 27406 5408 27412
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 5172 27396 5224 27402
rect 5172 27338 5224 27344
rect 5080 27124 5132 27130
rect 5080 27066 5132 27072
rect 5184 26994 5212 27338
rect 5460 26994 5488 27406
rect 5632 27328 5684 27334
rect 5632 27270 5684 27276
rect 4896 26988 4948 26994
rect 4896 26930 4948 26936
rect 5172 26988 5224 26994
rect 5172 26930 5224 26936
rect 5448 26988 5500 26994
rect 5448 26930 5500 26936
rect 4068 26318 4120 26324
rect 4618 26344 4674 26353
rect 4618 26279 4674 26288
rect 5078 26344 5134 26353
rect 5644 26314 5672 27270
rect 5078 26279 5134 26288
rect 5632 26308 5684 26314
rect 3976 26036 4028 26042
rect 3976 25978 4028 25984
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 3884 24948 3936 24954
rect 3884 24890 3936 24896
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 3252 22234 3280 23666
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 3792 23180 3844 23186
rect 3792 23122 3844 23128
rect 3804 22982 3832 23122
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3700 21956 3752 21962
rect 3700 21898 3752 21904
rect 3712 21690 3740 21898
rect 3700 21684 3752 21690
rect 3700 21626 3752 21632
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 3056 20528 3108 20534
rect 3056 20470 3108 20476
rect 3252 19990 3280 21286
rect 3240 19984 3292 19990
rect 3240 19926 3292 19932
rect 2872 19236 2924 19242
rect 2872 19178 2924 19184
rect 2884 18766 2912 19178
rect 3804 18902 3832 22918
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4160 21956 4212 21962
rect 4160 21898 4212 21904
rect 3976 21548 4028 21554
rect 4172 21536 4200 21898
rect 4632 21622 4660 22374
rect 5092 21962 5120 26279
rect 5632 26250 5684 26256
rect 5736 24818 5764 33798
rect 5908 31272 5960 31278
rect 5908 31214 5960 31220
rect 5920 30938 5948 31214
rect 5908 30932 5960 30938
rect 5908 30874 5960 30880
rect 6104 25974 6132 34886
rect 6368 33584 6420 33590
rect 6368 33526 6420 33532
rect 6380 32434 6408 33526
rect 6564 32774 6592 35974
rect 6644 35488 6696 35494
rect 6644 35430 6696 35436
rect 6656 35018 6684 35430
rect 6644 35012 6696 35018
rect 6644 34954 6696 34960
rect 6656 34746 6684 34954
rect 6644 34740 6696 34746
rect 6644 34682 6696 34688
rect 6552 32768 6604 32774
rect 6552 32710 6604 32716
rect 6368 32428 6420 32434
rect 6368 32370 6420 32376
rect 6460 32428 6512 32434
rect 6460 32370 6512 32376
rect 6380 32026 6408 32370
rect 6368 32020 6420 32026
rect 6368 31962 6420 31968
rect 6276 30660 6328 30666
rect 6276 30602 6328 30608
rect 6288 30138 6316 30602
rect 6380 30326 6408 31962
rect 6472 30938 6500 32370
rect 6460 30932 6512 30938
rect 6460 30874 6512 30880
rect 6368 30320 6420 30326
rect 6368 30262 6420 30268
rect 6288 30110 6408 30138
rect 6380 30054 6408 30110
rect 6368 30048 6420 30054
rect 6368 29990 6420 29996
rect 6380 28150 6408 29990
rect 6368 28144 6420 28150
rect 6368 28086 6420 28092
rect 6564 26874 6592 32710
rect 6748 32230 6776 37862
rect 7012 37188 7064 37194
rect 7012 37130 7064 37136
rect 7024 36378 7052 37130
rect 7196 36576 7248 36582
rect 7196 36518 7248 36524
rect 7472 36576 7524 36582
rect 7472 36518 7524 36524
rect 7012 36372 7064 36378
rect 7012 36314 7064 36320
rect 6828 34944 6880 34950
rect 6828 34886 6880 34892
rect 6840 34134 6868 34886
rect 6828 34128 6880 34134
rect 6828 34070 6880 34076
rect 6736 32224 6788 32230
rect 6736 32166 6788 32172
rect 6748 31754 6776 32166
rect 6656 31726 6776 31754
rect 6656 30734 6684 31726
rect 6840 31414 6868 34070
rect 6920 33516 6972 33522
rect 6920 33458 6972 33464
rect 6932 33114 6960 33458
rect 6920 33108 6972 33114
rect 6920 33050 6972 33056
rect 6828 31408 6880 31414
rect 6828 31350 6880 31356
rect 6840 30870 6868 31350
rect 7104 31340 7156 31346
rect 7104 31282 7156 31288
rect 6828 30864 6880 30870
rect 6828 30806 6880 30812
rect 7116 30734 7144 31282
rect 6644 30728 6696 30734
rect 6644 30670 6696 30676
rect 7104 30728 7156 30734
rect 7104 30670 7156 30676
rect 6920 30660 6972 30666
rect 6920 30602 6972 30608
rect 6828 30320 6880 30326
rect 6828 30262 6880 30268
rect 6840 29170 6868 30262
rect 6932 29510 6960 30602
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6828 29164 6880 29170
rect 6828 29106 6880 29112
rect 6644 28960 6696 28966
rect 6644 28902 6696 28908
rect 6656 28082 6684 28902
rect 6644 28076 6696 28082
rect 6644 28018 6696 28024
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 6920 28076 6972 28082
rect 6920 28018 6972 28024
rect 6748 27470 6776 28018
rect 6736 27464 6788 27470
rect 6736 27406 6788 27412
rect 6748 27130 6776 27406
rect 6932 27402 6960 28018
rect 6920 27396 6972 27402
rect 6920 27338 6972 27344
rect 6736 27124 6788 27130
rect 6736 27066 6788 27072
rect 6736 26988 6788 26994
rect 6736 26930 6788 26936
rect 6564 26846 6684 26874
rect 6184 26308 6236 26314
rect 6184 26250 6236 26256
rect 6092 25968 6144 25974
rect 6092 25910 6144 25916
rect 6196 25498 6224 26250
rect 6276 26240 6328 26246
rect 6552 26240 6604 26246
rect 6328 26188 6408 26194
rect 6276 26182 6408 26188
rect 6552 26182 6604 26188
rect 6288 26166 6408 26182
rect 6380 26042 6408 26166
rect 6368 26036 6420 26042
rect 6368 25978 6420 25984
rect 6380 25906 6408 25978
rect 6564 25906 6592 26182
rect 6368 25900 6420 25906
rect 6368 25842 6420 25848
rect 6552 25900 6604 25906
rect 6552 25842 6604 25848
rect 6184 25492 6236 25498
rect 6184 25434 6236 25440
rect 6368 25288 6420 25294
rect 6368 25230 6420 25236
rect 5908 25220 5960 25226
rect 5908 25162 5960 25168
rect 5920 24954 5948 25162
rect 5908 24948 5960 24954
rect 5908 24890 5960 24896
rect 5724 24812 5776 24818
rect 5724 24754 5776 24760
rect 6000 22772 6052 22778
rect 6000 22714 6052 22720
rect 5172 22704 5224 22710
rect 5172 22646 5224 22652
rect 5080 21956 5132 21962
rect 5080 21898 5132 21904
rect 5092 21622 5120 21898
rect 5184 21894 5212 22646
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 5184 21622 5212 21830
rect 4620 21616 4672 21622
rect 4620 21558 4672 21564
rect 5080 21616 5132 21622
rect 5080 21558 5132 21564
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 4028 21508 4200 21536
rect 3976 21490 4028 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4804 20460 4856 20466
rect 4804 20402 4856 20408
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4816 19854 4844 20402
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3792 18896 3844 18902
rect 3792 18838 3844 18844
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2228 18148 2280 18154
rect 2228 18090 2280 18096
rect 2240 15502 2268 18090
rect 2884 17202 2912 18702
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 3804 18358 3832 18566
rect 3792 18352 3844 18358
rect 3792 18294 3844 18300
rect 4540 18170 4568 18566
rect 4632 18426 4660 19314
rect 4816 19258 4844 19790
rect 4724 19230 4844 19258
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 4724 18766 4752 19230
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4540 18142 4660 18170
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3712 17270 3740 18022
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 16114 2360 16390
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2516 15706 2544 16526
rect 2884 16182 2912 17138
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 2872 16176 2924 16182
rect 2872 16118 2924 16124
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 3896 15502 3924 15846
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 2148 14550 2176 14962
rect 2240 14958 2268 15438
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2228 14952 2280 14958
rect 2228 14894 2280 14900
rect 2688 14952 2740 14958
rect 2688 14894 2740 14900
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2608 14414 2636 14758
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2700 14074 2728 14894
rect 2884 14618 2912 14962
rect 3792 14816 3844 14822
rect 3792 14758 3844 14764
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2688 14068 2740 14074
rect 2688 14010 2740 14016
rect 2700 12782 2728 14010
rect 3804 13870 3832 14758
rect 3792 13864 3844 13870
rect 3792 13806 3844 13812
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2148 11762 2176 12582
rect 2884 12238 2912 12718
rect 3804 12306 3832 13806
rect 3988 12434 4016 16458
rect 3896 12406 4016 12434
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2884 10062 2912 12174
rect 3804 11830 3832 12242
rect 3792 11824 3844 11830
rect 3792 11766 3844 11772
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9586 1716 9862
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1596 2446 1624 8774
rect 1688 8498 1716 8774
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1872 8430 1900 9454
rect 2884 9042 2912 9998
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1688 3194 1716 3878
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1780 3058 1808 7686
rect 1872 5710 1900 8366
rect 2332 8090 2360 8910
rect 3896 8838 3924 12406
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3988 9042 4016 9318
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2044 6112 2096 6118
rect 2044 6054 2096 6060
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 1860 5704 1912 5710
rect 1860 5646 1912 5652
rect 1872 3534 1900 5646
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 2056 3233 2084 6054
rect 2148 5710 2176 6054
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2516 5370 2544 6258
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2148 3466 2176 3878
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2136 3460 2188 3466
rect 2136 3402 2188 3408
rect 2042 3224 2098 3233
rect 2042 3159 2098 3168
rect 2424 3058 2452 3470
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 1780 2961 1808 2994
rect 1766 2952 1822 2961
rect 1766 2887 1822 2896
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1596 1766 1624 2382
rect 2608 2378 2636 7142
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2700 5234 2728 5578
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2792 4146 2820 8774
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2884 7954 2912 8230
rect 2962 7984 3018 7993
rect 2872 7948 2924 7954
rect 2962 7919 3018 7928
rect 2872 7890 2924 7896
rect 2976 7886 3004 7919
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 3068 4622 3096 6666
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 3160 4146 3188 7142
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3252 5710 3280 6598
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3344 4622 3372 6734
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 2792 3398 2820 4082
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 3160 3097 3188 4082
rect 3252 3641 3280 4422
rect 3238 3632 3294 3641
rect 3238 3567 3294 3576
rect 3344 3516 3372 4558
rect 3436 3670 3464 7414
rect 3700 7404 3752 7410
rect 3700 7346 3752 7352
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3344 3488 3464 3516
rect 3146 3088 3202 3097
rect 3146 3023 3202 3032
rect 3436 2990 3464 3488
rect 3528 3126 3556 7142
rect 3606 4176 3662 4185
rect 3606 4111 3662 4120
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 3620 2854 3648 4111
rect 3712 3194 3740 7346
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6390 3832 6598
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3790 4040 3846 4049
rect 3790 3975 3846 3984
rect 3804 3942 3832 3975
rect 3792 3936 3844 3942
rect 3792 3878 3844 3884
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3700 3188 3752 3194
rect 3700 3130 3752 3136
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3238 2680 3294 2689
rect 3238 2615 3294 2624
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 1780 1970 1808 2246
rect 1768 1964 1820 1970
rect 1768 1906 1820 1912
rect 1584 1760 1636 1766
rect 1584 1702 1636 1708
rect 2976 1426 3004 2518
rect 3252 2446 3280 2615
rect 3804 2514 3832 3606
rect 3792 2508 3844 2514
rect 3792 2450 3844 2456
rect 3896 2446 3924 8774
rect 3976 8288 4028 8294
rect 3976 8230 4028 8236
rect 3988 7993 4016 8230
rect 3974 7984 4030 7993
rect 3974 7919 4030 7928
rect 3976 7744 4028 7750
rect 3976 7686 4028 7692
rect 3988 7410 4016 7686
rect 4080 7410 4108 17818
rect 4632 17338 4660 18142
rect 4724 17814 4752 18702
rect 4816 18222 4844 19110
rect 4908 18834 4936 19246
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4712 17808 4764 17814
rect 4712 17750 4764 17756
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4724 17134 4752 17478
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4356 16250 4384 16526
rect 4724 16454 4752 17070
rect 4712 16448 4764 16454
rect 4712 16390 4764 16396
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4712 16040 4764 16046
rect 4908 16028 4936 18770
rect 5092 18154 5120 21558
rect 6012 20942 6040 22714
rect 6380 22642 6408 25230
rect 6368 22636 6420 22642
rect 6368 22578 6420 22584
rect 6368 22432 6420 22438
rect 6368 22374 6420 22380
rect 6092 22092 6144 22098
rect 6092 22034 6144 22040
rect 6104 21690 6132 22034
rect 6380 22030 6408 22374
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6552 22024 6604 22030
rect 6656 22012 6684 26846
rect 6748 26382 6776 26930
rect 6828 26784 6880 26790
rect 6828 26726 6880 26732
rect 6736 26376 6788 26382
rect 6736 26318 6788 26324
rect 6736 25900 6788 25906
rect 6736 25842 6788 25848
rect 6604 21984 6684 22012
rect 6552 21966 6604 21972
rect 6092 21684 6144 21690
rect 6092 21626 6144 21632
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6196 20942 6224 21626
rect 6656 21078 6684 21984
rect 6748 21894 6776 25842
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6644 21072 6696 21078
rect 6644 21014 6696 21020
rect 6000 20936 6052 20942
rect 6000 20878 6052 20884
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5908 19712 5960 19718
rect 5908 19654 5960 19660
rect 5644 19514 5672 19654
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5920 19446 5948 19654
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5276 18970 5304 19314
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 5080 18148 5132 18154
rect 5080 18090 5132 18096
rect 5276 17814 5304 18906
rect 5356 18692 5408 18698
rect 5356 18634 5408 18640
rect 5368 18086 5396 18634
rect 5920 18290 5948 19382
rect 6012 18698 6040 19722
rect 6656 18970 6684 21014
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 6000 18692 6052 18698
rect 6000 18634 6052 18640
rect 6184 18692 6236 18698
rect 6184 18634 6236 18640
rect 5908 18284 5960 18290
rect 5908 18226 5960 18232
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 4988 17808 5040 17814
rect 4988 17750 5040 17756
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 4764 16000 4936 16028
rect 4712 15982 4764 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 12782 4660 13874
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12170 4660 12718
rect 4724 12714 4752 15982
rect 5000 14906 5028 17750
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5080 15428 5132 15434
rect 5080 15370 5132 15376
rect 4816 14878 5028 14906
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 8906 4660 10610
rect 4724 9110 4752 12650
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4632 8566 4660 8842
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7818 4660 8502
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6866 4016 7142
rect 4080 7002 4108 7346
rect 4264 7206 4292 7346
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 3988 5234 4016 6802
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4540 6662 4568 6734
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 4528 5160 4580 5166
rect 4526 5128 4528 5137
rect 4580 5128 4582 5137
rect 4526 5063 4582 5072
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4826 4660 6734
rect 4724 5778 4752 9046
rect 4816 5846 4844 14878
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 4896 14544 4948 14550
rect 4896 14486 4948 14492
rect 4908 11665 4936 14486
rect 5000 14482 5028 14758
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4894 11656 4950 11665
rect 4894 11591 4950 11600
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 10606 4936 11494
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5000 8430 5028 8910
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 5000 7818 5028 8366
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 4896 7268 4948 7274
rect 4896 7210 4948 7216
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4712 5160 4764 5166
rect 4712 5102 4764 5108
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4724 4622 4752 5102
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 3988 2650 4016 4490
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4356 4146 4384 4422
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4080 3738 4108 4082
rect 4540 4078 4568 4422
rect 4724 4282 4752 4558
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4816 3194 4844 5170
rect 4908 4214 4936 7210
rect 5000 5574 5028 7754
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5000 5370 5028 5510
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 5000 4729 5028 5170
rect 4986 4720 5042 4729
rect 4986 4655 5042 4664
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3738 4936 3878
rect 4896 3732 4948 3738
rect 4896 3674 4948 3680
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4080 2514 4108 3130
rect 4908 2825 4936 3334
rect 4894 2816 4950 2825
rect 4214 2748 4522 2757
rect 4894 2751 4950 2760
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5000 2514 5028 4655
rect 5092 3058 5120 15370
rect 5276 14958 5304 16390
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 5276 11694 5304 14894
rect 5368 12850 5396 18022
rect 5460 17882 5488 18158
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5644 17134 5672 17614
rect 5920 17542 5948 18226
rect 6196 18086 6224 18634
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 18290 6776 18566
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5644 16726 5672 17070
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5644 15026 5672 16662
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5368 12306 5396 12786
rect 5448 12776 5500 12782
rect 5448 12718 5500 12724
rect 5356 12300 5408 12306
rect 5356 12242 5408 12248
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5276 9042 5304 11630
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 5184 6662 5212 8434
rect 5368 8242 5396 12242
rect 5460 11558 5488 12718
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5552 11762 5580 12038
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5644 11218 5672 14962
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5828 14618 5856 14758
rect 5816 14612 5868 14618
rect 5816 14554 5868 14560
rect 5816 14272 5868 14278
rect 5814 14240 5816 14249
rect 5868 14240 5870 14249
rect 5814 14175 5870 14184
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5632 10532 5684 10538
rect 5632 10474 5684 10480
rect 5644 10130 5672 10474
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5460 9586 5488 9862
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5552 8294 5580 9590
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5540 8288 5592 8294
rect 5368 8214 5488 8242
rect 5540 8230 5592 8236
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5368 7342 5396 8026
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 4622 5212 6598
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5276 3466 5304 7210
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5368 5234 5396 6258
rect 5460 5574 5488 8214
rect 5552 7954 5580 8230
rect 5540 7948 5592 7954
rect 5540 7890 5592 7896
rect 5644 7886 5672 9454
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5920 7342 5948 17478
rect 6196 16250 6224 18022
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6184 16244 6236 16250
rect 6184 16186 6236 16192
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6368 15020 6420 15026
rect 6368 14962 6420 14968
rect 6000 14476 6052 14482
rect 6000 14418 6052 14424
rect 6012 12714 6040 14418
rect 6380 13938 6408 14962
rect 6368 13932 6420 13938
rect 6196 13892 6368 13920
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 6012 10538 6040 12650
rect 6196 12238 6224 13892
rect 6368 13874 6420 13880
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6380 12442 6408 12582
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6276 12368 6328 12374
rect 6276 12310 6328 12316
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6196 11830 6224 12174
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 6196 10062 6224 11086
rect 6288 10810 6316 12310
rect 6472 12238 6500 15574
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6564 15026 6592 15302
rect 6656 15026 6684 16934
rect 6748 15434 6776 18226
rect 6840 15706 6868 26726
rect 6932 26518 6960 27338
rect 7208 26994 7236 36518
rect 7484 36174 7512 36518
rect 7380 36168 7432 36174
rect 7380 36110 7432 36116
rect 7472 36168 7524 36174
rect 7472 36110 7524 36116
rect 7392 35222 7420 36110
rect 7472 35692 7524 35698
rect 7472 35634 7524 35640
rect 7484 35290 7512 35634
rect 7472 35284 7524 35290
rect 7472 35226 7524 35232
rect 7380 35216 7432 35222
rect 7380 35158 7432 35164
rect 7392 34202 7420 35158
rect 7576 35086 7604 40326
rect 7748 40044 7800 40050
rect 8312 40032 8340 40870
rect 7800 40004 8340 40032
rect 7748 39986 7800 39992
rect 8852 39840 8904 39846
rect 8852 39782 8904 39788
rect 8116 39296 8168 39302
rect 8116 39238 8168 39244
rect 8128 37262 8156 39238
rect 8392 39092 8444 39098
rect 8392 39034 8444 39040
rect 8404 38350 8432 39034
rect 8864 38350 8892 39782
rect 9692 38486 9720 40938
rect 9876 40934 9904 41074
rect 9864 40928 9916 40934
rect 9864 40870 9916 40876
rect 9864 40520 9916 40526
rect 9864 40462 9916 40468
rect 9876 40118 9904 40462
rect 9864 40112 9916 40118
rect 9864 40054 9916 40060
rect 9876 39438 9904 40054
rect 9864 39432 9916 39438
rect 9864 39374 9916 39380
rect 9876 38758 9904 39374
rect 10048 39364 10100 39370
rect 10048 39306 10100 39312
rect 9864 38752 9916 38758
rect 9864 38694 9916 38700
rect 9680 38480 9732 38486
rect 9680 38422 9732 38428
rect 8392 38344 8444 38350
rect 8392 38286 8444 38292
rect 8852 38344 8904 38350
rect 8852 38286 8904 38292
rect 9404 38344 9456 38350
rect 9404 38286 9456 38292
rect 7840 37256 7892 37262
rect 7840 37198 7892 37204
rect 8116 37256 8168 37262
rect 8116 37198 8168 37204
rect 8208 37256 8260 37262
rect 8208 37198 8260 37204
rect 7852 36854 7880 37198
rect 7932 37188 7984 37194
rect 7932 37130 7984 37136
rect 7840 36848 7892 36854
rect 7840 36790 7892 36796
rect 7944 36718 7972 37130
rect 8220 36854 8248 37198
rect 8300 37120 8352 37126
rect 8300 37062 8352 37068
rect 8208 36848 8260 36854
rect 8208 36790 8260 36796
rect 8024 36780 8076 36786
rect 8024 36722 8076 36728
rect 7932 36712 7984 36718
rect 7932 36654 7984 36660
rect 8036 35630 8064 36722
rect 8024 35624 8076 35630
rect 8024 35566 8076 35572
rect 7564 35080 7616 35086
rect 7564 35022 7616 35028
rect 7576 34542 7604 35022
rect 8312 34678 8340 37062
rect 8300 34672 8352 34678
rect 8300 34614 8352 34620
rect 8208 34604 8260 34610
rect 8208 34546 8260 34552
rect 7564 34536 7616 34542
rect 7564 34478 7616 34484
rect 7748 34536 7800 34542
rect 7748 34478 7800 34484
rect 7380 34196 7432 34202
rect 7380 34138 7432 34144
rect 7472 32904 7524 32910
rect 7472 32846 7524 32852
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 7288 32020 7340 32026
rect 7288 31962 7340 31968
rect 7300 31822 7328 31962
rect 7288 31816 7340 31822
rect 7288 31758 7340 31764
rect 7300 31482 7328 31758
rect 7288 31476 7340 31482
rect 7288 31418 7340 31424
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 6920 26512 6972 26518
rect 6920 26454 6972 26460
rect 7012 25696 7064 25702
rect 7012 25638 7064 25644
rect 7024 25294 7052 25638
rect 7012 25288 7064 25294
rect 7012 25230 7064 25236
rect 7300 25226 7328 31418
rect 7392 27402 7420 32710
rect 7484 32570 7512 32846
rect 7472 32564 7524 32570
rect 7472 32506 7524 32512
rect 7564 31816 7616 31822
rect 7564 31758 7616 31764
rect 7470 31376 7526 31385
rect 7470 31311 7472 31320
rect 7524 31311 7526 31320
rect 7472 31282 7524 31288
rect 7576 30802 7604 31758
rect 7656 31136 7708 31142
rect 7656 31078 7708 31084
rect 7564 30796 7616 30802
rect 7564 30738 7616 30744
rect 7668 30258 7696 31078
rect 7656 30252 7708 30258
rect 7656 30194 7708 30200
rect 7760 29578 7788 34478
rect 8220 33658 8248 34546
rect 8208 33652 8260 33658
rect 8208 33594 8260 33600
rect 7932 32972 7984 32978
rect 7932 32914 7984 32920
rect 7944 30938 7972 32914
rect 8220 32910 8248 33594
rect 8208 32904 8260 32910
rect 8208 32846 8260 32852
rect 8208 32768 8260 32774
rect 8208 32710 8260 32716
rect 8220 32434 8248 32710
rect 8208 32428 8260 32434
rect 8208 32370 8260 32376
rect 8116 32224 8168 32230
rect 8116 32166 8168 32172
rect 8128 31754 8156 32166
rect 8116 31748 8168 31754
rect 8116 31690 8168 31696
rect 7932 30932 7984 30938
rect 7932 30874 7984 30880
rect 7748 29572 7800 29578
rect 7748 29514 7800 29520
rect 7472 28076 7524 28082
rect 7472 28018 7524 28024
rect 7484 27538 7512 28018
rect 7748 27600 7800 27606
rect 7748 27542 7800 27548
rect 7472 27532 7524 27538
rect 7472 27474 7524 27480
rect 7484 27402 7512 27474
rect 7380 27396 7432 27402
rect 7380 27338 7432 27344
rect 7472 27396 7524 27402
rect 7472 27338 7524 27344
rect 7392 26586 7420 27338
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 7484 26382 7512 27338
rect 7656 26512 7708 26518
rect 7656 26454 7708 26460
rect 7472 26376 7524 26382
rect 7472 26318 7524 26324
rect 7288 25220 7340 25226
rect 7288 25162 7340 25168
rect 7300 24954 7328 25162
rect 7288 24948 7340 24954
rect 7288 24890 7340 24896
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7208 24682 7236 24754
rect 7196 24676 7248 24682
rect 7196 24618 7248 24624
rect 7012 23656 7064 23662
rect 7012 23598 7064 23604
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6932 22098 6960 22578
rect 6920 22092 6972 22098
rect 6920 22034 6972 22040
rect 7024 22030 7052 23598
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 6920 21956 6972 21962
rect 6920 21898 6972 21904
rect 6932 21554 6960 21898
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 7208 20058 7236 24618
rect 7288 23112 7340 23118
rect 7288 23054 7340 23060
rect 7300 22030 7328 23054
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7472 22024 7524 22030
rect 7472 21966 7524 21972
rect 7484 21146 7512 21966
rect 7472 21140 7524 21146
rect 7472 21082 7524 21088
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 6920 18692 6972 18698
rect 6920 18634 6972 18640
rect 6932 18358 6960 18634
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 7484 18290 7512 19110
rect 7196 18284 7248 18290
rect 7481 18284 7533 18290
rect 7248 18244 7328 18272
rect 7196 18226 7248 18232
rect 7300 18204 7328 18244
rect 7481 18226 7533 18232
rect 7300 18176 7420 18204
rect 7196 16992 7248 16998
rect 7196 16934 7248 16940
rect 7208 16522 7236 16934
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7300 16590 7328 16730
rect 7392 16726 7420 18176
rect 7380 16720 7432 16726
rect 7380 16662 7432 16668
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 7116 15570 7144 15846
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6748 14550 6776 15030
rect 7392 14958 7420 16662
rect 7472 16584 7524 16590
rect 7576 16574 7604 19450
rect 7668 19242 7696 26454
rect 7760 22094 7788 27542
rect 7944 27130 7972 30874
rect 8024 29504 8076 29510
rect 8024 29446 8076 29452
rect 7932 27124 7984 27130
rect 7852 27084 7932 27112
rect 7852 25838 7880 27084
rect 7932 27066 7984 27072
rect 7932 26988 7984 26994
rect 7932 26930 7984 26936
rect 7944 26382 7972 26930
rect 7932 26376 7984 26382
rect 7930 26344 7932 26353
rect 7984 26344 7986 26353
rect 7930 26279 7986 26288
rect 7840 25832 7892 25838
rect 7840 25774 7892 25780
rect 7840 24132 7892 24138
rect 7840 24074 7892 24080
rect 7852 23730 7880 24074
rect 7840 23724 7892 23730
rect 7840 23666 7892 23672
rect 8036 22094 8064 29446
rect 8128 26314 8156 31690
rect 8404 29238 8432 38286
rect 9416 37874 9444 38286
rect 9496 38208 9548 38214
rect 9496 38150 9548 38156
rect 9404 37868 9456 37874
rect 9404 37810 9456 37816
rect 9508 36378 9536 38150
rect 9496 36372 9548 36378
rect 9496 36314 9548 36320
rect 9876 36174 9904 38694
rect 10060 38554 10088 39306
rect 10048 38548 10100 38554
rect 10048 38490 10100 38496
rect 10428 38486 10456 41210
rect 10968 41132 11020 41138
rect 10968 41074 11020 41080
rect 10980 40050 11008 41074
rect 11428 40928 11480 40934
rect 11428 40870 11480 40876
rect 11440 40526 11468 40870
rect 11428 40520 11480 40526
rect 11428 40462 11480 40468
rect 11336 40180 11388 40186
rect 11336 40122 11388 40128
rect 10968 40044 11020 40050
rect 10968 39986 11020 39992
rect 10416 38480 10468 38486
rect 10416 38422 10468 38428
rect 10232 38344 10284 38350
rect 10232 38286 10284 38292
rect 10244 38010 10272 38286
rect 10232 38004 10284 38010
rect 10232 37946 10284 37952
rect 9956 36780 10008 36786
rect 9956 36722 10008 36728
rect 8944 36168 8996 36174
rect 8944 36110 8996 36116
rect 9864 36168 9916 36174
rect 9864 36110 9916 36116
rect 8956 35630 8984 36110
rect 9772 35828 9824 35834
rect 9772 35770 9824 35776
rect 8944 35624 8996 35630
rect 8944 35566 8996 35572
rect 8484 34740 8536 34746
rect 8484 34682 8536 34688
rect 8852 34740 8904 34746
rect 8852 34682 8904 34688
rect 8496 34610 8524 34682
rect 8484 34604 8536 34610
rect 8484 34546 8536 34552
rect 8576 31272 8628 31278
rect 8576 31214 8628 31220
rect 8392 29232 8444 29238
rect 8392 29174 8444 29180
rect 8404 28626 8432 29174
rect 8392 28620 8444 28626
rect 8392 28562 8444 28568
rect 8300 28552 8352 28558
rect 8300 28494 8352 28500
rect 8482 28520 8538 28529
rect 8312 27538 8340 28494
rect 8482 28455 8538 28464
rect 8496 28218 8524 28455
rect 8484 28212 8536 28218
rect 8484 28154 8536 28160
rect 8300 27532 8352 27538
rect 8300 27474 8352 27480
rect 8116 26308 8168 26314
rect 8116 26250 8168 26256
rect 8208 26308 8260 26314
rect 8208 26250 8260 26256
rect 8220 26042 8248 26250
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8588 25498 8616 31214
rect 8668 27328 8720 27334
rect 8668 27270 8720 27276
rect 8680 26994 8708 27270
rect 8668 26988 8720 26994
rect 8668 26930 8720 26936
rect 8576 25492 8628 25498
rect 8576 25434 8628 25440
rect 8588 25294 8616 25434
rect 8576 25288 8628 25294
rect 8496 25248 8576 25276
rect 8116 22568 8168 22574
rect 8116 22510 8168 22516
rect 8128 22234 8156 22510
rect 8392 22432 8444 22438
rect 8392 22374 8444 22380
rect 8116 22228 8168 22234
rect 8116 22170 8168 22176
rect 7760 22066 7880 22094
rect 8036 22066 8156 22094
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7760 16794 7788 18158
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7524 16546 7604 16574
rect 7472 16526 7524 16532
rect 7564 15564 7616 15570
rect 7564 15506 7616 15512
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 7116 14414 7144 14758
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 12322 6868 12718
rect 6564 12294 6868 12322
rect 7392 12306 7420 14894
rect 7576 13841 7604 15506
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7668 13977 7696 15438
rect 7760 15314 7788 16730
rect 7852 15706 7880 22066
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7944 21622 7972 21830
rect 7932 21616 7984 21622
rect 7932 21558 7984 21564
rect 8128 21418 8156 22066
rect 8404 22030 8432 22374
rect 8496 22094 8524 25248
rect 8576 25230 8628 25236
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 8588 23730 8616 25094
rect 8576 23724 8628 23730
rect 8576 23666 8628 23672
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8680 22234 8708 22578
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8496 22066 8616 22094
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 8312 21622 8340 21898
rect 8300 21616 8352 21622
rect 8352 21576 8524 21604
rect 8300 21558 8352 21564
rect 8300 21480 8352 21486
rect 8300 21422 8352 21428
rect 8116 21412 8168 21418
rect 8116 21354 8168 21360
rect 8128 21078 8156 21354
rect 8116 21072 8168 21078
rect 8116 21014 8168 21020
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 7944 19446 7972 20198
rect 8312 19854 8340 21422
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8404 20262 8432 20810
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8300 19848 8352 19854
rect 8300 19790 8352 19796
rect 7932 19440 7984 19446
rect 7932 19382 7984 19388
rect 7944 18290 7972 19382
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 8128 18737 8156 19246
rect 8312 18834 8340 19790
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 19310 8432 19654
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8114 18728 8170 18737
rect 8114 18663 8170 18672
rect 8496 18358 8524 21576
rect 8588 19446 8616 22066
rect 8576 19440 8628 19446
rect 8576 19382 8628 19388
rect 8864 19174 8892 34682
rect 8956 32502 8984 35566
rect 9588 35080 9640 35086
rect 9588 35022 9640 35028
rect 9600 33930 9628 35022
rect 9680 34604 9732 34610
rect 9680 34546 9732 34552
rect 9692 34134 9720 34546
rect 9680 34128 9732 34134
rect 9680 34070 9732 34076
rect 9588 33924 9640 33930
rect 9588 33866 9640 33872
rect 8944 32496 8996 32502
rect 8944 32438 8996 32444
rect 8956 29850 8984 32438
rect 9600 31278 9628 33866
rect 9784 32570 9812 35770
rect 9876 35698 9904 36110
rect 9968 35698 9996 36722
rect 10324 36100 10376 36106
rect 10324 36042 10376 36048
rect 10140 36032 10192 36038
rect 10140 35974 10192 35980
rect 10152 35698 10180 35974
rect 9864 35692 9916 35698
rect 9864 35634 9916 35640
rect 9956 35692 10008 35698
rect 9956 35634 10008 35640
rect 10140 35692 10192 35698
rect 10140 35634 10192 35640
rect 9968 34610 9996 35634
rect 10336 34746 10364 36042
rect 10428 35154 10456 38422
rect 10980 38350 11008 39986
rect 11348 39370 11376 40122
rect 11808 40050 11836 41210
rect 12176 40730 12204 41482
rect 12532 41472 12584 41478
rect 12532 41414 12584 41420
rect 12624 41472 12676 41478
rect 12624 41414 12676 41420
rect 12544 41206 12572 41414
rect 12532 41200 12584 41206
rect 12532 41142 12584 41148
rect 12164 40724 12216 40730
rect 12164 40666 12216 40672
rect 11796 40044 11848 40050
rect 11796 39986 11848 39992
rect 11520 39908 11572 39914
rect 11520 39850 11572 39856
rect 11796 39908 11848 39914
rect 11796 39850 11848 39856
rect 11532 39642 11560 39850
rect 11520 39636 11572 39642
rect 11520 39578 11572 39584
rect 11152 39364 11204 39370
rect 11152 39306 11204 39312
rect 11336 39364 11388 39370
rect 11336 39306 11388 39312
rect 10968 38344 11020 38350
rect 10968 38286 11020 38292
rect 10784 38004 10836 38010
rect 10784 37946 10836 37952
rect 10796 37670 10824 37946
rect 10784 37664 10836 37670
rect 10784 37606 10836 37612
rect 10980 35698 11008 38286
rect 11164 38282 11192 39306
rect 11244 39296 11296 39302
rect 11244 39238 11296 39244
rect 11256 38350 11284 39238
rect 11808 38758 11836 39850
rect 11980 39364 12032 39370
rect 11980 39306 12032 39312
rect 11796 38752 11848 38758
rect 11796 38694 11848 38700
rect 11244 38344 11296 38350
rect 11244 38286 11296 38292
rect 11152 38276 11204 38282
rect 11152 38218 11204 38224
rect 11520 38276 11572 38282
rect 11520 38218 11572 38224
rect 11428 36372 11480 36378
rect 11428 36314 11480 36320
rect 11336 36032 11388 36038
rect 11336 35974 11388 35980
rect 11060 35760 11112 35766
rect 11060 35702 11112 35708
rect 10784 35692 10836 35698
rect 10784 35634 10836 35640
rect 10968 35692 11020 35698
rect 10968 35634 11020 35640
rect 10416 35148 10468 35154
rect 10416 35090 10468 35096
rect 10692 35148 10744 35154
rect 10692 35090 10744 35096
rect 10704 34746 10732 35090
rect 10796 35086 10824 35634
rect 10968 35488 11020 35494
rect 10968 35430 11020 35436
rect 10980 35086 11008 35430
rect 10784 35080 10836 35086
rect 10784 35022 10836 35028
rect 10968 35080 11020 35086
rect 10968 35022 11020 35028
rect 10968 34944 11020 34950
rect 10968 34886 11020 34892
rect 10324 34740 10376 34746
rect 10324 34682 10376 34688
rect 10692 34740 10744 34746
rect 10692 34682 10744 34688
rect 10416 34672 10468 34678
rect 10416 34614 10468 34620
rect 9956 34604 10008 34610
rect 9956 34546 10008 34552
rect 10232 34604 10284 34610
rect 10232 34546 10284 34552
rect 9864 34400 9916 34406
rect 9864 34342 9916 34348
rect 9772 32564 9824 32570
rect 9772 32506 9824 32512
rect 9680 31748 9732 31754
rect 9680 31690 9732 31696
rect 9692 31482 9720 31690
rect 9680 31476 9732 31482
rect 9680 31418 9732 31424
rect 9588 31272 9640 31278
rect 9588 31214 9640 31220
rect 8944 29844 8996 29850
rect 8944 29786 8996 29792
rect 8956 28150 8984 29786
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9324 29306 9352 29582
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9036 29164 9088 29170
rect 9036 29106 9088 29112
rect 9048 28762 9076 29106
rect 9220 28960 9272 28966
rect 9220 28902 9272 28908
rect 9036 28756 9088 28762
rect 9036 28698 9088 28704
rect 9232 28150 9260 28902
rect 8944 28144 8996 28150
rect 8944 28086 8996 28092
rect 9220 28144 9272 28150
rect 9220 28086 9272 28092
rect 9324 28014 9352 29242
rect 9600 28994 9628 31214
rect 9680 30796 9732 30802
rect 9680 30738 9732 30744
rect 9692 29238 9720 30738
rect 9680 29232 9732 29238
rect 9680 29174 9732 29180
rect 9416 28966 9628 28994
rect 9416 28558 9444 28966
rect 9588 28620 9640 28626
rect 9588 28562 9640 28568
rect 9404 28552 9456 28558
rect 9402 28520 9404 28529
rect 9496 28552 9548 28558
rect 9456 28520 9458 28529
rect 9496 28494 9548 28500
rect 9402 28455 9458 28464
rect 9508 28218 9536 28494
rect 9496 28212 9548 28218
rect 9496 28154 9548 28160
rect 9600 28150 9628 28562
rect 9588 28144 9640 28150
rect 9588 28086 9640 28092
rect 9404 28076 9456 28082
rect 9404 28018 9456 28024
rect 9312 28008 9364 28014
rect 9312 27950 9364 27956
rect 9312 27872 9364 27878
rect 9312 27814 9364 27820
rect 9036 26988 9088 26994
rect 9036 26930 9088 26936
rect 9048 26042 9076 26930
rect 9036 26036 9088 26042
rect 9036 25978 9088 25984
rect 9036 24812 9088 24818
rect 9036 24754 9088 24760
rect 9048 24070 9076 24754
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8484 18352 8536 18358
rect 8484 18294 8536 18300
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 7944 17542 7972 18226
rect 8496 18222 8524 18294
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7840 15700 7892 15706
rect 7840 15642 7892 15648
rect 7760 15286 7880 15314
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7760 14793 7788 15098
rect 7746 14784 7802 14793
rect 7746 14719 7802 14728
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7654 13968 7710 13977
rect 7654 13903 7710 13912
rect 7760 13870 7788 14350
rect 7748 13864 7800 13870
rect 7562 13832 7618 13841
rect 7748 13806 7800 13812
rect 7562 13767 7618 13776
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 12986 7696 13670
rect 7760 13326 7788 13806
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7668 12617 7696 12922
rect 7852 12850 7880 15286
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7654 12608 7710 12617
rect 7654 12543 7710 12552
rect 7852 12306 7880 12786
rect 7944 12434 7972 17478
rect 8680 17202 8708 18770
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9048 17882 9076 18362
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8036 16794 8064 17138
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12646 8340 13126
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 7944 12406 8064 12434
rect 7380 12300 7432 12306
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6564 12102 6592 12294
rect 7380 12242 7432 12248
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6196 7546 6224 9998
rect 6472 9994 6500 11630
rect 7024 11626 7052 12174
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11830 7144 12038
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 7012 11620 7064 11626
rect 7012 11562 7064 11568
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6564 10674 6592 11154
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6368 9920 6420 9926
rect 6368 9862 6420 9868
rect 6380 9382 6408 9862
rect 6472 9518 6500 9930
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6288 8906 6316 9318
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6276 8900 6328 8906
rect 6276 8842 6328 8848
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6564 7886 6592 8774
rect 6656 8498 6684 9114
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 6288 6390 6316 7822
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 6276 6384 6328 6390
rect 6276 6326 6328 6332
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4826 5396 4966
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5368 3534 5396 4150
rect 5460 3942 5488 5510
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5448 3596 5500 3602
rect 5552 3584 5580 6326
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5644 5370 5672 6054
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5500 3556 5580 3584
rect 5448 3538 5500 3544
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 5538 3496 5594 3505
rect 5264 3460 5316 3466
rect 5644 3466 5672 4762
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5828 4146 5856 4626
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5920 4321 5948 4422
rect 5906 4312 5962 4321
rect 5906 4247 5962 4256
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5814 4040 5870 4049
rect 5814 3975 5870 3984
rect 5908 4004 5960 4010
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5538 3431 5594 3440
rect 5632 3460 5684 3466
rect 5264 3402 5316 3408
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4988 2508 5040 2514
rect 4988 2450 5040 2456
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 5460 1902 5488 2858
rect 5448 1896 5500 1902
rect 5448 1838 5500 1844
rect 2964 1420 3016 1426
rect 2964 1362 3016 1368
rect 5552 800 5580 3431
rect 5632 3402 5684 3408
rect 5736 3040 5764 3674
rect 5828 3058 5856 3975
rect 5908 3946 5960 3952
rect 5920 3738 5948 3946
rect 6012 3942 6040 6122
rect 6380 5710 6408 7346
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 6472 6458 6500 6734
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6564 5778 6592 7482
rect 6644 7268 6696 7274
rect 6644 7210 6696 7216
rect 6552 5772 6604 5778
rect 6552 5714 6604 5720
rect 6368 5704 6420 5710
rect 6196 5664 6368 5692
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6104 3738 6132 4218
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 5908 3392 5960 3398
rect 5906 3360 5908 3369
rect 5960 3360 5962 3369
rect 5906 3295 5962 3304
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5644 3012 5764 3040
rect 5816 3052 5868 3058
rect 5644 2774 5672 3012
rect 5816 2994 5868 3000
rect 5814 2816 5870 2825
rect 5644 2746 5764 2774
rect 5814 2751 5870 2760
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 5644 800 5672 2586
rect 5736 800 5764 2746
rect 5828 800 5856 2751
rect 5920 800 5948 3130
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6090 2952 6146 2961
rect 6012 1562 6040 2926
rect 6090 2887 6146 2896
rect 6000 1556 6052 1562
rect 6000 1498 6052 1504
rect 6104 1442 6132 2887
rect 6012 1414 6132 1442
rect 6012 800 6040 1414
rect 6090 1320 6146 1329
rect 6090 1255 6146 1264
rect 6104 800 6132 1255
rect 6196 800 6224 5664
rect 6368 5646 6420 5652
rect 6564 5370 6592 5714
rect 6656 5642 6684 7210
rect 6644 5636 6696 5642
rect 6644 5578 6696 5584
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6380 5234 6408 5306
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6472 5114 6500 5170
rect 6288 5098 6500 5114
rect 6276 5092 6500 5098
rect 6328 5086 6500 5092
rect 6276 5034 6328 5040
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6276 4752 6328 4758
rect 6276 4694 6328 4700
rect 6288 2990 6316 4694
rect 6368 4208 6420 4214
rect 6366 4176 6368 4185
rect 6420 4176 6422 4185
rect 6366 4111 6422 4120
rect 6472 3602 6500 4966
rect 6748 4622 6776 11562
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6840 7342 6868 9862
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 7585 6960 9318
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 7024 8634 7052 8910
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7116 7886 7144 11630
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7300 9654 7328 10610
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7300 8090 7328 9590
rect 7392 9382 7420 12242
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7668 11898 7696 12106
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 6918 7576 6974 7585
rect 6918 7511 6974 7520
rect 7116 7410 7144 7822
rect 7392 7478 7420 9318
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7576 8294 7604 8570
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7576 7478 7604 8230
rect 7944 8090 7972 8366
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7944 7410 7972 8026
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6828 6248 6880 6254
rect 6828 6190 6880 6196
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6552 4480 6604 4486
rect 6552 4422 6604 4428
rect 6564 3618 6592 4422
rect 6736 3936 6788 3942
rect 6734 3904 6736 3913
rect 6788 3904 6790 3913
rect 6734 3839 6790 3848
rect 6460 3596 6512 3602
rect 6564 3590 6684 3618
rect 6840 3602 6868 6190
rect 6932 5914 6960 7346
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7024 5642 7052 6598
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6932 4826 6960 5170
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6460 3538 6512 3544
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 6288 1329 6316 2382
rect 6368 1556 6420 1562
rect 6368 1498 6420 1504
rect 6274 1320 6330 1329
rect 6274 1255 6330 1264
rect 6276 1216 6328 1222
rect 6276 1158 6328 1164
rect 6288 800 6316 1158
rect 6380 800 6408 1498
rect 6472 800 6500 3538
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6564 800 6592 3402
rect 6656 800 6684 3590
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6734 3224 6790 3233
rect 6734 3159 6790 3168
rect 6748 3058 6776 3159
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6748 2446 6776 2994
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6736 2304 6788 2310
rect 6734 2272 6736 2281
rect 6788 2272 6790 2281
rect 6734 2207 6790 2216
rect 6748 1970 6776 2207
rect 6736 1964 6788 1970
rect 6736 1906 6788 1912
rect 6840 800 6868 2926
rect 7024 2774 7052 5578
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7116 4826 7144 5034
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7288 4752 7340 4758
rect 7286 4720 7288 4729
rect 7340 4720 7342 4729
rect 7104 4684 7156 4690
rect 7286 4655 7342 4664
rect 7104 4626 7156 4632
rect 7116 4554 7144 4626
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 2990 7144 4490
rect 7194 4312 7250 4321
rect 7194 4247 7250 4256
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 6932 2746 7052 2774
rect 6932 800 6960 2746
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 7024 800 7052 2518
rect 7208 2106 7236 4247
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 7196 1760 7248 1766
rect 7196 1702 7248 1708
rect 7208 800 7236 1702
rect 7300 800 7328 4082
rect 7392 4026 7420 6258
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 7484 4826 7512 5170
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7576 4622 7604 6054
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7484 4146 7512 4558
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7392 3998 7512 4026
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7392 800 7420 2858
rect 7484 2774 7512 3998
rect 7576 3942 7604 4558
rect 7564 3936 7616 3942
rect 7564 3878 7616 3884
rect 7576 3670 7604 3878
rect 7668 3777 7696 6258
rect 7654 3768 7710 3777
rect 7654 3703 7710 3712
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7668 2990 7696 3703
rect 7760 3534 7788 7142
rect 8036 6254 8064 12406
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8220 9586 8248 10134
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7852 5302 7880 6054
rect 7840 5296 7892 5302
rect 7840 5238 7892 5244
rect 7852 4622 7880 5238
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8036 5137 8064 5170
rect 8022 5128 8078 5137
rect 8022 5063 8078 5072
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7944 4826 7972 4966
rect 7932 4820 7984 4826
rect 7932 4762 7984 4768
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7852 4078 7880 4558
rect 7944 4282 7972 4762
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 8036 4162 8064 5063
rect 7944 4134 8064 4162
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7944 3176 7972 4134
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 7760 3148 7972 3176
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7760 2836 7788 3148
rect 7838 3088 7894 3097
rect 8036 3058 8064 3946
rect 7838 3023 7894 3032
rect 7932 3052 7984 3058
rect 7668 2808 7788 2836
rect 7484 2746 7604 2774
rect 7576 800 7604 2746
rect 7668 800 7696 2808
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 7760 800 7788 2314
rect 7852 800 7880 3023
rect 7932 2994 7984 3000
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7944 800 7972 2994
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8036 800 8064 2790
rect 8128 2446 8156 8774
rect 8312 8090 8340 12582
rect 8404 9926 8432 15302
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8496 8514 8524 16390
rect 8760 13320 8812 13326
rect 8760 13262 8812 13268
rect 8772 11762 8800 13262
rect 9048 13190 9076 17818
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9140 15026 9168 17138
rect 9128 15020 9180 15026
rect 9128 14962 9180 14968
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 9232 12434 9260 22578
rect 9324 15706 9352 27814
rect 9416 26382 9444 28018
rect 9496 27464 9548 27470
rect 9496 27406 9548 27412
rect 9508 27130 9536 27406
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 9600 26382 9628 26862
rect 9692 26586 9720 29174
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9784 26450 9812 32506
rect 9876 29170 9904 34342
rect 10140 32224 10192 32230
rect 10140 32166 10192 32172
rect 10152 31346 10180 32166
rect 10244 31754 10272 34546
rect 10428 33590 10456 34614
rect 10980 34610 11008 34886
rect 10784 34604 10836 34610
rect 10784 34546 10836 34552
rect 10968 34604 11020 34610
rect 10968 34546 11020 34552
rect 10796 34202 10824 34546
rect 10784 34196 10836 34202
rect 10784 34138 10836 34144
rect 10416 33584 10468 33590
rect 10416 33526 10468 33532
rect 10876 32564 10928 32570
rect 10876 32506 10928 32512
rect 10244 31726 10364 31754
rect 10232 31476 10284 31482
rect 10232 31418 10284 31424
rect 10140 31340 10192 31346
rect 10140 31282 10192 31288
rect 10244 31249 10272 31418
rect 10230 31240 10286 31249
rect 10230 31175 10286 31184
rect 9956 30184 10008 30190
rect 9956 30126 10008 30132
rect 9968 29714 9996 30126
rect 9956 29708 10008 29714
rect 9956 29650 10008 29656
rect 9864 29164 9916 29170
rect 9864 29106 9916 29112
rect 9864 27872 9916 27878
rect 9864 27814 9916 27820
rect 9772 26444 9824 26450
rect 9772 26386 9824 26392
rect 9404 26376 9456 26382
rect 9404 26318 9456 26324
rect 9588 26376 9640 26382
rect 9588 26318 9640 26324
rect 9416 25838 9444 26318
rect 9404 25832 9456 25838
rect 9404 25774 9456 25780
rect 9876 25294 9904 27814
rect 10244 27538 10272 31175
rect 10232 27532 10284 27538
rect 10232 27474 10284 27480
rect 10232 27396 10284 27402
rect 10232 27338 10284 27344
rect 10244 27062 10272 27338
rect 10232 27056 10284 27062
rect 10232 26998 10284 27004
rect 9956 25356 10008 25362
rect 9956 25298 10008 25304
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9588 24812 9640 24818
rect 9588 24754 9640 24760
rect 9600 23662 9628 24754
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9692 24206 9720 24550
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9784 23866 9812 25230
rect 9968 24682 9996 25298
rect 9956 24676 10008 24682
rect 9956 24618 10008 24624
rect 10140 24676 10192 24682
rect 10140 24618 10192 24624
rect 9968 24410 9996 24618
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 10152 24138 10180 24618
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9772 23860 9824 23866
rect 9772 23802 9824 23808
rect 9588 23656 9640 23662
rect 9588 23598 9640 23604
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 9876 19938 9904 22918
rect 9968 22030 9996 24006
rect 10140 23724 10192 23730
rect 10140 23666 10192 23672
rect 10152 23526 10180 23666
rect 10140 23520 10192 23526
rect 10140 23462 10192 23468
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 10048 21956 10100 21962
rect 10048 21898 10100 21904
rect 10060 21554 10088 21898
rect 10152 21622 10180 23462
rect 10140 21616 10192 21622
rect 10140 21558 10192 21564
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 9416 17882 9444 19926
rect 9876 19910 10180 19938
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9600 18426 9628 18770
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9680 15904 9732 15910
rect 9680 15846 9732 15852
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9402 15600 9458 15609
rect 9402 15535 9458 15544
rect 9416 15502 9444 15535
rect 9692 15502 9720 15846
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 10152 15026 10180 19910
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9692 14278 9720 14418
rect 9680 14272 9732 14278
rect 9678 14240 9680 14249
rect 9732 14240 9734 14249
rect 9678 14175 9734 14184
rect 9784 13410 9812 14826
rect 10060 14618 10088 14894
rect 10244 14618 10272 26998
rect 10336 26382 10364 31726
rect 10888 31482 10916 32506
rect 10876 31476 10928 31482
rect 10876 31418 10928 31424
rect 10784 31340 10836 31346
rect 10980 31328 11008 34546
rect 11072 33930 11100 35702
rect 11348 35086 11376 35974
rect 11336 35080 11388 35086
rect 11336 35022 11388 35028
rect 11244 34468 11296 34474
rect 11244 34410 11296 34416
rect 11256 34202 11284 34410
rect 11244 34196 11296 34202
rect 11244 34138 11296 34144
rect 11060 33924 11112 33930
rect 11060 33866 11112 33872
rect 11256 33658 11284 34138
rect 11348 33998 11376 35022
rect 11440 34542 11468 36314
rect 11532 35766 11560 38218
rect 11612 37868 11664 37874
rect 11612 37810 11664 37816
rect 11624 37194 11652 37810
rect 11808 37738 11836 38694
rect 11992 37874 12020 39306
rect 12176 37942 12204 40666
rect 12636 40526 12664 41414
rect 12624 40520 12676 40526
rect 12624 40462 12676 40468
rect 12820 40390 12848 42230
rect 13820 42220 13872 42226
rect 13820 42162 13872 42168
rect 14924 42220 14976 42226
rect 14924 42162 14976 42168
rect 13360 42016 13412 42022
rect 13360 41958 13412 41964
rect 13372 41614 13400 41958
rect 13832 41614 13860 42162
rect 14936 41614 14964 42162
rect 13360 41608 13412 41614
rect 13360 41550 13412 41556
rect 13544 41608 13596 41614
rect 13544 41550 13596 41556
rect 13820 41608 13872 41614
rect 13820 41550 13872 41556
rect 14924 41608 14976 41614
rect 14924 41550 14976 41556
rect 13556 41414 13584 41550
rect 13636 41540 13688 41546
rect 13636 41482 13688 41488
rect 13464 41386 13584 41414
rect 13464 41138 13492 41386
rect 13452 41132 13504 41138
rect 13452 41074 13504 41080
rect 12348 40384 12400 40390
rect 12348 40326 12400 40332
rect 12808 40384 12860 40390
rect 12808 40326 12860 40332
rect 12164 37936 12216 37942
rect 12164 37878 12216 37884
rect 11888 37868 11940 37874
rect 11888 37810 11940 37816
rect 11980 37868 12032 37874
rect 11980 37810 12032 37816
rect 11796 37732 11848 37738
rect 11796 37674 11848 37680
rect 11612 37188 11664 37194
rect 11612 37130 11664 37136
rect 11624 35766 11652 37130
rect 11808 37126 11836 37674
rect 11900 37262 11928 37810
rect 11888 37256 11940 37262
rect 11888 37198 11940 37204
rect 11796 37120 11848 37126
rect 11796 37062 11848 37068
rect 11808 36106 11836 37062
rect 12360 36786 12388 40326
rect 12624 40044 12676 40050
rect 12624 39986 12676 39992
rect 12636 39846 12664 39986
rect 12624 39840 12676 39846
rect 12624 39782 12676 39788
rect 12636 38486 12664 39782
rect 12716 39296 12768 39302
rect 12716 39238 12768 39244
rect 12728 38826 12756 39238
rect 12716 38820 12768 38826
rect 12716 38762 12768 38768
rect 12624 38480 12676 38486
rect 12624 38422 12676 38428
rect 12624 38344 12676 38350
rect 12624 38286 12676 38292
rect 12636 37806 12664 38286
rect 12624 37800 12676 37806
rect 12624 37742 12676 37748
rect 12348 36780 12400 36786
rect 12348 36722 12400 36728
rect 12360 36378 12388 36722
rect 12348 36372 12400 36378
rect 12348 36314 12400 36320
rect 11796 36100 11848 36106
rect 11796 36042 11848 36048
rect 11520 35760 11572 35766
rect 11520 35702 11572 35708
rect 11612 35760 11664 35766
rect 11612 35702 11664 35708
rect 11704 35692 11756 35698
rect 11704 35634 11756 35640
rect 11612 34944 11664 34950
rect 11612 34886 11664 34892
rect 11624 34610 11652 34886
rect 11716 34746 11744 35634
rect 11704 34740 11756 34746
rect 11704 34682 11756 34688
rect 11612 34604 11664 34610
rect 11612 34546 11664 34552
rect 11428 34536 11480 34542
rect 11428 34478 11480 34484
rect 11336 33992 11388 33998
rect 11336 33934 11388 33940
rect 11244 33652 11296 33658
rect 11244 33594 11296 33600
rect 11060 32428 11112 32434
rect 11060 32370 11112 32376
rect 11072 31958 11100 32370
rect 11060 31952 11112 31958
rect 11060 31894 11112 31900
rect 10836 31300 11008 31328
rect 10784 31282 10836 31288
rect 10416 31136 10468 31142
rect 10416 31078 10468 31084
rect 10428 29102 10456 31078
rect 10796 30054 10824 31282
rect 11072 30734 11100 31894
rect 11440 31890 11468 34478
rect 11704 34400 11756 34406
rect 11704 34342 11756 34348
rect 11716 34066 11744 34342
rect 11704 34060 11756 34066
rect 11704 34002 11756 34008
rect 11808 32026 11836 36042
rect 11980 35148 12032 35154
rect 11980 35090 12032 35096
rect 11992 34202 12020 35090
rect 12532 34944 12584 34950
rect 12532 34886 12584 34892
rect 11980 34196 12032 34202
rect 11980 34138 12032 34144
rect 12348 33516 12400 33522
rect 12348 33458 12400 33464
rect 12072 32360 12124 32366
rect 12072 32302 12124 32308
rect 12084 32026 12112 32302
rect 11796 32020 11848 32026
rect 11796 31962 11848 31968
rect 12072 32020 12124 32026
rect 12072 31962 12124 31968
rect 11428 31884 11480 31890
rect 11428 31826 11480 31832
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11060 30728 11112 30734
rect 11060 30670 11112 30676
rect 10784 30048 10836 30054
rect 10784 29990 10836 29996
rect 10692 29572 10744 29578
rect 10692 29514 10744 29520
rect 10416 29096 10468 29102
rect 10416 29038 10468 29044
rect 10416 28960 10468 28966
rect 10416 28902 10468 28908
rect 10428 28422 10456 28902
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 10324 26376 10376 26382
rect 10324 26318 10376 26324
rect 10336 25974 10364 26318
rect 10324 25968 10376 25974
rect 10324 25910 10376 25916
rect 10324 25356 10376 25362
rect 10324 25298 10376 25304
rect 10336 24818 10364 25298
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10428 22778 10456 28358
rect 10600 26512 10652 26518
rect 10600 26454 10652 26460
rect 10612 26042 10640 26454
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10704 23905 10732 29514
rect 10796 28558 10824 29990
rect 11716 29850 11744 31282
rect 11808 30938 11836 31962
rect 12084 31754 12112 31962
rect 11900 31726 12112 31754
rect 11900 31346 11928 31726
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 11796 30932 11848 30938
rect 11796 30874 11848 30880
rect 11900 30394 11928 31282
rect 11888 30388 11940 30394
rect 11888 30330 11940 30336
rect 12360 30258 12388 33458
rect 12440 31136 12492 31142
rect 12440 31078 12492 31084
rect 12452 30666 12480 31078
rect 12544 30666 12572 34886
rect 12636 32502 12664 37742
rect 12728 37126 12756 38762
rect 12716 37120 12768 37126
rect 12716 37062 12768 37068
rect 12624 32496 12676 32502
rect 12624 32438 12676 32444
rect 12440 30660 12492 30666
rect 12440 30602 12492 30608
rect 12532 30660 12584 30666
rect 12532 30602 12584 30608
rect 12348 30252 12400 30258
rect 12348 30194 12400 30200
rect 11704 29844 11756 29850
rect 11704 29786 11756 29792
rect 11980 29844 12032 29850
rect 11980 29786 12032 29792
rect 10968 29572 11020 29578
rect 10968 29514 11020 29520
rect 10980 29306 11008 29514
rect 10968 29300 11020 29306
rect 10968 29242 11020 29248
rect 11704 28688 11756 28694
rect 11704 28630 11756 28636
rect 10784 28552 10836 28558
rect 10784 28494 10836 28500
rect 11520 28416 11572 28422
rect 11520 28358 11572 28364
rect 11152 28008 11204 28014
rect 11152 27950 11204 27956
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10888 26314 10916 26930
rect 11164 26926 11192 27950
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 10876 26308 10928 26314
rect 10876 26250 10928 26256
rect 10690 23896 10746 23905
rect 10690 23831 10746 23840
rect 10416 22772 10468 22778
rect 10416 22714 10468 22720
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10336 22438 10364 22578
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10336 22166 10364 22374
rect 10324 22160 10376 22166
rect 10324 22102 10376 22108
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10520 19378 10548 19654
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10336 16114 10364 16390
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10520 15502 10548 19314
rect 10612 15502 10640 21830
rect 10704 21146 10732 23831
rect 10888 21434 10916 26250
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 11072 24274 11100 25298
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 11072 23798 11100 24210
rect 11060 23792 11112 23798
rect 11060 23734 11112 23740
rect 11072 23118 11100 23734
rect 11060 23112 11112 23118
rect 11060 23054 11112 23060
rect 11060 22568 11112 22574
rect 11060 22510 11112 22516
rect 11072 22030 11100 22510
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 11072 21554 11100 21966
rect 11060 21548 11112 21554
rect 11060 21490 11112 21496
rect 10796 21406 10916 21434
rect 10692 21140 10744 21146
rect 10692 21082 10744 21088
rect 10796 15978 10824 21406
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10980 18154 11008 20810
rect 11060 18420 11112 18426
rect 11060 18362 11112 18368
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10980 18057 11008 18090
rect 10966 18048 11022 18057
rect 10966 17983 11022 17992
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10888 16250 10916 17818
rect 10876 16244 10928 16250
rect 10876 16186 10928 16192
rect 10784 15972 10836 15978
rect 10784 15914 10836 15920
rect 11072 15570 11100 18362
rect 11164 17882 11192 26862
rect 11336 25764 11388 25770
rect 11336 25706 11388 25712
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11256 24070 11284 24142
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 11256 20602 11284 24006
rect 11348 23322 11376 25706
rect 11336 23316 11388 23322
rect 11336 23258 11388 23264
rect 11532 22094 11560 28358
rect 11716 28082 11744 28630
rect 11992 28150 12020 29786
rect 12164 29640 12216 29646
rect 12164 29582 12216 29588
rect 11980 28144 12032 28150
rect 11980 28086 12032 28092
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 11716 27674 11744 28018
rect 11704 27668 11756 27674
rect 11704 27610 11756 27616
rect 12176 27538 12204 29582
rect 12360 28014 12388 30194
rect 12452 29073 12480 30602
rect 12438 29064 12494 29073
rect 12438 28999 12494 29008
rect 12544 28558 12572 30602
rect 12624 29572 12676 29578
rect 12624 29514 12676 29520
rect 12532 28552 12584 28558
rect 12532 28494 12584 28500
rect 12348 28008 12400 28014
rect 12348 27950 12400 27956
rect 12164 27532 12216 27538
rect 12164 27474 12216 27480
rect 12176 26858 12204 27474
rect 12164 26852 12216 26858
rect 12164 26794 12216 26800
rect 12176 25362 12204 26794
rect 12360 26586 12388 27950
rect 12544 26994 12572 28494
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 12164 25356 12216 25362
rect 12164 25298 12216 25304
rect 12440 24744 12492 24750
rect 12440 24686 12492 24692
rect 12256 24608 12308 24614
rect 12256 24550 12308 24556
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 11900 24206 11928 24346
rect 12268 24206 12296 24550
rect 12452 24206 12480 24686
rect 12636 24682 12664 29514
rect 12624 24676 12676 24682
rect 12624 24618 12676 24624
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 12072 24200 12124 24206
rect 12072 24142 12124 24148
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12440 24200 12492 24206
rect 12440 24142 12492 24148
rect 11612 24064 11664 24070
rect 11612 24006 11664 24012
rect 11624 23118 11652 24006
rect 12084 23866 12112 24142
rect 12072 23860 12124 23866
rect 12072 23802 12124 23808
rect 11980 23724 12032 23730
rect 11980 23666 12032 23672
rect 11888 23520 11940 23526
rect 11888 23462 11940 23468
rect 11612 23112 11664 23118
rect 11612 23054 11664 23060
rect 11704 23044 11756 23050
rect 11704 22986 11756 22992
rect 11716 22642 11744 22986
rect 11900 22642 11928 23462
rect 11992 23322 12020 23666
rect 11980 23316 12032 23322
rect 11980 23258 12032 23264
rect 11992 22710 12020 23258
rect 11980 22704 12032 22710
rect 11980 22646 12032 22652
rect 11704 22636 11756 22642
rect 11704 22578 11756 22584
rect 11888 22636 11940 22642
rect 11888 22578 11940 22584
rect 11532 22066 11652 22094
rect 11428 21344 11480 21350
rect 11428 21286 11480 21292
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11336 19848 11388 19854
rect 11256 19796 11336 19802
rect 11256 19790 11388 19796
rect 11256 19774 11376 19790
rect 11256 19174 11284 19774
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11348 19514 11376 19654
rect 11336 19508 11388 19514
rect 11336 19450 11388 19456
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11256 18766 11284 19110
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11256 18154 11284 18702
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11164 16046 11192 16390
rect 11440 16114 11468 21286
rect 11624 21078 11652 22066
rect 11716 21894 11744 22578
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 12452 21418 12480 24142
rect 12636 23118 12664 24618
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12728 22094 12756 37062
rect 12820 35086 12848 40326
rect 13464 39506 13492 41074
rect 13648 41070 13676 41482
rect 13832 41478 13860 41550
rect 15200 41540 15252 41546
rect 15200 41482 15252 41488
rect 13820 41472 13872 41478
rect 13820 41414 13872 41420
rect 13636 41064 13688 41070
rect 13636 41006 13688 41012
rect 13452 39500 13504 39506
rect 13452 39442 13504 39448
rect 13648 39370 13676 41006
rect 13728 40520 13780 40526
rect 13728 40462 13780 40468
rect 13740 40186 13768 40462
rect 13832 40458 13860 41414
rect 13912 40996 13964 41002
rect 13912 40938 13964 40944
rect 13820 40452 13872 40458
rect 13820 40394 13872 40400
rect 13728 40180 13780 40186
rect 13728 40122 13780 40128
rect 13636 39364 13688 39370
rect 13636 39306 13688 39312
rect 13648 38962 13676 39306
rect 13636 38956 13688 38962
rect 13636 38898 13688 38904
rect 13360 38344 13412 38350
rect 13360 38286 13412 38292
rect 13176 38276 13228 38282
rect 13176 38218 13228 38224
rect 13188 38010 13216 38218
rect 13176 38004 13228 38010
rect 13176 37946 13228 37952
rect 13268 37868 13320 37874
rect 13372 37856 13400 38286
rect 13320 37828 13400 37856
rect 13268 37810 13320 37816
rect 13280 37262 13308 37810
rect 13636 37664 13688 37670
rect 13636 37606 13688 37612
rect 13360 37324 13412 37330
rect 13360 37266 13412 37272
rect 13268 37256 13320 37262
rect 13268 37198 13320 37204
rect 13280 36718 13308 37198
rect 13268 36712 13320 36718
rect 13268 36654 13320 36660
rect 12992 36644 13044 36650
rect 12992 36586 13044 36592
rect 13004 35086 13032 36586
rect 13372 35766 13400 37266
rect 13648 37194 13676 37606
rect 13636 37188 13688 37194
rect 13636 37130 13688 37136
rect 13360 35760 13412 35766
rect 13360 35702 13412 35708
rect 13636 35760 13688 35766
rect 13636 35702 13688 35708
rect 13544 35624 13596 35630
rect 13544 35566 13596 35572
rect 12808 35080 12860 35086
rect 12808 35022 12860 35028
rect 12992 35080 13044 35086
rect 12992 35022 13044 35028
rect 13004 34542 13032 35022
rect 13556 35018 13584 35566
rect 13544 35012 13596 35018
rect 13544 34954 13596 34960
rect 13556 34678 13584 34954
rect 13544 34672 13596 34678
rect 13544 34614 13596 34620
rect 12992 34536 13044 34542
rect 12992 34478 13044 34484
rect 12900 32428 12952 32434
rect 12900 32370 12952 32376
rect 12808 31816 12860 31822
rect 12808 31758 12860 31764
rect 12820 31482 12848 31758
rect 12912 31686 12940 32370
rect 12900 31680 12952 31686
rect 12900 31622 12952 31628
rect 12808 31476 12860 31482
rect 12808 31418 12860 31424
rect 12912 30734 12940 31622
rect 13004 30734 13032 34478
rect 13084 32496 13136 32502
rect 13084 32438 13136 32444
rect 13452 32496 13504 32502
rect 13452 32438 13504 32444
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 13004 28994 13032 30670
rect 12820 28966 13032 28994
rect 12820 28558 12848 28966
rect 12808 28552 12860 28558
rect 12808 28494 12860 28500
rect 12820 26994 12848 28494
rect 13096 28422 13124 32438
rect 13360 32224 13412 32230
rect 13360 32166 13412 32172
rect 13268 31476 13320 31482
rect 13268 31418 13320 31424
rect 13176 31204 13228 31210
rect 13176 31146 13228 31152
rect 13188 29646 13216 31146
rect 13176 29640 13228 29646
rect 13176 29582 13228 29588
rect 13280 29238 13308 31418
rect 13372 31346 13400 32166
rect 13360 31340 13412 31346
rect 13360 31282 13412 31288
rect 13464 30802 13492 32438
rect 13648 31754 13676 35702
rect 13740 34746 13768 40122
rect 13924 37738 13952 40938
rect 15016 40928 15068 40934
rect 15016 40870 15068 40876
rect 14280 40452 14332 40458
rect 14280 40394 14332 40400
rect 14292 38554 14320 40394
rect 14924 40384 14976 40390
rect 14924 40326 14976 40332
rect 14556 40044 14608 40050
rect 14556 39986 14608 39992
rect 14568 39642 14596 39986
rect 14556 39636 14608 39642
rect 14556 39578 14608 39584
rect 14936 39438 14964 40326
rect 15028 40186 15056 40870
rect 15212 40390 15240 41482
rect 15200 40384 15252 40390
rect 15200 40326 15252 40332
rect 15016 40180 15068 40186
rect 15016 40122 15068 40128
rect 14556 39432 14608 39438
rect 14556 39374 14608 39380
rect 14924 39432 14976 39438
rect 14924 39374 14976 39380
rect 14568 39302 14596 39374
rect 14556 39296 14608 39302
rect 14556 39238 14608 39244
rect 14280 38548 14332 38554
rect 14280 38490 14332 38496
rect 13912 37732 13964 37738
rect 13912 37674 13964 37680
rect 14740 36780 14792 36786
rect 14740 36722 14792 36728
rect 14752 36378 14780 36722
rect 14740 36372 14792 36378
rect 14740 36314 14792 36320
rect 15028 36174 15056 40122
rect 14096 36168 14148 36174
rect 14096 36110 14148 36116
rect 14372 36168 14424 36174
rect 14372 36110 14424 36116
rect 15016 36168 15068 36174
rect 15016 36110 15068 36116
rect 14108 35834 14136 36110
rect 14096 35828 14148 35834
rect 14096 35770 14148 35776
rect 13728 34740 13780 34746
rect 13728 34682 13780 34688
rect 14384 34202 14412 36110
rect 15028 35766 15056 36110
rect 15016 35760 15068 35766
rect 15016 35702 15068 35708
rect 14924 34944 14976 34950
rect 14924 34886 14976 34892
rect 14372 34196 14424 34202
rect 14372 34138 14424 34144
rect 14372 33924 14424 33930
rect 14372 33866 14424 33872
rect 13820 33108 13872 33114
rect 13820 33050 13872 33056
rect 13832 32434 13860 33050
rect 14096 32904 14148 32910
rect 14096 32846 14148 32852
rect 13820 32428 13872 32434
rect 13820 32370 13872 32376
rect 13648 31726 13768 31754
rect 13740 31346 13768 31726
rect 13728 31340 13780 31346
rect 13728 31282 13780 31288
rect 13740 31142 13768 31282
rect 13728 31136 13780 31142
rect 13728 31078 13780 31084
rect 13452 30796 13504 30802
rect 13452 30738 13504 30744
rect 13268 29232 13320 29238
rect 13268 29174 13320 29180
rect 13740 29170 13768 31078
rect 14108 30802 14136 32846
rect 14188 32564 14240 32570
rect 14188 32506 14240 32512
rect 14200 32434 14228 32506
rect 14384 32502 14412 33866
rect 14556 33448 14608 33454
rect 14556 33390 14608 33396
rect 14464 32836 14516 32842
rect 14464 32778 14516 32784
rect 14476 32570 14504 32778
rect 14464 32564 14516 32570
rect 14464 32506 14516 32512
rect 14372 32496 14424 32502
rect 14372 32438 14424 32444
rect 14568 32434 14596 33390
rect 14936 32910 14964 34886
rect 14924 32904 14976 32910
rect 14924 32846 14976 32852
rect 15200 32768 15252 32774
rect 15200 32710 15252 32716
rect 15212 32502 15240 32710
rect 15200 32496 15252 32502
rect 15200 32438 15252 32444
rect 14188 32428 14240 32434
rect 14188 32370 14240 32376
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 14924 32428 14976 32434
rect 14924 32370 14976 32376
rect 14200 31958 14228 32370
rect 14936 32026 14964 32370
rect 14924 32020 14976 32026
rect 14924 31962 14976 31968
rect 14188 31952 14240 31958
rect 14188 31894 14240 31900
rect 14096 30796 14148 30802
rect 14096 30738 14148 30744
rect 14004 30592 14056 30598
rect 14004 30534 14056 30540
rect 14016 30258 14044 30534
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 14004 30116 14056 30122
rect 14004 30058 14056 30064
rect 13452 29164 13504 29170
rect 13452 29106 13504 29112
rect 13728 29164 13780 29170
rect 13728 29106 13780 29112
rect 13464 29034 13492 29106
rect 13176 29028 13228 29034
rect 13176 28970 13228 28976
rect 13452 29028 13504 29034
rect 13452 28970 13504 28976
rect 12992 28416 13044 28422
rect 12992 28358 13044 28364
rect 13084 28416 13136 28422
rect 13084 28358 13136 28364
rect 13004 28082 13032 28358
rect 13096 28218 13124 28358
rect 13084 28212 13136 28218
rect 13084 28154 13136 28160
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 13188 27470 13216 28970
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 12900 27396 12952 27402
rect 12900 27338 12952 27344
rect 12808 26988 12860 26994
rect 12808 26930 12860 26936
rect 12912 26926 12940 27338
rect 12900 26920 12952 26926
rect 12900 26862 12952 26868
rect 13464 26042 13492 28970
rect 13740 28762 13768 29106
rect 13728 28756 13780 28762
rect 13728 28698 13780 28704
rect 13544 28484 13596 28490
rect 13544 28426 13596 28432
rect 13556 27674 13584 28426
rect 14016 28082 14044 30058
rect 14200 29782 14228 31894
rect 15304 31754 15332 47534
rect 16672 42220 16724 42226
rect 16672 42162 16724 42168
rect 15568 42016 15620 42022
rect 15568 41958 15620 41964
rect 15384 41608 15436 41614
rect 15384 41550 15436 41556
rect 15396 41138 15424 41550
rect 15580 41274 15608 41958
rect 15752 41608 15804 41614
rect 15752 41550 15804 41556
rect 15568 41268 15620 41274
rect 15568 41210 15620 41216
rect 15384 41132 15436 41138
rect 15384 41074 15436 41080
rect 15764 41002 15792 41550
rect 15752 40996 15804 41002
rect 15752 40938 15804 40944
rect 16580 40520 16632 40526
rect 16500 40480 16580 40508
rect 16028 40384 16080 40390
rect 16028 40326 16080 40332
rect 15660 39976 15712 39982
rect 15660 39918 15712 39924
rect 15672 37262 15700 39918
rect 16040 37874 16068 40326
rect 16500 39982 16528 40480
rect 16580 40462 16632 40468
rect 16488 39976 16540 39982
rect 16488 39918 16540 39924
rect 16500 39438 16528 39918
rect 16488 39432 16540 39438
rect 16488 39374 16540 39380
rect 16684 39302 16712 42162
rect 16764 41540 16816 41546
rect 16764 41482 16816 41488
rect 16776 40458 16804 41482
rect 17328 41414 17356 55762
rect 17420 55214 17448 56306
rect 18052 55616 18104 55622
rect 18050 55584 18052 55593
rect 18104 55584 18106 55593
rect 18050 55519 18106 55528
rect 18708 55418 18736 56306
rect 18788 56160 18840 56166
rect 18788 56102 18840 56108
rect 18696 55412 18748 55418
rect 18696 55354 18748 55360
rect 17420 55186 17540 55214
rect 17512 41414 17540 55186
rect 18420 41540 18472 41546
rect 18420 41482 18472 41488
rect 17684 41472 17736 41478
rect 17684 41414 17736 41420
rect 17236 41386 17356 41414
rect 17420 41386 17540 41414
rect 16764 40452 16816 40458
rect 16764 40394 16816 40400
rect 16672 39296 16724 39302
rect 16672 39238 16724 39244
rect 16684 38282 16712 39238
rect 16672 38276 16724 38282
rect 16672 38218 16724 38224
rect 17132 38208 17184 38214
rect 17132 38150 17184 38156
rect 17144 37874 17172 38150
rect 16028 37868 16080 37874
rect 16028 37810 16080 37816
rect 17132 37868 17184 37874
rect 17132 37810 17184 37816
rect 17040 37800 17092 37806
rect 17040 37742 17092 37748
rect 16948 37664 17000 37670
rect 16948 37606 17000 37612
rect 15660 37256 15712 37262
rect 15660 37198 15712 37204
rect 16672 37188 16724 37194
rect 16672 37130 16724 37136
rect 15476 37120 15528 37126
rect 15476 37062 15528 37068
rect 15488 36922 15516 37062
rect 16684 36922 16712 37130
rect 15476 36916 15528 36922
rect 15476 36858 15528 36864
rect 16672 36916 16724 36922
rect 16672 36858 16724 36864
rect 15488 36174 15516 36858
rect 16960 36786 16988 37606
rect 17052 37126 17080 37742
rect 17040 37120 17092 37126
rect 17040 37062 17092 37068
rect 16948 36780 17000 36786
rect 16948 36722 17000 36728
rect 16856 36712 16908 36718
rect 16856 36654 16908 36660
rect 16868 36242 16896 36654
rect 16856 36236 16908 36242
rect 16856 36178 16908 36184
rect 15476 36168 15528 36174
rect 15476 36110 15528 36116
rect 15660 36100 15712 36106
rect 15660 36042 15712 36048
rect 15476 34672 15528 34678
rect 15476 34614 15528 34620
rect 15488 33590 15516 34614
rect 15568 33856 15620 33862
rect 15568 33798 15620 33804
rect 15580 33590 15608 33798
rect 15476 33584 15528 33590
rect 15476 33526 15528 33532
rect 15568 33584 15620 33590
rect 15568 33526 15620 33532
rect 15672 33454 15700 36042
rect 16960 36038 16988 36722
rect 17052 36174 17080 37062
rect 17132 36780 17184 36786
rect 17132 36722 17184 36728
rect 17144 36378 17172 36722
rect 17132 36372 17184 36378
rect 17132 36314 17184 36320
rect 17040 36168 17092 36174
rect 17040 36110 17092 36116
rect 16948 36032 17000 36038
rect 16948 35974 17000 35980
rect 17040 35556 17092 35562
rect 17040 35498 17092 35504
rect 16948 35148 17000 35154
rect 16948 35090 17000 35096
rect 16960 34746 16988 35090
rect 16948 34740 17000 34746
rect 16948 34682 17000 34688
rect 16960 34610 16988 34682
rect 16948 34604 17000 34610
rect 16948 34546 17000 34552
rect 16396 33992 16448 33998
rect 16396 33934 16448 33940
rect 16304 33584 16356 33590
rect 16304 33526 16356 33532
rect 15660 33448 15712 33454
rect 15660 33390 15712 33396
rect 15844 33040 15896 33046
rect 15844 32982 15896 32988
rect 15384 32496 15436 32502
rect 15384 32438 15436 32444
rect 15212 31726 15332 31754
rect 14280 31340 14332 31346
rect 14280 31282 14332 31288
rect 14292 30870 14320 31282
rect 15016 31272 15068 31278
rect 15014 31240 15016 31249
rect 15068 31240 15070 31249
rect 15014 31175 15070 31184
rect 14924 31136 14976 31142
rect 14924 31078 14976 31084
rect 14280 30864 14332 30870
rect 14280 30806 14332 30812
rect 14832 30796 14884 30802
rect 14832 30738 14884 30744
rect 14844 30394 14872 30738
rect 14936 30734 14964 31078
rect 14924 30728 14976 30734
rect 14924 30670 14976 30676
rect 14924 30592 14976 30598
rect 14924 30534 14976 30540
rect 14832 30388 14884 30394
rect 14832 30330 14884 30336
rect 14188 29776 14240 29782
rect 14188 29718 14240 29724
rect 14188 29504 14240 29510
rect 14188 29446 14240 29452
rect 14200 29034 14228 29446
rect 14464 29096 14516 29102
rect 14464 29038 14516 29044
rect 14188 29028 14240 29034
rect 14188 28970 14240 28976
rect 14476 28762 14504 29038
rect 14464 28756 14516 28762
rect 14464 28698 14516 28704
rect 14844 28150 14872 30330
rect 14936 29646 14964 30534
rect 14924 29640 14976 29646
rect 14924 29582 14976 29588
rect 14936 29238 14964 29582
rect 14924 29232 14976 29238
rect 14924 29174 14976 29180
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 14924 28552 14976 28558
rect 14924 28494 14976 28500
rect 14832 28144 14884 28150
rect 14832 28086 14884 28092
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 13544 27668 13596 27674
rect 13544 27610 13596 27616
rect 14016 27606 14044 28018
rect 14936 27946 14964 28494
rect 15120 28218 15148 29106
rect 15108 28212 15160 28218
rect 15108 28154 15160 28160
rect 14924 27940 14976 27946
rect 14924 27882 14976 27888
rect 15016 27872 15068 27878
rect 15016 27814 15068 27820
rect 14004 27600 14056 27606
rect 14004 27542 14056 27548
rect 13636 26920 13688 26926
rect 13636 26862 13688 26868
rect 13452 26036 13504 26042
rect 13452 25978 13504 25984
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 12820 25702 12848 25842
rect 12808 25696 12860 25702
rect 12808 25638 12860 25644
rect 12820 22166 12848 25638
rect 13360 25288 13412 25294
rect 13360 25230 13412 25236
rect 13176 24608 13228 24614
rect 13176 24550 13228 24556
rect 13188 24206 13216 24550
rect 13372 24206 13400 25230
rect 13544 24336 13596 24342
rect 13544 24278 13596 24284
rect 13176 24200 13228 24206
rect 13176 24142 13228 24148
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12912 23730 12940 24006
rect 13556 23730 13584 24278
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 13544 23724 13596 23730
rect 13544 23666 13596 23672
rect 12900 22432 12952 22438
rect 12900 22374 12952 22380
rect 12808 22160 12860 22166
rect 12808 22102 12860 22108
rect 12636 22066 12756 22094
rect 12440 21412 12492 21418
rect 12440 21354 12492 21360
rect 11612 21072 11664 21078
rect 11612 21014 11664 21020
rect 11624 20602 11652 21014
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11900 19854 11928 20538
rect 12440 19916 12492 19922
rect 12440 19858 12492 19864
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 11716 19514 11744 19790
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11704 19236 11756 19242
rect 11704 19178 11756 19184
rect 11520 18692 11572 18698
rect 11520 18634 11572 18640
rect 11532 18426 11560 18634
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11532 17542 11560 18226
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11532 16998 11560 17478
rect 11520 16992 11572 16998
rect 11520 16934 11572 16940
rect 11624 16114 11652 18566
rect 11716 18426 11744 19178
rect 12176 18970 12204 19790
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11992 18290 12020 18566
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 12084 17610 12112 18294
rect 12176 18290 12204 18906
rect 12452 18358 12480 19858
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12544 18766 12572 19314
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12452 18170 12480 18294
rect 12544 18272 12572 18702
rect 12636 18340 12664 22066
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12728 20058 12756 20402
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12728 19174 12756 19790
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12728 18902 12756 19110
rect 12716 18896 12768 18902
rect 12716 18838 12768 18844
rect 12636 18312 12756 18340
rect 12544 18244 12664 18272
rect 12452 18154 12572 18170
rect 12452 18148 12584 18154
rect 12452 18142 12532 18148
rect 12532 18090 12584 18096
rect 12636 17678 12664 18244
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11702 16688 11758 16697
rect 11702 16623 11758 16632
rect 11428 16108 11480 16114
rect 11428 16050 11480 16056
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11716 16046 11744 16623
rect 11796 16108 11848 16114
rect 11796 16050 11848 16056
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 10876 15564 10928 15570
rect 10876 15506 10928 15512
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 14006 10824 14214
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 9692 13382 9812 13410
rect 9692 12782 9720 13382
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9232 12406 9628 12434
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9232 10470 9260 10678
rect 9220 10464 9272 10470
rect 9272 10424 9352 10452
rect 9220 10406 9272 10412
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8956 9722 8984 9998
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 9140 9654 9168 9862
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8404 8486 8524 8514
rect 8864 8498 8892 9454
rect 8852 8492 8904 8498
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8220 4486 8248 6598
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8220 4146 8248 4422
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8312 3942 8340 5578
rect 8404 4826 8432 8486
rect 8852 8434 8904 8440
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8588 6798 8616 7142
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 6322 8524 6598
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8482 5128 8538 5137
rect 8482 5063 8484 5072
rect 8536 5063 8538 5072
rect 8484 5034 8536 5040
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8588 4706 8616 6734
rect 8680 6186 8708 6802
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8668 6180 8720 6186
rect 8668 6122 8720 6128
rect 8404 4678 8616 4706
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8298 3768 8354 3777
rect 8298 3703 8300 3712
rect 8352 3703 8354 3712
rect 8300 3674 8352 3680
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8128 1766 8156 2382
rect 8116 1760 8168 1766
rect 8116 1702 8168 1708
rect 8116 1624 8168 1630
rect 8116 1566 8168 1572
rect 8128 800 8156 1566
rect 8220 800 8248 3470
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 8312 800 8340 3402
rect 8404 800 8432 4678
rect 8482 3632 8538 3641
rect 8680 3602 8708 6122
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8760 5160 8812 5166
rect 8760 5102 8812 5108
rect 8772 4282 8800 5102
rect 8864 5030 8892 6054
rect 8852 5024 8904 5030
rect 8852 4966 8904 4972
rect 8864 4622 8892 4966
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8956 4282 8984 4762
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8772 3670 8800 4014
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 8482 3567 8538 3576
rect 8668 3596 8720 3602
rect 8496 2378 8524 3567
rect 8668 3538 8720 3544
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8496 800 8524 2314
rect 8588 800 8616 3334
rect 8864 3126 8892 4082
rect 8942 4040 8998 4049
rect 8942 3975 8998 3984
rect 8956 3194 8984 3975
rect 9048 3670 9076 6258
rect 9140 3738 9168 6598
rect 9232 4146 9260 7686
rect 9324 4826 9352 10424
rect 9600 9654 9628 12406
rect 9692 12186 9720 12718
rect 9784 12442 9812 13194
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 9772 12436 9824 12442
rect 10520 12434 10548 13126
rect 10520 12406 10732 12434
rect 9772 12378 9824 12384
rect 10704 12238 10732 12406
rect 10692 12232 10744 12238
rect 9692 12170 9812 12186
rect 10692 12174 10744 12180
rect 9692 12164 9824 12170
rect 9692 12158 9772 12164
rect 9772 12106 9824 12112
rect 9784 11150 9812 12106
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10606 9720 10950
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9508 8498 9536 8910
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9416 8022 9444 8434
rect 9600 8294 9628 9590
rect 9784 9042 9812 11086
rect 10140 11076 10192 11082
rect 10140 11018 10192 11024
rect 10152 10674 10180 11018
rect 9956 10668 10008 10674
rect 9956 10610 10008 10616
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 9864 9104 9916 9110
rect 9864 9046 9916 9052
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9784 8838 9812 8978
rect 9876 8974 9904 9046
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9692 8566 9720 8774
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9416 6322 9444 7958
rect 9508 7750 9536 8026
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 6730 9536 7686
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9220 4140 9272 4146
rect 9272 4100 9352 4128
rect 9220 4082 9272 4088
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9036 3664 9088 3670
rect 9036 3606 9088 3612
rect 9140 3346 9168 3674
rect 9232 3398 9260 3946
rect 9048 3318 9168 3346
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8760 3120 8812 3126
rect 8760 3062 8812 3068
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 8772 800 8800 3062
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8956 2774 8984 2926
rect 9048 2922 9076 3318
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 8956 2746 9076 2774
rect 8852 1420 8904 1426
rect 8852 1362 8904 1368
rect 8864 800 8892 1362
rect 9048 800 9076 2746
rect 9140 800 9168 3130
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9232 2514 9260 3062
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9324 800 9352 4100
rect 9416 3534 9444 4626
rect 9600 3738 9628 8230
rect 9784 7993 9812 8230
rect 9770 7984 9826 7993
rect 9770 7919 9826 7928
rect 9784 4282 9812 7919
rect 9876 6934 9904 8910
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9968 6798 9996 10610
rect 10428 10130 10456 10610
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10324 9920 10376 9926
rect 10322 9888 10324 9897
rect 10376 9888 10378 9897
rect 10322 9823 10378 9832
rect 10428 9722 10456 10066
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10244 8906 10272 9114
rect 10336 9110 10364 9318
rect 10324 9104 10376 9110
rect 10324 9046 10376 9052
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10048 7268 10100 7274
rect 10048 7210 10100 7216
rect 10060 6866 10088 7210
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10138 6896 10194 6905
rect 10048 6860 10100 6866
rect 10138 6831 10194 6840
rect 10048 6802 10100 6808
rect 10152 6798 10180 6831
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9876 6390 9904 6598
rect 9864 6384 9916 6390
rect 9864 6326 9916 6332
rect 10232 5772 10284 5778
rect 10232 5714 10284 5720
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9772 4276 9824 4282
rect 9772 4218 9824 4224
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9508 2854 9536 3674
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 9416 800 9444 2518
rect 9508 2038 9536 2790
rect 9496 2032 9548 2038
rect 9496 1974 9548 1980
rect 9600 800 9628 3470
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9784 1442 9812 2790
rect 9692 1414 9812 1442
rect 9692 800 9720 1414
rect 9968 800 9996 5646
rect 10046 4040 10102 4049
rect 10046 3975 10102 3984
rect 10060 3058 10088 3975
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10244 800 10272 5714
rect 10336 3534 10364 7142
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10428 3058 10456 9318
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10414 2680 10470 2689
rect 10414 2615 10416 2624
rect 10468 2615 10470 2624
rect 10416 2586 10468 2592
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 10336 2106 10364 2314
rect 10324 2100 10376 2106
rect 10324 2042 10376 2048
rect 10428 2038 10456 2586
rect 10416 2032 10468 2038
rect 10416 1974 10468 1980
rect 10520 800 10548 6734
rect 10612 4146 10640 12038
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10704 3534 10732 12174
rect 10796 10962 10824 13942
rect 10888 11626 10916 15506
rect 11716 15314 11744 15982
rect 11808 15434 11836 16050
rect 11900 15502 11928 17478
rect 12176 16794 12204 17614
rect 12360 17338 12388 17614
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12636 17270 12664 17614
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12440 17196 12492 17202
rect 12440 17138 12492 17144
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 11980 16108 12032 16114
rect 11980 16050 12032 16056
rect 11992 15706 12020 16050
rect 12452 15706 12480 17138
rect 12624 16652 12676 16658
rect 12624 16594 12676 16600
rect 12636 16114 12664 16594
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11796 15428 11848 15434
rect 11796 15370 11848 15376
rect 11716 15286 11836 15314
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11072 12918 11100 14962
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11532 12238 11560 12582
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11716 12102 11744 12786
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 10796 10934 10916 10962
rect 10888 10606 10916 10934
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10888 7750 10916 10542
rect 11348 9058 11376 11018
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11256 9042 11376 9058
rect 11244 9036 11376 9042
rect 11296 9030 11376 9036
rect 11244 8978 11296 8984
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11256 8634 11284 8842
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7206 10916 7686
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10784 5840 10836 5846
rect 10784 5782 10836 5788
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 10600 2644 10652 2650
rect 10600 2586 10652 2592
rect 10612 1426 10640 2586
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 10704 1902 10732 2042
rect 10692 1896 10744 1902
rect 10692 1838 10744 1844
rect 10600 1420 10652 1426
rect 10600 1362 10652 1368
rect 10796 800 10824 5782
rect 10888 4826 10916 7142
rect 11060 6724 11112 6730
rect 11060 6666 11112 6672
rect 11072 6186 11100 6666
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11348 5846 11376 9030
rect 11532 8566 11560 10542
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11532 5710 11560 6394
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11336 5704 11388 5710
rect 11336 5646 11388 5652
rect 11520 5704 11572 5710
rect 11520 5646 11572 5652
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10874 3224 10930 3233
rect 10874 3159 10930 3168
rect 10888 3058 10916 3159
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10980 2774 11008 5170
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11256 4622 11284 5102
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11256 3942 11284 4558
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11256 3126 11284 3878
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 10980 2746 11100 2774
rect 11072 800 11100 2746
rect 11348 800 11376 5646
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11440 4010 11468 4762
rect 11532 4758 11560 5170
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11532 4554 11560 4694
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11532 4146 11560 4490
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11624 800 11652 6054
rect 11716 2446 11744 8298
rect 11808 4826 11836 15286
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11992 14414 12020 14962
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11992 13002 12020 14350
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12084 13938 12112 14214
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 11992 12974 12112 13002
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 9042 11928 10950
rect 11992 10810 12020 12718
rect 12084 12170 12112 12974
rect 12544 12442 12572 13330
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12072 12164 12124 12170
rect 12072 12106 12124 12112
rect 12348 12164 12400 12170
rect 12348 12106 12400 12112
rect 12084 11762 12112 12106
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12360 11694 12388 12106
rect 12544 11830 12572 12174
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 11992 9994 12020 10542
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 7478 11928 8774
rect 11992 8430 12020 9930
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 11888 7472 11940 7478
rect 11888 7414 11940 7420
rect 12084 7410 12112 7958
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 12360 6798 12388 11630
rect 12544 11218 12572 11766
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12636 10742 12664 16050
rect 12728 11082 12756 18312
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12820 16114 12848 16390
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12820 15910 12848 16050
rect 12808 15904 12860 15910
rect 12808 15846 12860 15852
rect 12820 15162 12848 15846
rect 12912 15502 12940 22374
rect 13648 22094 13676 26862
rect 14096 26308 14148 26314
rect 14096 26250 14148 26256
rect 14108 25906 14136 26250
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 13820 25832 13872 25838
rect 13820 25774 13872 25780
rect 13912 25832 13964 25838
rect 13912 25774 13964 25780
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 13740 24342 13768 24754
rect 13728 24336 13780 24342
rect 13728 24278 13780 24284
rect 13740 23866 13768 24278
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 13832 23186 13860 25774
rect 13924 24274 13952 25774
rect 14108 25158 14136 25842
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 13912 24268 13964 24274
rect 13912 24210 13964 24216
rect 13924 24070 13952 24210
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13820 23180 13872 23186
rect 13820 23122 13872 23128
rect 13648 22066 13768 22094
rect 13636 21412 13688 21418
rect 13636 21354 13688 21360
rect 13452 21004 13504 21010
rect 13452 20946 13504 20952
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13268 20800 13320 20806
rect 13268 20742 13320 20748
rect 13280 19854 13308 20742
rect 13372 20466 13400 20878
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13372 19378 13400 20402
rect 13464 19854 13492 20946
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13464 18290 13492 19790
rect 13648 19446 13676 21354
rect 13636 19440 13688 19446
rect 13636 19382 13688 19388
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13464 17678 13492 18226
rect 13648 17882 13676 18226
rect 13636 17876 13688 17882
rect 13636 17818 13688 17824
rect 13452 17672 13504 17678
rect 13452 17614 13504 17620
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 17270 13124 17478
rect 13084 17264 13136 17270
rect 13084 17206 13136 17212
rect 13740 16250 13768 22066
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 13912 21072 13964 21078
rect 13912 21014 13964 21020
rect 13924 20942 13952 21014
rect 13912 20936 13964 20942
rect 13912 20878 13964 20884
rect 13924 20482 13952 20878
rect 14016 20874 14044 21422
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 14016 20602 14044 20810
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 13924 20454 14044 20482
rect 13912 19712 13964 19718
rect 13912 19654 13964 19660
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13832 18290 13860 18702
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13924 17338 13952 19654
rect 13912 17332 13964 17338
rect 13912 17274 13964 17280
rect 14016 17218 14044 20454
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13924 17190 14044 17218
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13832 16114 13860 17138
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13832 15502 13860 16050
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 13820 15496 13872 15502
rect 13820 15438 13872 15444
rect 13268 15428 13320 15434
rect 13188 15388 13268 15416
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 11150 13032 11494
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12544 9382 12572 9522
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12544 8265 12572 9318
rect 12530 8256 12586 8265
rect 12530 8191 12586 8200
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 11992 6458 12020 6734
rect 11980 6452 12032 6458
rect 11980 6394 12032 6400
rect 11980 6180 12032 6186
rect 11980 6122 12032 6128
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 11900 800 11928 4966
rect 11992 3058 12020 6122
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12084 4690 12112 5170
rect 12072 4684 12124 4690
rect 12072 4626 12124 4632
rect 12084 4078 12112 4626
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12176 800 12204 6054
rect 12452 5914 12480 6734
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12268 4758 12296 4966
rect 12256 4752 12308 4758
rect 12256 4694 12308 4700
rect 12452 800 12480 5102
rect 12544 3534 12572 7482
rect 12728 5710 12756 7686
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12636 3602 12664 3946
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12728 800 12756 4082
rect 12912 3913 12940 6666
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12898 3904 12954 3913
rect 12898 3839 12954 3848
rect 13004 800 13032 6054
rect 13096 4078 13124 15098
rect 13188 13734 13216 15388
rect 13268 15370 13320 15376
rect 13832 14890 13860 15438
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13188 12850 13216 13670
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11762 13308 12038
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13464 11354 13492 11698
rect 13452 11348 13504 11354
rect 13452 11290 13504 11296
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13556 9518 13584 10066
rect 13544 9512 13596 9518
rect 13544 9454 13596 9460
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13188 8974 13216 9318
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 13464 7206 13492 8842
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13452 7200 13504 7206
rect 13452 7142 13504 7148
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13188 3534 13216 7142
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13268 5704 13320 5710
rect 13268 5646 13320 5652
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13188 2854 13216 3470
rect 13176 2848 13228 2854
rect 13176 2790 13228 2796
rect 13280 800 13308 5646
rect 13372 4622 13400 6802
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13464 3126 13492 7142
rect 13556 6798 13584 8298
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13450 2680 13506 2689
rect 13450 2615 13452 2624
rect 13504 2615 13506 2624
rect 13452 2586 13504 2592
rect 13556 800 13584 4626
rect 13648 4010 13676 14214
rect 13924 12434 13952 17190
rect 14108 12442 14136 25094
rect 14372 24812 14424 24818
rect 14372 24754 14424 24760
rect 14188 24744 14240 24750
rect 14188 24686 14240 24692
rect 14200 23866 14228 24686
rect 14384 24410 14412 24754
rect 14372 24404 14424 24410
rect 14372 24346 14424 24352
rect 14844 24206 14872 25094
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14660 23905 14688 24142
rect 14646 23896 14702 23905
rect 14188 23860 14240 23866
rect 14646 23831 14648 23840
rect 14188 23802 14240 23808
rect 14700 23831 14702 23840
rect 14648 23802 14700 23808
rect 14200 22710 14228 23802
rect 14660 23526 14688 23802
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 14372 23180 14424 23186
rect 14372 23122 14424 23128
rect 14188 22704 14240 22710
rect 14188 22646 14240 22652
rect 14280 21344 14332 21350
rect 14280 21286 14332 21292
rect 14292 20942 14320 21286
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14200 19514 14228 19790
rect 14384 19514 14412 23122
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14924 23112 14976 23118
rect 14924 23054 14976 23060
rect 14740 22976 14792 22982
rect 14740 22918 14792 22924
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14464 22432 14516 22438
rect 14464 22374 14516 22380
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14292 17626 14320 19314
rect 14384 18970 14412 19450
rect 14372 18964 14424 18970
rect 14372 18906 14424 18912
rect 14200 17598 14320 17626
rect 14200 17270 14228 17598
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14292 17202 14320 17478
rect 14476 17202 14504 22374
rect 14660 21690 14688 22578
rect 14752 22438 14780 22918
rect 14844 22506 14872 23054
rect 14936 22710 14964 23054
rect 14924 22704 14976 22710
rect 14924 22646 14976 22652
rect 14832 22500 14884 22506
rect 14832 22442 14884 22448
rect 14740 22432 14792 22438
rect 14740 22374 14792 22380
rect 14936 22234 14964 22646
rect 14924 22228 14976 22234
rect 14924 22170 14976 22176
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14188 16516 14240 16522
rect 14188 16458 14240 16464
rect 14200 15978 14228 16458
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14188 15972 14240 15978
rect 14188 15914 14240 15920
rect 14200 15502 14228 15914
rect 14292 15706 14320 16050
rect 14568 16046 14596 17206
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14660 16114 14688 17070
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14556 16040 14608 16046
rect 14556 15982 14608 15988
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14568 15570 14596 15982
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14372 15428 14424 15434
rect 14372 15370 14424 15376
rect 14384 14822 14412 15370
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14384 14414 14412 14758
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14292 13530 14320 13874
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14096 12436 14148 12442
rect 13924 12406 14044 12434
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13832 11762 13860 12310
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13912 9444 13964 9450
rect 13912 9386 13964 9392
rect 13924 8838 13952 9386
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13740 8265 13768 8570
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13726 8256 13782 8265
rect 13726 8191 13782 8200
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13740 2582 13768 7686
rect 13832 5114 13860 8502
rect 13924 8498 13952 8774
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13910 6760 13966 6769
rect 14016 6746 14044 12406
rect 14096 12378 14148 12384
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11082 14228 12038
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 14108 9994 14136 10474
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 14108 7392 14136 9930
rect 14292 9586 14320 13262
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14200 9110 14228 9522
rect 14384 9466 14412 14350
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 14556 13184 14608 13190
rect 14556 13126 14608 13132
rect 14740 13184 14792 13190
rect 14740 13126 14792 13132
rect 14568 12170 14596 13126
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14464 11688 14516 11694
rect 14568 11676 14596 12106
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 11762 14688 12038
rect 14752 11898 14780 13126
rect 14844 12986 14872 13262
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14936 12434 14964 19450
rect 15028 19174 15056 27814
rect 15212 26874 15240 31726
rect 15292 30252 15344 30258
rect 15396 30240 15424 32438
rect 15568 32428 15620 32434
rect 15568 32370 15620 32376
rect 15476 31204 15528 31210
rect 15476 31146 15528 31152
rect 15344 30212 15424 30240
rect 15292 30194 15344 30200
rect 15488 29850 15516 31146
rect 15580 31142 15608 32370
rect 15856 31754 15884 32982
rect 16316 32910 16344 33526
rect 16408 32978 16436 33934
rect 16488 33516 16540 33522
rect 16488 33458 16540 33464
rect 16396 32972 16448 32978
rect 16396 32914 16448 32920
rect 16304 32904 16356 32910
rect 16304 32846 16356 32852
rect 15672 31726 15884 31754
rect 16408 31754 16436 32914
rect 16500 32910 16528 33458
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 16960 32366 16988 34546
rect 16948 32360 17000 32366
rect 16948 32302 17000 32308
rect 17052 32298 17080 35498
rect 17132 33448 17184 33454
rect 17132 33390 17184 33396
rect 17144 32978 17172 33390
rect 17132 32972 17184 32978
rect 17132 32914 17184 32920
rect 17132 32428 17184 32434
rect 17132 32370 17184 32376
rect 17040 32292 17092 32298
rect 17040 32234 17092 32240
rect 17144 32026 17172 32370
rect 17132 32020 17184 32026
rect 17052 31980 17132 32008
rect 16672 31816 16724 31822
rect 16672 31758 16724 31764
rect 16408 31726 16528 31754
rect 15672 31346 15700 31726
rect 16304 31476 16356 31482
rect 16304 31418 16356 31424
rect 15660 31340 15712 31346
rect 15660 31282 15712 31288
rect 15568 31136 15620 31142
rect 15568 31078 15620 31084
rect 15476 29844 15528 29850
rect 15476 29786 15528 29792
rect 15384 29232 15436 29238
rect 15384 29174 15436 29180
rect 15396 29034 15424 29174
rect 15384 29028 15436 29034
rect 15384 28970 15436 28976
rect 15292 28960 15344 28966
rect 15292 28902 15344 28908
rect 15304 28694 15332 28902
rect 15292 28688 15344 28694
rect 15292 28630 15344 28636
rect 15396 28558 15424 28970
rect 15580 28558 15608 31078
rect 15672 28762 15700 31282
rect 15936 31204 15988 31210
rect 15936 31146 15988 31152
rect 15752 30320 15804 30326
rect 15752 30262 15804 30268
rect 15764 29646 15792 30262
rect 15844 30116 15896 30122
rect 15844 30058 15896 30064
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15660 28756 15712 28762
rect 15660 28698 15712 28704
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15568 28552 15620 28558
rect 15568 28494 15620 28500
rect 15568 28416 15620 28422
rect 15568 28358 15620 28364
rect 15580 28082 15608 28358
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 15382 27432 15438 27441
rect 15382 27367 15384 27376
rect 15436 27367 15438 27376
rect 15752 27396 15804 27402
rect 15384 27338 15436 27344
rect 15752 27338 15804 27344
rect 15212 26846 15424 26874
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15212 23798 15240 24550
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 15396 23202 15424 26846
rect 15764 25906 15792 27338
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15856 25786 15884 30058
rect 15764 25758 15884 25786
rect 15568 25696 15620 25702
rect 15568 25638 15620 25644
rect 15580 25226 15608 25638
rect 15568 25220 15620 25226
rect 15568 25162 15620 25168
rect 15580 24342 15608 25162
rect 15568 24336 15620 24342
rect 15568 24278 15620 24284
rect 15212 23174 15424 23202
rect 15212 22930 15240 23174
rect 15384 22976 15436 22982
rect 15212 22902 15332 22930
rect 15384 22918 15436 22924
rect 15200 22228 15252 22234
rect 15200 22170 15252 22176
rect 15212 22030 15240 22170
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15212 17678 15240 18022
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 15028 13818 15056 16118
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15120 14958 15148 15438
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15120 13938 15148 14894
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15028 13790 15148 13818
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 14844 12406 14964 12434
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14516 11648 14596 11676
rect 14464 11630 14516 11636
rect 14464 9580 14516 9586
rect 14464 9522 14516 9528
rect 14292 9438 14412 9466
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14200 8294 14228 8774
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14188 7404 14240 7410
rect 14108 7364 14188 7392
rect 14188 7346 14240 7352
rect 14096 7200 14148 7206
rect 14096 7142 14148 7148
rect 14108 7002 14136 7142
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 13966 6718 14044 6746
rect 14096 6724 14148 6730
rect 13910 6695 13966 6704
rect 13924 6662 13952 6695
rect 14200 6712 14228 7346
rect 14148 6684 14228 6712
rect 14096 6666 14148 6672
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 14004 6656 14056 6662
rect 14004 6598 14056 6604
rect 14016 6322 14044 6598
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14096 5704 14148 5710
rect 14096 5646 14148 5652
rect 13832 5086 14044 5114
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 13832 800 13860 4966
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13924 3602 13952 4422
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 14016 3058 14044 5086
rect 14108 4146 14136 5646
rect 14292 5370 14320 9438
rect 14372 9376 14424 9382
rect 14372 9318 14424 9324
rect 14384 8974 14412 9318
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14476 8838 14504 9522
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14752 7750 14780 8434
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14568 7342 14596 7373
rect 14556 7336 14608 7342
rect 14554 7304 14556 7313
rect 14608 7304 14610 7313
rect 14554 7239 14610 7248
rect 14568 6798 14596 7239
rect 14556 6792 14608 6798
rect 14556 6734 14608 6740
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 14568 5642 14596 6734
rect 14660 6458 14688 6734
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14752 5658 14780 7686
rect 14844 6905 14872 12406
rect 15028 12374 15056 13262
rect 15120 13190 15148 13790
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15120 12850 15148 13126
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15016 12368 15068 12374
rect 15016 12310 15068 12316
rect 15120 12238 15148 12582
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15212 12170 15240 12242
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14936 8294 14964 11018
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 10810 15056 10950
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15016 8356 15068 8362
rect 15016 8298 15068 8304
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14830 6896 14886 6905
rect 14830 6831 14886 6840
rect 14936 6798 14964 7346
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14936 6662 14964 6734
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14936 5710 14964 6598
rect 14924 5704 14976 5710
rect 14830 5672 14886 5681
rect 14556 5636 14608 5642
rect 14752 5630 14830 5658
rect 14924 5646 14976 5652
rect 14830 5607 14886 5616
rect 14556 5578 14608 5584
rect 14844 5574 14872 5607
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14280 5364 14332 5370
rect 14280 5306 14332 5312
rect 15028 5234 15056 8298
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14096 3392 14148 3398
rect 14094 3360 14096 3369
rect 14148 3360 14150 3369
rect 14094 3295 14150 3304
rect 14200 3210 14228 4966
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14108 3182 14228 3210
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 14016 2106 14044 2382
rect 14004 2100 14056 2106
rect 14004 2042 14056 2048
rect 14108 800 14136 3182
rect 14292 2774 14320 4558
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14200 2746 14320 2774
rect 14200 800 14228 2746
rect 14384 800 14412 3674
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14476 800 14504 3470
rect 14554 3224 14610 3233
rect 14554 3159 14556 3168
rect 14608 3159 14610 3168
rect 14556 3130 14608 3136
rect 14554 2680 14610 2689
rect 14554 2615 14556 2624
rect 14608 2615 14610 2624
rect 14556 2586 14608 2592
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14568 2038 14596 2382
rect 14556 2032 14608 2038
rect 14556 1974 14608 1980
rect 14660 800 14688 3878
rect 14752 800 14780 5170
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14844 3466 14872 4966
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 15120 3058 15148 7822
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15120 2854 15148 2994
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15108 2848 15160 2854
rect 15108 2790 15160 2796
rect 14924 2508 14976 2514
rect 14924 2450 14976 2456
rect 14936 800 14964 2450
rect 15028 800 15056 2790
rect 15212 800 15240 3946
rect 15304 3194 15332 22902
rect 15396 21554 15424 22918
rect 15660 21888 15712 21894
rect 15660 21830 15712 21836
rect 15764 21842 15792 25758
rect 15948 25294 15976 31146
rect 16316 31142 16344 31418
rect 16304 31136 16356 31142
rect 16304 31078 16356 31084
rect 16212 30592 16264 30598
rect 16212 30534 16264 30540
rect 16224 30326 16252 30534
rect 16212 30320 16264 30326
rect 16212 30262 16264 30268
rect 16212 28960 16264 28966
rect 16212 28902 16264 28908
rect 16224 28490 16252 28902
rect 16212 28484 16264 28490
rect 16212 28426 16264 28432
rect 16224 28218 16252 28426
rect 16212 28212 16264 28218
rect 16212 28154 16264 28160
rect 16212 27124 16264 27130
rect 16212 27066 16264 27072
rect 16028 25764 16080 25770
rect 16028 25706 16080 25712
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15856 24614 15884 25094
rect 15844 24608 15896 24614
rect 15844 24550 15896 24556
rect 15856 23050 15884 24550
rect 15948 24410 15976 25230
rect 16040 25226 16068 25706
rect 16028 25220 16080 25226
rect 16028 25162 16080 25168
rect 15936 24404 15988 24410
rect 15936 24346 15988 24352
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 15844 23044 15896 23050
rect 15844 22986 15896 22992
rect 16132 22778 16160 23054
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15856 22001 15884 22034
rect 16120 22024 16172 22030
rect 15842 21992 15898 22001
rect 16120 21966 16172 21972
rect 15842 21927 15898 21936
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15568 20324 15620 20330
rect 15568 20266 15620 20272
rect 15580 20058 15608 20266
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15396 15502 15424 16390
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 11286 15516 11494
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15672 11014 15700 21830
rect 15764 21814 15884 21842
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15764 19854 15792 20402
rect 15856 19854 15884 21814
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 15752 19848 15804 19854
rect 15752 19790 15804 19796
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15764 17202 15792 19790
rect 15856 19174 15884 19790
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18086 15884 19110
rect 15844 18080 15896 18086
rect 15844 18022 15896 18028
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15948 17134 15976 21626
rect 16028 20868 16080 20874
rect 16028 20810 16080 20816
rect 16040 20602 16068 20810
rect 16028 20596 16080 20602
rect 16028 20538 16080 20544
rect 15936 17128 15988 17134
rect 15936 17070 15988 17076
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15764 16590 15792 16730
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15948 16250 15976 16526
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 16040 12986 16068 20538
rect 16132 19922 16160 21966
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 16132 16182 16160 16526
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15764 12170 15792 12922
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15752 12164 15804 12170
rect 15752 12106 15804 12112
rect 16040 11558 16068 12174
rect 16132 11558 16160 12242
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16040 11064 16068 11494
rect 16040 11036 16160 11064
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15568 9376 15620 9382
rect 15568 9318 15620 9324
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15488 6769 15516 6802
rect 15474 6760 15530 6769
rect 15474 6695 15530 6704
rect 15476 5704 15528 5710
rect 15474 5672 15476 5681
rect 15528 5672 15530 5681
rect 15474 5607 15530 5616
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15304 800 15332 2994
rect 15396 800 15424 4558
rect 15580 2938 15608 9318
rect 15948 8974 15976 9318
rect 16132 9110 16160 11036
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15672 7546 15700 7754
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15948 7274 15976 8910
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 16040 6458 16068 6734
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 15752 6180 15804 6186
rect 15752 6122 15804 6128
rect 15764 5778 15792 6122
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 15844 5092 15896 5098
rect 15844 5034 15896 5040
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15488 2910 15608 2938
rect 15488 2446 15516 2910
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15580 800 15608 2790
rect 15672 800 15700 4966
rect 15856 3602 15884 5034
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15844 3596 15896 3602
rect 15844 3538 15896 3544
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15764 1442 15792 3470
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15856 2446 15884 2586
rect 15844 2440 15896 2446
rect 15844 2382 15896 2388
rect 15856 1902 15884 2382
rect 15844 1896 15896 1902
rect 15844 1838 15896 1844
rect 15764 1414 15884 1442
rect 15856 800 15884 1414
rect 15948 800 15976 4558
rect 16132 4078 16160 5510
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 16120 4072 16172 4078
rect 16120 4014 16172 4020
rect 16040 2774 16068 4014
rect 16118 3768 16174 3777
rect 16118 3703 16120 3712
rect 16172 3703 16174 3712
rect 16120 3674 16172 3680
rect 16118 3224 16174 3233
rect 16118 3159 16120 3168
rect 16172 3159 16174 3168
rect 16120 3130 16172 3136
rect 16040 2746 16160 2774
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 16040 1306 16068 2246
rect 16132 1442 16160 2746
rect 16224 2582 16252 27066
rect 16316 24614 16344 31078
rect 16500 30734 16528 31726
rect 16488 30728 16540 30734
rect 16488 30670 16540 30676
rect 16500 30258 16528 30670
rect 16684 30666 16712 31758
rect 17052 30938 17080 31980
rect 17132 31962 17184 31968
rect 17040 30932 17092 30938
rect 17040 30874 17092 30880
rect 16764 30864 16816 30870
rect 16764 30806 16816 30812
rect 16672 30660 16724 30666
rect 16672 30602 16724 30608
rect 16672 30388 16724 30394
rect 16592 30348 16672 30376
rect 16488 30252 16540 30258
rect 16488 30194 16540 30200
rect 16396 30048 16448 30054
rect 16396 29990 16448 29996
rect 16304 24608 16356 24614
rect 16304 24550 16356 24556
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16316 22506 16344 23258
rect 16304 22500 16356 22506
rect 16304 22442 16356 22448
rect 16316 22030 16344 22442
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16408 21706 16436 29990
rect 16592 26382 16620 30348
rect 16672 30330 16724 30336
rect 16672 28008 16724 28014
rect 16672 27950 16724 27956
rect 16580 26376 16632 26382
rect 16580 26318 16632 26324
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 16500 22642 16528 24618
rect 16592 24070 16620 24754
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16316 21690 16436 21706
rect 16304 21684 16436 21690
rect 16356 21678 16436 21684
rect 16304 21626 16356 21632
rect 16396 21616 16448 21622
rect 16396 21558 16448 21564
rect 16304 21548 16356 21554
rect 16304 21490 16356 21496
rect 16316 21078 16344 21490
rect 16304 21072 16356 21078
rect 16304 21014 16356 21020
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16316 16658 16344 16730
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16408 13326 16436 21558
rect 16500 21554 16528 22578
rect 16592 22234 16620 24006
rect 16684 22574 16712 27950
rect 16776 27606 16804 30806
rect 17040 30728 17092 30734
rect 17040 30670 17092 30676
rect 17052 30394 17080 30670
rect 17040 30388 17092 30394
rect 17040 30330 17092 30336
rect 16948 29640 17000 29646
rect 16948 29582 17000 29588
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16868 27674 16896 27814
rect 16856 27668 16908 27674
rect 16856 27610 16908 27616
rect 16764 27600 16816 27606
rect 16764 27542 16816 27548
rect 16776 26450 16804 27542
rect 16960 26874 16988 29582
rect 17040 27464 17092 27470
rect 17040 27406 17092 27412
rect 16868 26846 16988 26874
rect 16764 26444 16816 26450
rect 16764 26386 16816 26392
rect 16868 23322 16896 26846
rect 17052 26382 17080 27406
rect 17236 27130 17264 41386
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17328 34066 17356 35022
rect 17316 34060 17368 34066
rect 17316 34002 17368 34008
rect 17328 32570 17356 34002
rect 17316 32564 17368 32570
rect 17316 32506 17368 32512
rect 17316 32360 17368 32366
rect 17316 32302 17368 32308
rect 17328 31958 17356 32302
rect 17316 31952 17368 31958
rect 17316 31894 17368 31900
rect 17328 30870 17356 31894
rect 17316 30864 17368 30870
rect 17316 30806 17368 30812
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 17224 27124 17276 27130
rect 17224 27066 17276 27072
rect 17328 27010 17356 30534
rect 17144 26982 17356 27010
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 16948 25220 17000 25226
rect 16948 25162 17000 25168
rect 16960 24342 16988 25162
rect 16948 24336 17000 24342
rect 17000 24296 17080 24324
rect 16948 24278 17000 24284
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16684 22094 16712 22510
rect 16592 22066 16712 22094
rect 16868 22094 16896 23258
rect 16868 22066 16988 22094
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16500 21146 16528 21490
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16500 20534 16528 21082
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16500 19378 16528 20470
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16500 17746 16528 19314
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16592 14618 16620 22066
rect 16960 22030 16988 22066
rect 16948 22024 17000 22030
rect 16946 21992 16948 22001
rect 17000 21992 17002 22001
rect 16946 21927 17002 21936
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 16960 21622 16988 21830
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16960 20806 16988 21286
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16960 20602 16988 20742
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16764 19372 16816 19378
rect 16764 19314 16816 19320
rect 16776 18970 16804 19314
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 17052 18766 17080 24296
rect 17144 22098 17172 26982
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17132 22092 17184 22098
rect 17132 22034 17184 22040
rect 17224 22024 17276 22030
rect 17224 21966 17276 21972
rect 17236 21554 17264 21966
rect 17224 21548 17276 21554
rect 17224 21490 17276 21496
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 16776 18358 16804 18702
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 17040 17264 17092 17270
rect 17040 17206 17092 17212
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16684 15094 16712 17138
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 16764 16720 16816 16726
rect 16762 16688 16764 16697
rect 16816 16688 16818 16697
rect 16762 16623 16818 16632
rect 16960 16590 16988 17002
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16776 16250 16804 16526
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16960 15366 16988 16050
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16408 12714 16436 13262
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16684 12782 16712 13194
rect 16868 12918 16896 14894
rect 16960 14550 16988 15302
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 16856 12912 16908 12918
rect 16856 12854 16908 12860
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16684 12374 16712 12718
rect 16672 12368 16724 12374
rect 16672 12310 16724 12316
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16500 10266 16528 10950
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16592 8090 16620 12106
rect 16684 11150 16712 12310
rect 16868 12102 16896 12854
rect 17052 12434 17080 17206
rect 17224 16448 17276 16454
rect 17224 16390 17276 16396
rect 17236 15094 17264 16390
rect 17224 15088 17276 15094
rect 17224 15030 17276 15036
rect 17052 12406 17172 12434
rect 17144 12306 17172 12406
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16868 11830 16896 12038
rect 17144 11898 17172 12242
rect 17328 11898 17356 26250
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 16856 11824 16908 11830
rect 16856 11766 16908 11772
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16672 8832 16724 8838
rect 16672 8774 16724 8780
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16592 6322 16620 8026
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16408 4049 16436 4218
rect 16684 4162 16712 8774
rect 16776 8566 16804 9590
rect 16868 9042 16896 11766
rect 17328 10742 17356 11834
rect 17316 10736 17368 10742
rect 17316 10678 17368 10684
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17144 9994 17172 10610
rect 17132 9988 17184 9994
rect 17132 9930 17184 9936
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 16856 9036 16908 9042
rect 16856 8978 16908 8984
rect 17052 8838 17080 9046
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7478 16804 7686
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16868 6905 16896 8570
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16854 6896 16910 6905
rect 16854 6831 16910 6840
rect 17052 6254 17080 7346
rect 17040 6248 17092 6254
rect 17040 6190 17092 6196
rect 17052 5642 17080 6190
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 16592 4134 16712 4162
rect 16394 4040 16450 4049
rect 16394 3975 16450 3984
rect 16592 3534 16620 4134
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16684 3398 16712 3946
rect 17052 3754 17080 4626
rect 17130 4040 17186 4049
rect 17130 3975 17186 3984
rect 16776 3726 17080 3754
rect 17144 3738 17172 3975
rect 17132 3732 17184 3738
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16396 2032 16448 2038
rect 16396 1974 16448 1980
rect 16132 1414 16252 1442
rect 16040 1278 16160 1306
rect 16132 800 16160 1278
rect 16224 800 16252 1414
rect 16408 800 16436 1974
rect 16500 800 16528 2858
rect 16684 800 16712 2994
rect 16776 800 16804 3726
rect 17132 3674 17184 3680
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 16868 3534 16896 3606
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 16868 1442 16896 3470
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16960 1850 16988 3334
rect 17236 3058 17264 9318
rect 17316 8900 17368 8906
rect 17316 8842 17368 8848
rect 17328 8634 17356 8842
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17224 3052 17276 3058
rect 17224 2994 17276 3000
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17224 2372 17276 2378
rect 17224 2314 17276 2320
rect 16960 1822 17172 1850
rect 17144 1442 17172 1822
rect 16868 1414 16988 1442
rect 16960 800 16988 1414
rect 17052 1414 17172 1442
rect 17052 800 17080 1414
rect 17236 800 17264 2314
rect 17328 800 17356 2926
rect 17420 2650 17448 41386
rect 17500 40928 17552 40934
rect 17500 40870 17552 40876
rect 17512 40526 17540 40870
rect 17500 40520 17552 40526
rect 17500 40462 17552 40468
rect 17512 37874 17540 40462
rect 17500 37868 17552 37874
rect 17500 37810 17552 37816
rect 17500 37664 17552 37670
rect 17500 37606 17552 37612
rect 17512 31754 17540 37606
rect 17592 35012 17644 35018
rect 17592 34954 17644 34960
rect 17604 34746 17632 34954
rect 17592 34740 17644 34746
rect 17592 34682 17644 34688
rect 17592 33992 17644 33998
rect 17592 33934 17644 33940
rect 17604 33590 17632 33934
rect 17592 33584 17644 33590
rect 17592 33526 17644 33532
rect 17604 33318 17632 33526
rect 17592 33312 17644 33318
rect 17592 33254 17644 33260
rect 17696 32910 17724 41414
rect 17776 40996 17828 41002
rect 17776 40938 17828 40944
rect 17788 39370 17816 40938
rect 18432 40458 18460 41482
rect 18604 40928 18656 40934
rect 18604 40870 18656 40876
rect 18420 40452 18472 40458
rect 18420 40394 18472 40400
rect 18432 40118 18460 40394
rect 18420 40112 18472 40118
rect 18420 40054 18472 40060
rect 18328 39976 18380 39982
rect 18328 39918 18380 39924
rect 18340 39438 18368 39918
rect 18328 39432 18380 39438
rect 18328 39374 18380 39380
rect 17776 39364 17828 39370
rect 17776 39306 17828 39312
rect 18144 38480 18196 38486
rect 18144 38422 18196 38428
rect 18156 36786 18184 38422
rect 18328 38004 18380 38010
rect 18328 37946 18380 37952
rect 18340 37806 18368 37946
rect 18512 37868 18564 37874
rect 18512 37810 18564 37816
rect 18328 37800 18380 37806
rect 18328 37742 18380 37748
rect 18340 37194 18368 37742
rect 18524 37262 18552 37810
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 18328 37188 18380 37194
rect 18328 37130 18380 37136
rect 18236 36848 18288 36854
rect 18236 36790 18288 36796
rect 18144 36780 18196 36786
rect 18064 36740 18144 36768
rect 18064 36378 18092 36740
rect 18144 36722 18196 36728
rect 18144 36644 18196 36650
rect 18144 36586 18196 36592
rect 18052 36372 18104 36378
rect 18052 36314 18104 36320
rect 18052 35692 18104 35698
rect 18052 35634 18104 35640
rect 17960 35488 18012 35494
rect 17960 35430 18012 35436
rect 17972 34610 18000 35430
rect 18064 35290 18092 35634
rect 18052 35284 18104 35290
rect 18052 35226 18104 35232
rect 18064 34678 18092 35226
rect 18052 34672 18104 34678
rect 18052 34614 18104 34620
rect 18156 34610 18184 36586
rect 18248 36106 18276 36790
rect 18236 36100 18288 36106
rect 18236 36042 18288 36048
rect 18248 35766 18276 36042
rect 18236 35760 18288 35766
rect 18236 35702 18288 35708
rect 18236 35012 18288 35018
rect 18236 34954 18288 34960
rect 17868 34604 17920 34610
rect 17868 34546 17920 34552
rect 17960 34604 18012 34610
rect 17960 34546 18012 34552
rect 18144 34604 18196 34610
rect 18144 34546 18196 34552
rect 17880 34202 17908 34546
rect 17868 34196 17920 34202
rect 17868 34138 17920 34144
rect 18156 33998 18184 34546
rect 17868 33992 17920 33998
rect 17868 33934 17920 33940
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 17880 33658 17908 33934
rect 17868 33652 17920 33658
rect 17868 33594 17920 33600
rect 17960 33516 18012 33522
rect 17960 33458 18012 33464
rect 17592 32904 17644 32910
rect 17592 32846 17644 32852
rect 17684 32904 17736 32910
rect 17684 32846 17736 32852
rect 17604 32502 17632 32846
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17592 32496 17644 32502
rect 17592 32438 17644 32444
rect 17604 32366 17632 32438
rect 17592 32360 17644 32366
rect 17592 32302 17644 32308
rect 17512 31726 17632 31754
rect 17500 27396 17552 27402
rect 17500 27338 17552 27344
rect 17512 26586 17540 27338
rect 17500 26580 17552 26586
rect 17500 26522 17552 26528
rect 17512 25906 17540 26522
rect 17500 25900 17552 25906
rect 17500 25842 17552 25848
rect 17604 22166 17632 31726
rect 17776 27940 17828 27946
rect 17776 27882 17828 27888
rect 17788 27470 17816 27882
rect 17776 27464 17828 27470
rect 17776 27406 17828 27412
rect 17788 27130 17816 27406
rect 17776 27124 17828 27130
rect 17776 27066 17828 27072
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17696 26042 17724 26930
rect 17776 26376 17828 26382
rect 17776 26318 17828 26324
rect 17684 26036 17736 26042
rect 17684 25978 17736 25984
rect 17788 24750 17816 26318
rect 17776 24744 17828 24750
rect 17776 24686 17828 24692
rect 17788 23594 17816 24686
rect 17776 23588 17828 23594
rect 17776 23530 17828 23536
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17592 22160 17644 22166
rect 17592 22102 17644 22108
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17512 21146 17540 21966
rect 17592 21344 17644 21350
rect 17592 21286 17644 21292
rect 17500 21140 17552 21146
rect 17500 21082 17552 21088
rect 17604 20942 17632 21286
rect 17592 20936 17644 20942
rect 17592 20878 17644 20884
rect 17592 20256 17644 20262
rect 17592 20198 17644 20204
rect 17604 10810 17632 20198
rect 17696 13462 17724 22170
rect 17880 20262 17908 32710
rect 17972 31890 18000 33458
rect 18156 33402 18184 33934
rect 18064 33374 18184 33402
rect 18064 33114 18092 33374
rect 18248 33318 18276 34954
rect 18340 34746 18368 37130
rect 18328 34740 18380 34746
rect 18328 34682 18380 34688
rect 18524 33862 18552 37198
rect 18616 36038 18644 40870
rect 18800 37369 18828 56102
rect 18892 55214 18920 56374
rect 18972 56364 19024 56370
rect 18972 56306 19024 56312
rect 18984 55350 19012 56306
rect 19260 55962 19288 57394
rect 19352 56506 19380 57394
rect 20076 57248 20128 57254
rect 20074 57216 20076 57225
rect 20128 57216 20130 57225
rect 20074 57151 20130 57160
rect 19432 56976 19484 56982
rect 19432 56918 19484 56924
rect 19340 56500 19392 56506
rect 19340 56442 19392 56448
rect 19444 55962 19472 56918
rect 20088 56846 20116 57151
rect 20076 56840 20128 56846
rect 20076 56782 20128 56788
rect 19984 56704 20036 56710
rect 19984 56646 20036 56652
rect 20720 56704 20772 56710
rect 20720 56646 20772 56652
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 19996 56370 20024 56646
rect 20732 56370 20760 56646
rect 22204 56506 22232 57394
rect 22284 56704 22336 56710
rect 22284 56646 22336 56652
rect 22192 56500 22244 56506
rect 22192 56442 22244 56448
rect 22296 56370 22324 56646
rect 24412 56506 24440 57394
rect 25136 56704 25188 56710
rect 25134 56672 25136 56681
rect 25188 56672 25190 56681
rect 25134 56607 25190 56616
rect 24400 56500 24452 56506
rect 24400 56442 24452 56448
rect 19984 56364 20036 56370
rect 19984 56306 20036 56312
rect 20536 56364 20588 56370
rect 20536 56306 20588 56312
rect 20720 56364 20772 56370
rect 20720 56306 20772 56312
rect 21088 56364 21140 56370
rect 21088 56306 21140 56312
rect 21640 56364 21692 56370
rect 21640 56306 21692 56312
rect 22284 56364 22336 56370
rect 22284 56306 22336 56312
rect 22560 56364 22612 56370
rect 22560 56306 22612 56312
rect 23940 56364 23992 56370
rect 23940 56306 23992 56312
rect 24952 56364 25004 56370
rect 24952 56306 25004 56312
rect 19248 55956 19300 55962
rect 19248 55898 19300 55904
rect 19432 55956 19484 55962
rect 19432 55898 19484 55904
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 19156 55412 19208 55418
rect 19156 55354 19208 55360
rect 18972 55344 19024 55350
rect 18970 55312 18972 55321
rect 19024 55312 19026 55321
rect 18970 55247 19026 55256
rect 18892 55186 19012 55214
rect 18786 37360 18842 37369
rect 18786 37295 18842 37304
rect 18696 37120 18748 37126
rect 18696 37062 18748 37068
rect 18604 36032 18656 36038
rect 18604 35974 18656 35980
rect 18616 34898 18644 35974
rect 18708 35018 18736 37062
rect 18696 35012 18748 35018
rect 18696 34954 18748 34960
rect 18616 34870 18736 34898
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18604 33584 18656 33590
rect 18604 33526 18656 33532
rect 18236 33312 18288 33318
rect 18236 33254 18288 33260
rect 18052 33108 18104 33114
rect 18052 33050 18104 33056
rect 17960 31884 18012 31890
rect 17960 31826 18012 31832
rect 17960 30252 18012 30258
rect 17960 30194 18012 30200
rect 17972 29850 18000 30194
rect 17960 29844 18012 29850
rect 17960 29786 18012 29792
rect 18248 28490 18276 33254
rect 18616 32978 18644 33526
rect 18604 32972 18656 32978
rect 18604 32914 18656 32920
rect 18420 32768 18472 32774
rect 18420 32710 18472 32716
rect 18432 32586 18460 32710
rect 18432 32558 18552 32586
rect 18616 32570 18644 32914
rect 18524 32502 18552 32558
rect 18604 32564 18656 32570
rect 18604 32506 18656 32512
rect 18512 32496 18564 32502
rect 18512 32438 18564 32444
rect 18328 30864 18380 30870
rect 18328 30806 18380 30812
rect 18340 30326 18368 30806
rect 18512 30660 18564 30666
rect 18512 30602 18564 30608
rect 18524 30394 18552 30602
rect 18604 30592 18656 30598
rect 18604 30534 18656 30540
rect 18512 30388 18564 30394
rect 18512 30330 18564 30336
rect 18328 30320 18380 30326
rect 18328 30262 18380 30268
rect 18616 29646 18644 30534
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18236 28484 18288 28490
rect 18236 28426 18288 28432
rect 18420 28484 18472 28490
rect 18420 28426 18472 28432
rect 17960 27872 18012 27878
rect 17960 27814 18012 27820
rect 17972 25430 18000 27814
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18144 26308 18196 26314
rect 18144 26250 18196 26256
rect 18052 26240 18104 26246
rect 18052 26182 18104 26188
rect 18064 25906 18092 26182
rect 18052 25900 18104 25906
rect 18052 25842 18104 25848
rect 18064 25498 18092 25842
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 17960 25424 18012 25430
rect 17960 25366 18012 25372
rect 18064 24274 18092 25434
rect 18156 25294 18184 26250
rect 18248 26042 18276 26318
rect 18236 26036 18288 26042
rect 18236 25978 18288 25984
rect 18432 25974 18460 28426
rect 18708 26382 18736 34870
rect 18788 31136 18840 31142
rect 18788 31078 18840 31084
rect 18800 29578 18828 31078
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18788 29572 18840 29578
rect 18788 29514 18840 29520
rect 18788 29300 18840 29306
rect 18788 29242 18840 29248
rect 18696 26376 18748 26382
rect 18696 26318 18748 26324
rect 18420 25968 18472 25974
rect 18420 25910 18472 25916
rect 18604 25968 18656 25974
rect 18604 25910 18656 25916
rect 18236 25424 18288 25430
rect 18236 25366 18288 25372
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 18052 24268 18104 24274
rect 18052 24210 18104 24216
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17972 23050 18000 23666
rect 17960 23044 18012 23050
rect 17960 22986 18012 22992
rect 17972 20874 18000 22986
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18064 21690 18092 21966
rect 18052 21684 18104 21690
rect 18052 21626 18104 21632
rect 18052 21344 18104 21350
rect 18052 21286 18104 21292
rect 18064 20942 18092 21286
rect 18156 21010 18184 25230
rect 18248 24410 18276 25366
rect 18616 25158 18644 25910
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 18420 24200 18472 24206
rect 18420 24142 18472 24148
rect 18236 24132 18288 24138
rect 18236 24074 18288 24080
rect 18248 23866 18276 24074
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18432 21894 18460 24142
rect 18420 21888 18472 21894
rect 18420 21830 18472 21836
rect 18144 21004 18196 21010
rect 18144 20946 18196 20952
rect 18052 20936 18104 20942
rect 18052 20878 18104 20884
rect 17960 20868 18012 20874
rect 17960 20810 18012 20816
rect 17972 20330 18000 20810
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 18052 19984 18104 19990
rect 18052 19926 18104 19932
rect 18064 19174 18092 19926
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 17776 18828 17828 18834
rect 17776 18770 17828 18776
rect 17788 16522 17816 18770
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17880 18358 17908 18702
rect 17868 18352 17920 18358
rect 18064 18340 18092 19110
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 17868 18294 17920 18300
rect 17972 18312 18092 18340
rect 17972 18222 18000 18312
rect 18156 18222 18184 18702
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17880 18034 17908 18090
rect 17880 18006 18000 18034
rect 17972 17270 18000 18006
rect 17960 17264 18012 17270
rect 18012 17212 18092 17218
rect 17960 17206 18092 17212
rect 17972 17190 18092 17206
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17972 16658 18000 17002
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17776 16516 17828 16522
rect 17776 16458 17828 16464
rect 18064 16454 18092 17190
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18248 16250 18276 16526
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 18248 14890 18276 16050
rect 18524 15162 18552 24550
rect 18616 23866 18644 25094
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18800 22778 18828 29242
rect 18892 29034 18920 29582
rect 18880 29028 18932 29034
rect 18880 28970 18932 28976
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 18616 22030 18644 22714
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18800 22234 18828 22578
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18604 22024 18656 22030
rect 18604 21966 18656 21972
rect 18788 20528 18840 20534
rect 18788 20470 18840 20476
rect 18800 20262 18828 20470
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18800 18358 18828 18566
rect 18788 18352 18840 18358
rect 18788 18294 18840 18300
rect 18602 18048 18658 18057
rect 18602 17983 18658 17992
rect 18512 15156 18564 15162
rect 18512 15098 18564 15104
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 17684 13456 17736 13462
rect 17684 13398 17736 13404
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17696 9674 17724 13398
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18052 12844 18104 12850
rect 18052 12786 18104 12792
rect 18064 12170 18092 12786
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 18156 11354 18184 12174
rect 18432 11762 18460 12582
rect 18524 12238 18552 13126
rect 18616 12345 18644 17983
rect 18892 17202 18920 28970
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18892 17066 18920 17138
rect 18880 17060 18932 17066
rect 18880 17002 18932 17008
rect 18984 16946 19012 55186
rect 19064 38208 19116 38214
rect 19064 38150 19116 38156
rect 19076 37874 19104 38150
rect 19064 37868 19116 37874
rect 19064 37810 19116 37816
rect 19076 36854 19104 37810
rect 19064 36848 19116 36854
rect 19064 36790 19116 36796
rect 19064 33924 19116 33930
rect 19064 33866 19116 33872
rect 19076 33658 19104 33866
rect 19064 33652 19116 33658
rect 19064 33594 19116 33600
rect 19168 31754 19196 55354
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19432 41540 19484 41546
rect 19432 41482 19484 41488
rect 19340 41472 19392 41478
rect 19338 41440 19340 41449
rect 19392 41440 19394 41449
rect 19338 41375 19394 41384
rect 19444 41290 19472 41482
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19260 41262 19472 41290
rect 19260 40372 19288 41262
rect 19338 41168 19394 41177
rect 19524 41132 19576 41138
rect 19338 41103 19394 41112
rect 19352 40526 19380 41103
rect 19444 41092 19524 41120
rect 19340 40520 19392 40526
rect 19340 40462 19392 40468
rect 19260 40344 19380 40372
rect 19248 40112 19300 40118
rect 19248 40054 19300 40060
rect 19260 37210 19288 40054
rect 19352 39642 19380 40344
rect 19444 39982 19472 41092
rect 19524 41074 19576 41080
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19432 39976 19484 39982
rect 19432 39918 19484 39924
rect 19340 39636 19392 39642
rect 19340 39578 19392 39584
rect 19352 38010 19380 39578
rect 19444 39438 19472 39918
rect 19432 39432 19484 39438
rect 19432 39374 19484 39380
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19432 38276 19484 38282
rect 19432 38218 19484 38224
rect 19340 38004 19392 38010
rect 19340 37946 19392 37952
rect 19260 37182 19380 37210
rect 19352 37126 19380 37182
rect 19340 37120 19392 37126
rect 19340 37062 19392 37068
rect 19248 34604 19300 34610
rect 19248 34546 19300 34552
rect 19260 33862 19288 34546
rect 19352 33998 19380 37062
rect 19444 36922 19472 38218
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19432 36916 19484 36922
rect 19432 36858 19484 36864
rect 19432 36576 19484 36582
rect 19432 36518 19484 36524
rect 19444 34950 19472 36518
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19432 34944 19484 34950
rect 19432 34886 19484 34892
rect 19444 34626 19472 34886
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19800 34672 19852 34678
rect 19444 34610 19564 34626
rect 19800 34614 19852 34620
rect 19444 34604 19576 34610
rect 19444 34598 19524 34604
rect 19524 34546 19576 34552
rect 19432 34536 19484 34542
rect 19432 34478 19484 34484
rect 19340 33992 19392 33998
rect 19340 33934 19392 33940
rect 19248 33856 19300 33862
rect 19248 33798 19300 33804
rect 19352 33590 19380 33934
rect 19340 33584 19392 33590
rect 19340 33526 19392 33532
rect 19444 32434 19472 34478
rect 19536 33930 19564 34546
rect 19812 33998 19840 34614
rect 19800 33992 19852 33998
rect 19800 33934 19852 33940
rect 19524 33924 19576 33930
rect 19524 33866 19576 33872
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19708 33516 19760 33522
rect 19708 33458 19760 33464
rect 19720 33318 19748 33458
rect 19708 33312 19760 33318
rect 19708 33254 19760 33260
rect 19720 32842 19748 33254
rect 19708 32836 19760 32842
rect 19708 32778 19760 32784
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19248 32428 19300 32434
rect 19248 32370 19300 32376
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19076 31726 19196 31754
rect 19076 22094 19104 31726
rect 19260 31278 19288 32370
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31340 19484 31346
rect 19432 31282 19484 31288
rect 19248 31272 19300 31278
rect 19248 31214 19300 31220
rect 19260 30870 19288 31214
rect 19248 30864 19300 30870
rect 19248 30806 19300 30812
rect 19444 30394 19472 31282
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19156 30388 19208 30394
rect 19156 30330 19208 30336
rect 19432 30388 19484 30394
rect 19432 30330 19484 30336
rect 19168 29170 19196 30330
rect 19248 30184 19300 30190
rect 19248 30126 19300 30132
rect 19260 29306 19288 30126
rect 19892 30116 19944 30122
rect 19892 30058 19944 30064
rect 19904 29578 19932 30058
rect 19432 29572 19484 29578
rect 19432 29514 19484 29520
rect 19892 29572 19944 29578
rect 19892 29514 19944 29520
rect 19248 29300 19300 29306
rect 19248 29242 19300 29248
rect 19156 29164 19208 29170
rect 19156 29106 19208 29112
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19352 28966 19380 29106
rect 19340 28960 19392 28966
rect 19340 28902 19392 28908
rect 19352 28082 19380 28902
rect 19444 28762 19472 29514
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 28756 19484 28762
rect 19432 28698 19484 28704
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 19260 26586 19288 26930
rect 19340 26784 19392 26790
rect 19392 26732 19472 26738
rect 19340 26726 19472 26732
rect 19352 26710 19472 26726
rect 19248 26580 19300 26586
rect 19248 26522 19300 26528
rect 19444 25906 19472 26710
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19248 25900 19300 25906
rect 19248 25842 19300 25848
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 19260 25770 19288 25842
rect 19248 25764 19300 25770
rect 19248 25706 19300 25712
rect 19156 25152 19208 25158
rect 19156 25094 19208 25100
rect 19168 24818 19196 25094
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 19260 24138 19288 25706
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19352 25158 19380 25230
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19248 24132 19300 24138
rect 19248 24074 19300 24080
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19352 22098 19380 22918
rect 19076 22066 19196 22094
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 18892 16918 19012 16946
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18708 15502 18736 16390
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18800 15026 18828 15302
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18800 14618 18828 14962
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 18708 12850 18736 13670
rect 18788 13524 18840 13530
rect 18788 13466 18840 13472
rect 18800 12986 18828 13466
rect 18788 12980 18840 12986
rect 18788 12922 18840 12928
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18602 12336 18658 12345
rect 18602 12271 18658 12280
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18708 12050 18736 12786
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18800 12170 18828 12718
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18524 12022 18736 12050
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18144 10464 18196 10470
rect 18144 10406 18196 10412
rect 17512 9646 17724 9674
rect 17512 8498 17540 9646
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17880 9382 17908 9522
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17604 6662 17632 7482
rect 17776 6792 17828 6798
rect 17776 6734 17828 6740
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17604 5370 17632 6598
rect 17788 5710 17816 6734
rect 17880 5778 17908 9318
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17972 7818 18000 8434
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 17960 7812 18012 7818
rect 17960 7754 18012 7760
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17604 5137 17632 5306
rect 17696 5166 17724 5578
rect 17788 5234 17816 5646
rect 18064 5386 18092 7890
rect 18156 7546 18184 10406
rect 18524 9382 18552 12022
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 11354 18736 11494
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18144 7336 18196 7342
rect 18142 7304 18144 7313
rect 18196 7304 18198 7313
rect 18142 7239 18198 7248
rect 18156 5642 18184 7239
rect 18248 6798 18276 8230
rect 18340 8090 18368 8366
rect 18328 8084 18380 8090
rect 18328 8026 18380 8032
rect 18524 7546 18552 9318
rect 18708 9110 18736 9522
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18616 8294 18644 8434
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18604 7812 18656 7818
rect 18708 7800 18736 9046
rect 18892 8514 18920 16918
rect 19076 13394 19104 21830
rect 19064 13388 19116 13394
rect 19064 13330 19116 13336
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 18984 12918 19012 13126
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 18984 12764 19012 12854
rect 18984 12736 19104 12764
rect 19076 12238 19104 12736
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19076 12102 19104 12174
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11354 19104 12038
rect 19064 11348 19116 11354
rect 19064 11290 19116 11296
rect 19168 9058 19196 22066
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 19246 20496 19302 20505
rect 19246 20431 19248 20440
rect 19300 20431 19302 20440
rect 19248 20402 19300 20408
rect 19352 19786 19380 20878
rect 19444 20466 19472 25842
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19892 24676 19944 24682
rect 19892 24618 19944 24624
rect 19904 24206 19932 24618
rect 19892 24200 19944 24206
rect 19892 24142 19944 24148
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 19904 19854 19932 20198
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19260 18358 19288 18702
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19248 18352 19300 18358
rect 19248 18294 19300 18300
rect 19260 15570 19288 18294
rect 19340 18284 19392 18290
rect 19340 18226 19392 18232
rect 19352 16182 19380 18226
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19340 16176 19392 16182
rect 19340 16118 19392 16124
rect 19444 16046 19472 16390
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19892 16176 19944 16182
rect 19892 16118 19944 16124
rect 19904 16046 19932 16118
rect 19432 16040 19484 16046
rect 19432 15982 19484 15988
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19352 14074 19380 14350
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 19260 12434 19288 12786
rect 19260 12406 19380 12434
rect 19246 12336 19302 12345
rect 19246 12271 19302 12280
rect 19260 11762 19288 12271
rect 19352 12238 19380 12406
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19260 10470 19288 11698
rect 19444 11014 19472 15982
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19628 14414 19656 14554
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19996 9722 20024 56306
rect 20352 55616 20404 55622
rect 20350 55584 20352 55593
rect 20404 55584 20406 55593
rect 20350 55519 20406 55528
rect 20168 41608 20220 41614
rect 20168 41550 20220 41556
rect 20076 40520 20128 40526
rect 20180 40508 20208 41550
rect 20260 41472 20312 41478
rect 20260 41414 20312 41420
rect 20272 40594 20300 41414
rect 20444 40996 20496 41002
rect 20444 40938 20496 40944
rect 20260 40588 20312 40594
rect 20260 40530 20312 40536
rect 20128 40480 20208 40508
rect 20076 40462 20128 40468
rect 20088 39914 20116 40462
rect 20272 40440 20300 40530
rect 20456 40458 20484 40938
rect 20180 40412 20300 40440
rect 20444 40452 20496 40458
rect 20076 39908 20128 39914
rect 20076 39850 20128 39856
rect 20076 39296 20128 39302
rect 20180 39284 20208 40412
rect 20444 40394 20496 40400
rect 20352 40384 20404 40390
rect 20352 40326 20404 40332
rect 20364 39370 20392 40326
rect 20260 39364 20312 39370
rect 20260 39306 20312 39312
rect 20352 39364 20404 39370
rect 20352 39306 20404 39312
rect 20128 39256 20208 39284
rect 20076 39238 20128 39244
rect 20088 37942 20116 39238
rect 20076 37936 20128 37942
rect 20076 37878 20128 37884
rect 20088 36582 20116 37878
rect 20168 37868 20220 37874
rect 20168 37810 20220 37816
rect 20180 37466 20208 37810
rect 20168 37460 20220 37466
rect 20168 37402 20220 37408
rect 20076 36576 20128 36582
rect 20076 36518 20128 36524
rect 20168 34740 20220 34746
rect 20168 34682 20220 34688
rect 20076 34604 20128 34610
rect 20076 34546 20128 34552
rect 20088 34202 20116 34546
rect 20076 34196 20128 34202
rect 20076 34138 20128 34144
rect 20180 31754 20208 34682
rect 20272 34610 20300 39306
rect 20456 37942 20484 40394
rect 20444 37936 20496 37942
rect 20444 37878 20496 37884
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 20456 34542 20484 37878
rect 20444 34536 20496 34542
rect 20444 34478 20496 34484
rect 20088 31726 20208 31754
rect 20088 29492 20116 31726
rect 20260 30932 20312 30938
rect 20260 30874 20312 30880
rect 20088 29464 20208 29492
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 20088 28082 20116 29106
rect 20076 28076 20128 28082
rect 20076 28018 20128 28024
rect 20076 27940 20128 27946
rect 20076 27882 20128 27888
rect 20088 24614 20116 27882
rect 20180 27418 20208 29464
rect 20272 27606 20300 30874
rect 20444 30728 20496 30734
rect 20444 30670 20496 30676
rect 20456 30258 20484 30670
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20444 30252 20496 30258
rect 20444 30194 20496 30200
rect 20364 29850 20392 30194
rect 20352 29844 20404 29850
rect 20352 29786 20404 29792
rect 20352 29572 20404 29578
rect 20352 29514 20404 29520
rect 20364 29186 20392 29514
rect 20456 29306 20484 30194
rect 20444 29300 20496 29306
rect 20444 29242 20496 29248
rect 20364 29158 20484 29186
rect 20352 29028 20404 29034
rect 20352 28970 20404 28976
rect 20260 27600 20312 27606
rect 20260 27542 20312 27548
rect 20180 27390 20300 27418
rect 20168 26920 20220 26926
rect 20168 26862 20220 26868
rect 20180 25226 20208 26862
rect 20168 25220 20220 25226
rect 20168 25162 20220 25168
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20076 23044 20128 23050
rect 20076 22986 20128 22992
rect 20088 22506 20116 22986
rect 20180 22778 20208 25162
rect 20272 23322 20300 27390
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 20168 22772 20220 22778
rect 20168 22714 20220 22720
rect 20076 22500 20128 22506
rect 20076 22442 20128 22448
rect 20260 21888 20312 21894
rect 20260 21830 20312 21836
rect 20168 20868 20220 20874
rect 20168 20810 20220 20816
rect 20180 20398 20208 20810
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 20088 19446 20116 20198
rect 20180 19854 20208 20334
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 20076 16108 20128 16114
rect 20180 16096 20208 19790
rect 20128 16068 20208 16096
rect 20076 16050 20128 16056
rect 20088 15026 20116 16050
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20168 14952 20220 14958
rect 20168 14894 20220 14900
rect 20180 14414 20208 14894
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20076 13728 20128 13734
rect 20076 13670 20128 13676
rect 20088 12850 20116 13670
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 19168 9030 19288 9058
rect 18972 8968 19024 8974
rect 18972 8910 19024 8916
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 18656 7772 18736 7800
rect 18800 8486 18920 8514
rect 18604 7754 18656 7760
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18328 6656 18380 6662
rect 18328 6598 18380 6604
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 17972 5358 18092 5386
rect 18248 5370 18276 5646
rect 18236 5364 18288 5370
rect 17776 5228 17828 5234
rect 17776 5170 17828 5176
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17684 5160 17736 5166
rect 17590 5128 17646 5137
rect 17684 5102 17736 5108
rect 17590 5063 17646 5072
rect 17880 5030 17908 5170
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17868 5024 17920 5030
rect 17868 4966 17920 4972
rect 17500 3596 17552 3602
rect 17500 3538 17552 3544
rect 17408 2644 17460 2650
rect 17408 2586 17460 2592
rect 17512 800 17540 3538
rect 17604 800 17632 4966
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17682 4176 17738 4185
rect 17682 4111 17738 4120
rect 17696 3194 17724 4111
rect 17774 3768 17830 3777
rect 17774 3703 17776 3712
rect 17828 3703 17830 3712
rect 17776 3674 17828 3680
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17788 3058 17816 3334
rect 17880 3126 17908 4422
rect 17972 3670 18000 5358
rect 18236 5306 18288 5312
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 17776 3052 17828 3058
rect 17776 2994 17828 3000
rect 17788 800 17816 2994
rect 18064 2774 18092 4490
rect 18142 4040 18198 4049
rect 18142 3975 18198 3984
rect 18156 3194 18184 3975
rect 18340 3534 18368 6598
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18512 6180 18564 6186
rect 18512 6122 18564 6128
rect 18524 5574 18552 6122
rect 18616 5914 18644 6190
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18708 5710 18736 6054
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18512 5568 18564 5574
rect 18512 5510 18564 5516
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18064 2746 18184 2774
rect 18050 2680 18106 2689
rect 18050 2615 18106 2624
rect 18064 2582 18092 2615
rect 18052 2576 18104 2582
rect 18052 2518 18104 2524
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17880 800 17908 2382
rect 18052 1896 18104 1902
rect 18052 1838 18104 1844
rect 18064 800 18092 1838
rect 18156 800 18184 2746
rect 18340 800 18368 3470
rect 18432 800 18460 3946
rect 18524 3942 18552 5510
rect 18696 4752 18748 4758
rect 18696 4694 18748 4700
rect 18602 4040 18658 4049
rect 18602 3975 18658 3984
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18616 3738 18644 3975
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18524 2310 18552 2994
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18524 1766 18552 2246
rect 18512 1760 18564 1766
rect 18512 1702 18564 1708
rect 18616 800 18644 3062
rect 18708 800 18736 4694
rect 18800 3738 18828 8486
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18892 7342 18920 8366
rect 18984 8362 19012 8910
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 19076 7886 19104 8910
rect 19156 8900 19208 8906
rect 19156 8842 19208 8848
rect 19168 8634 19196 8842
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19168 8294 19196 8434
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 19076 6390 19104 7822
rect 19260 7562 19288 9030
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 19444 7750 19472 8434
rect 20088 8430 20116 12786
rect 20168 12368 20220 12374
rect 20168 12310 20220 12316
rect 20180 12170 20208 12310
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20180 11354 20208 12106
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20076 8424 20128 8430
rect 20076 8366 20128 8372
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19168 7534 19288 7562
rect 19064 6384 19116 6390
rect 19064 6326 19116 6332
rect 19076 5778 19104 6326
rect 19064 5772 19116 5778
rect 19064 5714 19116 5720
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18786 3224 18842 3233
rect 18786 3159 18842 3168
rect 18800 3126 18828 3159
rect 18788 3120 18840 3126
rect 18788 3062 18840 3068
rect 18892 2854 18920 3878
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18880 1760 18932 1766
rect 18880 1702 18932 1708
rect 18892 800 18920 1702
rect 18984 800 19012 4626
rect 19076 4146 19104 5714
rect 19064 4140 19116 4146
rect 19064 4082 19116 4088
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 19076 1442 19104 3062
rect 19168 2582 19196 7534
rect 19444 7410 19472 7686
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 19260 6882 19288 7142
rect 19444 6934 19472 7346
rect 20180 7206 20208 7346
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 19432 6928 19484 6934
rect 19260 6854 19380 6882
rect 19432 6870 19484 6876
rect 20180 6866 20208 7142
rect 19352 6390 19380 6854
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19524 6384 19576 6390
rect 19524 6326 19576 6332
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19352 5098 19380 5578
rect 19340 5092 19392 5098
rect 19340 5034 19392 5040
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19156 2576 19208 2582
rect 19156 2518 19208 2524
rect 19076 1414 19196 1442
rect 19168 800 19196 1414
rect 19260 800 19288 4558
rect 19352 1358 19380 4558
rect 19444 4264 19472 5850
rect 19536 5556 19564 6326
rect 19505 5528 19564 5556
rect 19505 5302 19533 5528
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19505 5296 19576 5302
rect 19505 5256 19524 5296
rect 19524 5238 19576 5244
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19444 4236 19564 4264
rect 19536 4146 19564 4236
rect 19524 4140 19576 4146
rect 19524 4082 19576 4088
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 19444 3398 19472 3878
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19430 3224 19486 3233
rect 19574 3227 19882 3236
rect 19430 3159 19432 3168
rect 19484 3159 19486 3168
rect 19432 3130 19484 3136
rect 19522 3088 19578 3097
rect 19996 3058 20024 6598
rect 20076 6112 20128 6118
rect 20076 6054 20128 6060
rect 20088 5166 20116 6054
rect 20076 5160 20128 5166
rect 20076 5102 20128 5108
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19522 3023 19578 3032
rect 19984 3052 20036 3058
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19340 1352 19392 1358
rect 19340 1294 19392 1300
rect 19444 1290 19472 2858
rect 19536 2446 19564 3023
rect 19984 2994 20036 3000
rect 19524 2440 19576 2446
rect 19524 2382 19576 2388
rect 19536 2292 19564 2382
rect 19505 2264 19564 2292
rect 19505 2088 19533 2264
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19505 2060 19564 2088
rect 19432 1284 19484 1290
rect 19432 1226 19484 1232
rect 19536 1170 19564 2060
rect 19996 1442 20024 2994
rect 19444 1142 19564 1170
rect 19720 1414 20024 1442
rect 20088 1442 20116 4966
rect 20180 3126 20208 6666
rect 20272 3505 20300 21830
rect 20364 19922 20392 28970
rect 20456 28762 20484 29158
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20456 26926 20484 28698
rect 20444 26920 20496 26926
rect 20444 26862 20496 26868
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 20456 25974 20484 26726
rect 20444 25968 20496 25974
rect 20444 25910 20496 25916
rect 20444 25152 20496 25158
rect 20444 25094 20496 25100
rect 20456 24682 20484 25094
rect 20444 24676 20496 24682
rect 20444 24618 20496 24624
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20456 21418 20484 21490
rect 20444 21412 20496 21418
rect 20444 21354 20496 21360
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20456 20330 20484 20402
rect 20444 20324 20496 20330
rect 20444 20266 20496 20272
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20364 17202 20392 19654
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20364 14414 20392 14758
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20364 3942 20392 7686
rect 20456 7410 20484 18022
rect 20548 13705 20576 56306
rect 21100 55826 21128 56306
rect 21088 55820 21140 55826
rect 21088 55762 21140 55768
rect 20720 41472 20772 41478
rect 20720 41414 20772 41420
rect 20732 41138 20760 41414
rect 20720 41132 20772 41138
rect 20720 41074 20772 41080
rect 20628 40996 20680 41002
rect 20628 40938 20680 40944
rect 20640 40730 20668 40938
rect 20628 40724 20680 40730
rect 20628 40666 20680 40672
rect 20628 40520 20680 40526
rect 20628 40462 20680 40468
rect 20640 39438 20668 40462
rect 21456 40180 21508 40186
rect 21456 40122 21508 40128
rect 21468 40050 21496 40122
rect 21456 40044 21508 40050
rect 21456 39986 21508 39992
rect 20628 39432 20680 39438
rect 20628 39374 20680 39380
rect 20640 38418 20668 39374
rect 20628 38412 20680 38418
rect 20628 38354 20680 38360
rect 21272 37732 21324 37738
rect 21272 37674 21324 37680
rect 20996 37664 21048 37670
rect 20996 37606 21048 37612
rect 21008 37262 21036 37606
rect 20996 37256 21048 37262
rect 20996 37198 21048 37204
rect 20812 35148 20864 35154
rect 20812 35090 20864 35096
rect 20628 32020 20680 32026
rect 20628 31962 20680 31968
rect 20640 29322 20668 31962
rect 20824 31278 20852 35090
rect 21088 35012 21140 35018
rect 21088 34954 21140 34960
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20824 29782 20852 31214
rect 20904 31136 20956 31142
rect 20904 31078 20956 31084
rect 20916 30258 20944 31078
rect 20904 30252 20956 30258
rect 20904 30194 20956 30200
rect 20812 29776 20864 29782
rect 20812 29718 20864 29724
rect 20640 29294 20760 29322
rect 20732 28370 20760 29294
rect 20640 28342 20760 28370
rect 20996 28416 21048 28422
rect 20996 28358 21048 28364
rect 20640 23798 20668 28342
rect 20812 27124 20864 27130
rect 20812 27066 20864 27072
rect 20824 26994 20852 27066
rect 20812 26988 20864 26994
rect 20812 26930 20864 26936
rect 20824 26314 20852 26930
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 20812 26308 20864 26314
rect 20812 26250 20864 26256
rect 20628 23792 20680 23798
rect 20628 23734 20680 23740
rect 20628 22500 20680 22506
rect 20628 22442 20680 22448
rect 20640 20466 20668 22442
rect 20824 22234 20852 26250
rect 20916 25906 20944 26862
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 20904 24744 20956 24750
rect 20904 24686 20956 24692
rect 20916 24342 20944 24686
rect 20904 24336 20956 24342
rect 20904 24278 20956 24284
rect 20904 24064 20956 24070
rect 20904 24006 20956 24012
rect 20916 22642 20944 24006
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 21008 22386 21036 28358
rect 21100 22438 21128 34954
rect 21180 32360 21232 32366
rect 21180 32302 21232 32308
rect 21192 29646 21220 32302
rect 21180 29640 21232 29646
rect 21180 29582 21232 29588
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 20916 22358 21036 22386
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 20812 22228 20864 22234
rect 20812 22170 20864 22176
rect 20812 22092 20864 22098
rect 20812 22034 20864 22040
rect 20720 21956 20772 21962
rect 20720 21898 20772 21904
rect 20732 21690 20760 21898
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20824 20534 20852 22034
rect 20812 20528 20864 20534
rect 20812 20470 20864 20476
rect 20916 20466 20944 22358
rect 20996 22228 21048 22234
rect 20996 22170 21048 22176
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20720 19780 20772 19786
rect 20720 19722 20772 19728
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20640 15366 20668 15982
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20640 13938 20668 15302
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 20534 13696 20590 13705
rect 20534 13631 20590 13640
rect 20732 13138 20760 19722
rect 20904 18080 20956 18086
rect 20904 18022 20956 18028
rect 20916 17746 20944 18022
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20810 17640 20866 17649
rect 20810 17575 20812 17584
rect 20864 17575 20866 17584
rect 20812 17546 20864 17552
rect 20916 17320 20944 17682
rect 20824 17292 20944 17320
rect 20824 14822 20852 17292
rect 21008 17218 21036 22170
rect 21192 19854 21220 26726
rect 21284 24698 21312 37674
rect 21364 36576 21416 36582
rect 21364 36518 21416 36524
rect 21376 27962 21404 36518
rect 21468 31754 21496 39986
rect 21548 34944 21600 34950
rect 21548 34886 21600 34892
rect 21560 34678 21588 34886
rect 21548 34672 21600 34678
rect 21548 34614 21600 34620
rect 21548 34536 21600 34542
rect 21548 34478 21600 34484
rect 21560 33998 21588 34478
rect 21548 33992 21600 33998
rect 21548 33934 21600 33940
rect 21468 31726 21588 31754
rect 21456 30116 21508 30122
rect 21456 30058 21508 30064
rect 21468 29646 21496 30058
rect 21560 29850 21588 31726
rect 21652 30326 21680 56306
rect 22572 55622 22600 56306
rect 22560 55616 22612 55622
rect 22558 55584 22560 55593
rect 22612 55584 22614 55593
rect 22558 55519 22614 55528
rect 23480 41472 23532 41478
rect 23480 41414 23532 41420
rect 23492 41386 23704 41414
rect 23388 41200 23440 41206
rect 23388 41142 23440 41148
rect 22192 41132 22244 41138
rect 22192 41074 22244 41080
rect 23020 41132 23072 41138
rect 23020 41074 23072 41080
rect 23112 41132 23164 41138
rect 23112 41074 23164 41080
rect 22100 40656 22152 40662
rect 22100 40598 22152 40604
rect 21824 40452 21876 40458
rect 21824 40394 21876 40400
rect 21836 40186 21864 40394
rect 22112 40186 22140 40598
rect 22204 40390 22232 41074
rect 22928 41064 22980 41070
rect 22928 41006 22980 41012
rect 22284 40928 22336 40934
rect 22284 40870 22336 40876
rect 22192 40384 22244 40390
rect 22192 40326 22244 40332
rect 21824 40180 21876 40186
rect 21824 40122 21876 40128
rect 22100 40180 22152 40186
rect 22100 40122 22152 40128
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 21928 36854 21956 37198
rect 21916 36848 21968 36854
rect 21916 36790 21968 36796
rect 21928 34610 21956 36790
rect 22112 35222 22140 40122
rect 22296 40050 22324 40870
rect 22940 40526 22968 41006
rect 23032 40730 23060 41074
rect 23020 40724 23072 40730
rect 23020 40666 23072 40672
rect 23124 40662 23152 41074
rect 23296 40996 23348 41002
rect 23296 40938 23348 40944
rect 23112 40656 23164 40662
rect 23112 40598 23164 40604
rect 23308 40526 23336 40938
rect 22928 40520 22980 40526
rect 22928 40462 22980 40468
rect 23296 40520 23348 40526
rect 23296 40462 23348 40468
rect 22652 40384 22704 40390
rect 22652 40326 22704 40332
rect 22284 40044 22336 40050
rect 22284 39986 22336 39992
rect 22192 39908 22244 39914
rect 22192 39850 22244 39856
rect 22100 35216 22152 35222
rect 22100 35158 22152 35164
rect 22204 35086 22232 39850
rect 22284 37664 22336 37670
rect 22284 37606 22336 37612
rect 22296 37262 22324 37606
rect 22284 37256 22336 37262
rect 22284 37198 22336 37204
rect 22296 36786 22324 37198
rect 22664 36786 22692 40326
rect 22940 40050 22968 40462
rect 23020 40452 23072 40458
rect 23020 40394 23072 40400
rect 23032 40186 23060 40394
rect 23400 40186 23428 41142
rect 23676 41138 23704 41386
rect 23664 41132 23716 41138
rect 23664 41074 23716 41080
rect 23480 40928 23532 40934
rect 23480 40870 23532 40876
rect 23020 40180 23072 40186
rect 23388 40180 23440 40186
rect 23020 40122 23072 40128
rect 23308 40140 23388 40168
rect 22928 40044 22980 40050
rect 22928 39986 22980 39992
rect 23204 39908 23256 39914
rect 23204 39850 23256 39856
rect 23112 37664 23164 37670
rect 23112 37606 23164 37612
rect 23124 37194 23152 37606
rect 23216 37262 23244 39850
rect 23204 37256 23256 37262
rect 23204 37198 23256 37204
rect 23112 37188 23164 37194
rect 23112 37130 23164 37136
rect 22744 37120 22796 37126
rect 22744 37062 22796 37068
rect 22284 36780 22336 36786
rect 22284 36722 22336 36728
rect 22468 36780 22520 36786
rect 22468 36722 22520 36728
rect 22652 36780 22704 36786
rect 22652 36722 22704 36728
rect 22296 35850 22324 36722
rect 22480 36582 22508 36722
rect 22468 36576 22520 36582
rect 22468 36518 22520 36524
rect 22652 36576 22704 36582
rect 22652 36518 22704 36524
rect 22664 36038 22692 36518
rect 22652 36032 22704 36038
rect 22756 36009 22784 37062
rect 23124 36582 23152 37130
rect 23112 36576 23164 36582
rect 23112 36518 23164 36524
rect 23020 36032 23072 36038
rect 22652 35974 22704 35980
rect 22742 36000 22798 36009
rect 22296 35822 22416 35850
rect 22388 35698 22416 35822
rect 22664 35766 22692 35974
rect 23020 35974 23072 35980
rect 22742 35935 22798 35944
rect 22652 35760 22704 35766
rect 22652 35702 22704 35708
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 22388 35494 22416 35634
rect 22376 35488 22428 35494
rect 22376 35430 22428 35436
rect 22100 35080 22152 35086
rect 22100 35022 22152 35028
rect 22192 35080 22244 35086
rect 22192 35022 22244 35028
rect 21916 34604 21968 34610
rect 21916 34546 21968 34552
rect 21928 34490 21956 34546
rect 21928 34462 22048 34490
rect 22020 33998 22048 34462
rect 22112 34202 22140 35022
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 22100 33856 22152 33862
rect 22100 33798 22152 33804
rect 22112 31822 22140 33798
rect 22204 32366 22232 35022
rect 22192 32360 22244 32366
rect 22192 32302 22244 32308
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 22008 31136 22060 31142
rect 22008 31078 22060 31084
rect 22020 30734 22048 31078
rect 21732 30728 21784 30734
rect 21732 30670 21784 30676
rect 22008 30728 22060 30734
rect 22008 30670 22060 30676
rect 21640 30320 21692 30326
rect 21640 30262 21692 30268
rect 21640 30184 21692 30190
rect 21640 30126 21692 30132
rect 21548 29844 21600 29850
rect 21548 29786 21600 29792
rect 21456 29640 21508 29646
rect 21456 29582 21508 29588
rect 21468 29306 21496 29582
rect 21456 29300 21508 29306
rect 21456 29242 21508 29248
rect 21456 28552 21508 28558
rect 21456 28494 21508 28500
rect 21468 28082 21496 28494
rect 21456 28076 21508 28082
rect 21456 28018 21508 28024
rect 21376 27934 21496 27962
rect 21284 24670 21404 24698
rect 21272 24132 21324 24138
rect 21272 24074 21324 24080
rect 21284 23798 21312 24074
rect 21272 23792 21324 23798
rect 21272 23734 21324 23740
rect 21376 23322 21404 24670
rect 21468 24206 21496 27934
rect 21560 24970 21588 29786
rect 21652 29578 21680 30126
rect 21640 29572 21692 29578
rect 21640 29514 21692 29520
rect 21652 29170 21680 29514
rect 21640 29164 21692 29170
rect 21640 29106 21692 29112
rect 21652 28966 21680 29106
rect 21640 28960 21692 28966
rect 21640 28902 21692 28908
rect 21652 28558 21680 28902
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 21744 27402 21772 30670
rect 22112 30666 22140 31758
rect 22204 31226 22232 32302
rect 22284 31952 22336 31958
rect 22284 31894 22336 31900
rect 22296 31346 22324 31894
rect 22388 31754 22416 35430
rect 22664 31754 22692 35702
rect 23032 35698 23060 35974
rect 23020 35692 23072 35698
rect 23020 35634 23072 35640
rect 23112 35692 23164 35698
rect 23112 35634 23164 35640
rect 23020 35488 23072 35494
rect 23020 35430 23072 35436
rect 22836 34400 22888 34406
rect 22756 34348 22836 34354
rect 22756 34342 22888 34348
rect 22756 34326 22876 34342
rect 22756 33930 22784 34326
rect 22744 33924 22796 33930
rect 22744 33866 22796 33872
rect 22388 31726 22600 31754
rect 22468 31680 22520 31686
rect 22468 31622 22520 31628
rect 22572 31634 22600 31726
rect 22652 31748 22704 31754
rect 22652 31690 22704 31696
rect 22480 31346 22508 31622
rect 22572 31606 22692 31634
rect 22282 31340 22334 31346
rect 22282 31282 22334 31288
rect 22468 31340 22520 31346
rect 22468 31282 22520 31288
rect 22560 31272 22612 31278
rect 22204 31220 22560 31226
rect 22204 31214 22612 31220
rect 22204 31198 22600 31214
rect 22100 30660 22152 30666
rect 22100 30602 22152 30608
rect 22192 30592 22244 30598
rect 22192 30534 22244 30540
rect 22100 30320 22152 30326
rect 22100 30262 22152 30268
rect 21824 30252 21876 30258
rect 21824 30194 21876 30200
rect 21836 28558 21864 30194
rect 22112 29458 22140 30262
rect 22204 29646 22232 30534
rect 22284 30252 22336 30258
rect 22284 30194 22336 30200
rect 22296 29646 22324 30194
rect 22376 30048 22428 30054
rect 22376 29990 22428 29996
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 22284 29640 22336 29646
rect 22284 29582 22336 29588
rect 22112 29430 22232 29458
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 21732 27396 21784 27402
rect 21732 27338 21784 27344
rect 21744 27062 21772 27338
rect 21732 27056 21784 27062
rect 21732 26998 21784 27004
rect 21640 25900 21692 25906
rect 21640 25842 21692 25848
rect 21652 25158 21680 25842
rect 21744 25294 21772 26998
rect 21916 26852 21968 26858
rect 21916 26794 21968 26800
rect 21824 26376 21876 26382
rect 21824 26318 21876 26324
rect 21836 26042 21864 26318
rect 21824 26036 21876 26042
rect 21824 25978 21876 25984
rect 21836 25906 21864 25978
rect 21824 25900 21876 25906
rect 21824 25842 21876 25848
rect 21732 25288 21784 25294
rect 21732 25230 21784 25236
rect 21640 25152 21692 25158
rect 21640 25094 21692 25100
rect 21560 24942 21680 24970
rect 21652 24682 21680 24942
rect 21744 24818 21772 25230
rect 21732 24812 21784 24818
rect 21732 24754 21784 24760
rect 21640 24676 21692 24682
rect 21640 24618 21692 24624
rect 21548 24608 21600 24614
rect 21548 24550 21600 24556
rect 21560 24274 21588 24550
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21468 23730 21496 24006
rect 21732 23792 21784 23798
rect 21732 23734 21784 23740
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 21376 22506 21404 23258
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 21468 21078 21496 23666
rect 21640 22432 21692 22438
rect 21640 22374 21692 22380
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21456 21072 21508 21078
rect 21456 21014 21508 21020
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21192 19514 21220 19790
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21284 18222 21312 20810
rect 21456 19304 21508 19310
rect 21456 19246 21508 19252
rect 21272 18216 21324 18222
rect 21272 18158 21324 18164
rect 21364 17672 21416 17678
rect 21364 17614 21416 17620
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 20916 17190 21036 17218
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20640 13110 20760 13138
rect 20640 12918 20668 13110
rect 20824 13002 20852 14554
rect 20732 12974 20852 13002
rect 20628 12912 20680 12918
rect 20628 12854 20680 12860
rect 20732 9654 20760 12974
rect 20812 12912 20864 12918
rect 20812 12854 20864 12860
rect 20824 11898 20852 12854
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20916 11064 20944 17190
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 21008 16114 21036 16594
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21008 15570 21036 16050
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14618 21036 14758
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 21008 12306 21036 14554
rect 21100 12986 21128 17478
rect 21376 16998 21404 17614
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21180 16720 21232 16726
rect 21180 16662 21232 16668
rect 21192 16046 21220 16662
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21192 15434 21220 15982
rect 21468 15910 21496 19246
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21180 15428 21232 15434
rect 21180 15370 21232 15376
rect 21284 14074 21312 15438
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21376 13870 21404 14350
rect 21364 13864 21416 13870
rect 21364 13806 21416 13812
rect 21376 13190 21404 13806
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21192 12730 21220 12786
rect 21100 12702 21220 12730
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 21100 11150 21128 12702
rect 21376 11286 21404 13126
rect 21468 12850 21496 15846
rect 21560 15706 21588 21490
rect 21548 15700 21600 15706
rect 21548 15642 21600 15648
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21652 12782 21680 22374
rect 21744 20806 21772 23734
rect 21836 21622 21864 25842
rect 21928 24342 21956 26794
rect 22008 26784 22060 26790
rect 22008 26726 22060 26732
rect 22020 26382 22048 26726
rect 21987 26376 22048 26382
rect 22039 26336 22048 26376
rect 22100 26376 22152 26382
rect 21987 26318 22039 26324
rect 22100 26318 22152 26324
rect 22112 26246 22140 26318
rect 22100 26240 22152 26246
rect 22100 26182 22152 26188
rect 22204 26194 22232 29430
rect 22296 28150 22324 29582
rect 22284 28144 22336 28150
rect 22284 28086 22336 28092
rect 22112 25906 22140 26182
rect 22204 26166 22324 26194
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 22112 24206 22140 24754
rect 22192 24608 22244 24614
rect 22192 24550 22244 24556
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 21916 24064 21968 24070
rect 21916 24006 21968 24012
rect 21928 22030 21956 24006
rect 22204 22642 22232 24550
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22006 22264 22062 22273
rect 22006 22199 22008 22208
rect 22060 22199 22062 22208
rect 22008 22170 22060 22176
rect 21916 22024 21968 22030
rect 21916 21966 21968 21972
rect 21824 21616 21876 21622
rect 21824 21558 21876 21564
rect 21732 20800 21784 20806
rect 21732 20742 21784 20748
rect 21916 20392 21968 20398
rect 21916 20334 21968 20340
rect 21928 19446 21956 20334
rect 21916 19440 21968 19446
rect 21916 19382 21968 19388
rect 21824 19168 21876 19174
rect 21824 19110 21876 19116
rect 21836 17746 21864 19110
rect 21928 17882 21956 19382
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21824 17740 21876 17746
rect 21824 17682 21876 17688
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21732 14340 21784 14346
rect 21732 14282 21784 14288
rect 21744 13462 21772 14282
rect 21732 13456 21784 13462
rect 21732 13398 21784 13404
rect 21836 13410 21864 16934
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21928 14346 21956 15302
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 22020 13530 22048 22170
rect 22100 21956 22152 21962
rect 22100 21898 22152 21904
rect 22112 21010 22140 21898
rect 22192 21344 22244 21350
rect 22192 21286 22244 21292
rect 22100 21004 22152 21010
rect 22100 20946 22152 20952
rect 22112 20466 22140 20946
rect 22204 20874 22232 21286
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22112 18834 22140 19994
rect 22204 19854 22232 20810
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22204 18834 22232 19314
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22192 18828 22244 18834
rect 22192 18770 22244 18776
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 22112 15978 22140 16390
rect 22100 15972 22152 15978
rect 22100 15914 22152 15920
rect 22112 15502 22140 15914
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22204 15434 22232 15846
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22112 14074 22140 15030
rect 22204 14958 22232 15370
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 22204 14822 22232 14894
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22204 14006 22232 14758
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 22008 13524 22060 13530
rect 22008 13466 22060 13472
rect 21836 13382 22140 13410
rect 21640 12776 21692 12782
rect 21640 12718 21692 12724
rect 21916 12640 21968 12646
rect 21916 12582 21968 12588
rect 21456 12300 21508 12306
rect 21456 12242 21508 12248
rect 21468 11830 21496 12242
rect 21928 12238 21956 12582
rect 22008 12368 22060 12374
rect 22008 12310 22060 12316
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21456 11824 21508 11830
rect 21456 11766 21508 11772
rect 22020 11762 22048 12310
rect 22112 12238 22140 13382
rect 22192 13252 22244 13258
rect 22192 13194 22244 13200
rect 22204 12782 22232 13194
rect 22192 12776 22244 12782
rect 22192 12718 22244 12724
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22204 12170 22232 12718
rect 22192 12164 22244 12170
rect 22192 12106 22244 12112
rect 22204 11762 22232 12106
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21652 11354 21680 11630
rect 21916 11552 21968 11558
rect 21916 11494 21968 11500
rect 21640 11348 21692 11354
rect 21640 11290 21692 11296
rect 21364 11280 21416 11286
rect 21364 11222 21416 11228
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 20996 11076 21048 11082
rect 20916 11036 20996 11064
rect 20996 11018 21048 11024
rect 21008 10470 21036 11018
rect 21376 10606 21404 11222
rect 21652 11218 21680 11290
rect 21640 11212 21692 11218
rect 21640 11154 21692 11160
rect 21928 11150 21956 11494
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20640 8566 20668 9114
rect 20732 8974 20760 9590
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 21180 8900 21232 8906
rect 21180 8842 21232 8848
rect 21192 8786 21220 8842
rect 21100 8758 21220 8786
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 21100 8430 21128 8758
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 20536 7812 20588 7818
rect 20536 7754 20588 7760
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20444 7268 20496 7274
rect 20444 7210 20496 7216
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20350 3768 20406 3777
rect 20350 3703 20406 3712
rect 20364 3670 20392 3703
rect 20352 3664 20404 3670
rect 20352 3606 20404 3612
rect 20258 3496 20314 3505
rect 20258 3431 20314 3440
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20350 3360 20406 3369
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 20272 3074 20300 3334
rect 20350 3295 20406 3304
rect 20364 3194 20392 3295
rect 20352 3188 20404 3194
rect 20352 3130 20404 3136
rect 20272 3046 20392 3074
rect 20260 2984 20312 2990
rect 20260 2926 20312 2932
rect 20166 2680 20222 2689
rect 20166 2615 20222 2624
rect 20180 2582 20208 2615
rect 20168 2576 20220 2582
rect 20168 2518 20220 2524
rect 20272 2378 20300 2926
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20272 1630 20300 2314
rect 20260 1624 20312 1630
rect 20260 1566 20312 1572
rect 20364 1562 20392 3046
rect 20456 2990 20484 7210
rect 20548 3233 20576 7754
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 20640 5914 20668 6258
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20628 4616 20680 4622
rect 20628 4558 20680 4564
rect 20534 3224 20590 3233
rect 20534 3159 20590 3168
rect 20536 3120 20588 3126
rect 20536 3062 20588 3068
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20444 2848 20496 2854
rect 20444 2790 20496 2796
rect 20352 1556 20404 1562
rect 20352 1498 20404 1504
rect 20260 1488 20312 1494
rect 20088 1414 20208 1442
rect 20456 1442 20484 2790
rect 20260 1430 20312 1436
rect 19444 800 19472 1142
rect 19524 944 19576 950
rect 19524 886 19576 892
rect 19536 800 19564 886
rect 19720 800 19748 1414
rect 19800 1352 19852 1358
rect 19800 1294 19852 1300
rect 19984 1352 20036 1358
rect 19984 1294 20036 1300
rect 19812 800 19840 1294
rect 19996 800 20024 1294
rect 20180 1170 20208 1414
rect 20088 1142 20208 1170
rect 20088 800 20116 1142
rect 20272 800 20300 1430
rect 20364 1414 20484 1442
rect 20364 800 20392 1414
rect 20548 800 20576 3062
rect 20640 800 20668 4558
rect 20732 3126 20760 6598
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20824 3534 20852 6054
rect 20996 5364 21048 5370
rect 20996 5306 21048 5312
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20720 3120 20772 3126
rect 20720 3062 20772 3068
rect 20824 800 20852 3470
rect 20916 800 20944 4966
rect 21008 4146 21036 5306
rect 21100 4826 21128 8366
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21192 7002 21220 7346
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 21284 7002 21312 7142
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20994 4040 21050 4049
rect 20994 3975 21050 3984
rect 21008 3126 21036 3975
rect 20996 3120 21048 3126
rect 20996 3062 21048 3068
rect 21100 2774 21128 4558
rect 21192 3126 21220 6054
rect 21376 3670 21404 9658
rect 21652 7750 21680 10406
rect 22192 9512 22244 9518
rect 22192 9454 22244 9460
rect 22204 9042 22232 9454
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 21836 8498 21864 8978
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21652 7410 21680 7686
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21916 7200 21968 7206
rect 21914 7168 21916 7177
rect 21968 7168 21970 7177
rect 21914 7103 21970 7112
rect 21640 6792 21692 6798
rect 21640 6734 21692 6740
rect 21652 6254 21680 6734
rect 22008 6452 22060 6458
rect 22008 6394 22060 6400
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 22020 6186 22048 6394
rect 22204 6390 22232 7414
rect 22192 6384 22244 6390
rect 22192 6326 22244 6332
rect 22204 6254 22232 6326
rect 22192 6248 22244 6254
rect 22192 6190 22244 6196
rect 22008 6180 22060 6186
rect 22008 6122 22060 6128
rect 22204 5710 22232 6190
rect 22192 5704 22244 5710
rect 22192 5646 22244 5652
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21456 3596 21508 3602
rect 21456 3538 21508 3544
rect 21180 3120 21232 3126
rect 21232 3080 21404 3108
rect 21180 3062 21232 3068
rect 21272 2848 21324 2854
rect 21272 2790 21324 2796
rect 21100 2746 21220 2774
rect 21088 1692 21140 1698
rect 21088 1634 21140 1640
rect 21100 800 21128 1634
rect 21192 800 21220 2746
rect 21284 2446 21312 2790
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 21376 800 21404 3080
rect 21468 800 21496 3538
rect 21560 2378 21588 3946
rect 21652 3534 21680 5510
rect 21732 5024 21784 5030
rect 21732 4966 21784 4972
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21548 2372 21600 2378
rect 21548 2314 21600 2320
rect 21560 1698 21588 2314
rect 21548 1692 21600 1698
rect 21548 1634 21600 1640
rect 21652 800 21680 3470
rect 21744 800 21772 4966
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 22192 4616 22244 4622
rect 22192 4558 22244 4564
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21836 1442 21864 2790
rect 21928 1578 21956 4558
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 22112 2258 22140 3062
rect 22204 2360 22232 4558
rect 22296 3194 22324 26166
rect 22388 22098 22416 29990
rect 22560 29028 22612 29034
rect 22560 28970 22612 28976
rect 22468 26988 22520 26994
rect 22468 26930 22520 26936
rect 22480 26586 22508 26930
rect 22468 26580 22520 26586
rect 22468 26522 22520 26528
rect 22468 26308 22520 26314
rect 22468 26250 22520 26256
rect 22480 25974 22508 26250
rect 22468 25968 22520 25974
rect 22468 25910 22520 25916
rect 22468 25696 22520 25702
rect 22468 25638 22520 25644
rect 22480 25226 22508 25638
rect 22468 25220 22520 25226
rect 22468 25162 22520 25168
rect 22572 25106 22600 28970
rect 22664 27946 22692 31606
rect 22756 30258 22784 33866
rect 22836 31748 22888 31754
rect 22836 31690 22888 31696
rect 22744 30252 22796 30258
rect 22744 30194 22796 30200
rect 22848 29034 22876 31690
rect 22928 31680 22980 31686
rect 22928 31622 22980 31628
rect 22940 30598 22968 31622
rect 22928 30592 22980 30598
rect 22928 30534 22980 30540
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 22836 29028 22888 29034
rect 22836 28970 22888 28976
rect 22652 27940 22704 27946
rect 22652 27882 22704 27888
rect 22480 25078 22600 25106
rect 22480 23322 22508 25078
rect 22558 24848 22614 24857
rect 22558 24783 22614 24792
rect 22572 24342 22600 24783
rect 22560 24336 22612 24342
rect 22560 24278 22612 24284
rect 22560 23588 22612 23594
rect 22560 23530 22612 23536
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 22572 23118 22600 23530
rect 22560 23112 22612 23118
rect 22560 23054 22612 23060
rect 22664 23050 22692 27882
rect 22836 25152 22888 25158
rect 22836 25094 22888 25100
rect 22848 24818 22876 25094
rect 22744 24812 22796 24818
rect 22744 24754 22796 24760
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22756 24138 22784 24754
rect 22744 24132 22796 24138
rect 22744 24074 22796 24080
rect 22756 23798 22784 24074
rect 22744 23792 22796 23798
rect 22744 23734 22796 23740
rect 22940 23712 22968 29446
rect 23032 24818 23060 35430
rect 23124 35086 23152 35634
rect 23112 35080 23164 35086
rect 23112 35022 23164 35028
rect 23308 33930 23336 40140
rect 23388 40122 23440 40128
rect 23388 40044 23440 40050
rect 23388 39986 23440 39992
rect 23400 38758 23428 39986
rect 23492 39370 23520 40870
rect 23572 40384 23624 40390
rect 23572 40326 23624 40332
rect 23584 40118 23612 40326
rect 23572 40112 23624 40118
rect 23572 40054 23624 40060
rect 23676 40050 23704 41074
rect 23756 40180 23808 40186
rect 23756 40122 23808 40128
rect 23664 40044 23716 40050
rect 23664 39986 23716 39992
rect 23768 39914 23796 40122
rect 23848 39976 23900 39982
rect 23848 39918 23900 39924
rect 23756 39908 23808 39914
rect 23756 39850 23808 39856
rect 23860 39438 23888 39918
rect 23848 39432 23900 39438
rect 23848 39374 23900 39380
rect 23480 39364 23532 39370
rect 23480 39306 23532 39312
rect 23388 38752 23440 38758
rect 23388 38694 23440 38700
rect 23400 38554 23428 38694
rect 23388 38548 23440 38554
rect 23388 38490 23440 38496
rect 23296 33924 23348 33930
rect 23296 33866 23348 33872
rect 23756 33924 23808 33930
rect 23756 33866 23808 33872
rect 23480 33584 23532 33590
rect 23480 33526 23532 33532
rect 23492 32910 23520 33526
rect 23768 33046 23796 33866
rect 23756 33040 23808 33046
rect 23756 32982 23808 32988
rect 23480 32904 23532 32910
rect 23480 32846 23532 32852
rect 23492 32298 23520 32846
rect 23664 32836 23716 32842
rect 23664 32778 23716 32784
rect 23572 32768 23624 32774
rect 23572 32710 23624 32716
rect 23480 32292 23532 32298
rect 23480 32234 23532 32240
rect 23584 31754 23612 32710
rect 23676 32570 23704 32778
rect 23664 32564 23716 32570
rect 23664 32506 23716 32512
rect 23584 31748 23716 31754
rect 23584 31726 23664 31748
rect 23664 31690 23716 31696
rect 23676 31346 23704 31690
rect 23664 31340 23716 31346
rect 23664 31282 23716 31288
rect 23676 31142 23704 31282
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 23676 30598 23704 31078
rect 23664 30592 23716 30598
rect 23664 30534 23716 30540
rect 23296 29844 23348 29850
rect 23296 29786 23348 29792
rect 23308 29238 23336 29786
rect 23296 29232 23348 29238
rect 23296 29174 23348 29180
rect 23388 29232 23440 29238
rect 23388 29174 23440 29180
rect 23400 28422 23428 29174
rect 23572 28484 23624 28490
rect 23572 28426 23624 28432
rect 23388 28416 23440 28422
rect 23388 28358 23440 28364
rect 23584 27441 23612 28426
rect 23570 27432 23626 27441
rect 23570 27367 23626 27376
rect 23112 26784 23164 26790
rect 23112 26726 23164 26732
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 23124 23798 23152 26726
rect 23112 23792 23164 23798
rect 23112 23734 23164 23740
rect 23020 23724 23072 23730
rect 22940 23684 23020 23712
rect 23020 23666 23072 23672
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22376 22092 22428 22098
rect 22376 22034 22428 22040
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22388 18290 22416 19722
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22388 16658 22416 18226
rect 22376 16652 22428 16658
rect 22376 16594 22428 16600
rect 22376 13252 22428 13258
rect 22376 13194 22428 13200
rect 22388 12442 22416 13194
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22388 10810 22416 11698
rect 22480 11098 22508 22918
rect 23676 22658 23704 30534
rect 23768 28218 23796 32982
rect 23952 31754 23980 56306
rect 24964 55622 24992 56306
rect 25332 56234 25360 57394
rect 26608 56704 26660 56710
rect 26608 56646 26660 56652
rect 26620 56370 26648 56646
rect 26988 56506 27016 57394
rect 27620 57384 27672 57390
rect 27620 57326 27672 57332
rect 27632 56506 27660 57326
rect 26976 56500 27028 56506
rect 26976 56442 27028 56448
rect 27620 56500 27672 56506
rect 27620 56442 27672 56448
rect 25596 56364 25648 56370
rect 25596 56306 25648 56312
rect 26608 56364 26660 56370
rect 26608 56306 26660 56312
rect 27160 56364 27212 56370
rect 27160 56306 27212 56312
rect 25320 56228 25372 56234
rect 25320 56170 25372 56176
rect 25136 56160 25188 56166
rect 25136 56102 25188 56108
rect 25148 55962 25176 56102
rect 25136 55956 25188 55962
rect 25136 55898 25188 55904
rect 25608 55622 25636 56306
rect 26332 55752 26384 55758
rect 26332 55694 26384 55700
rect 24952 55616 25004 55622
rect 24952 55558 25004 55564
rect 25596 55616 25648 55622
rect 25596 55558 25648 55564
rect 26148 55616 26200 55622
rect 26148 55558 26200 55564
rect 24964 44985 24992 55558
rect 24950 44976 25006 44985
rect 24950 44911 25006 44920
rect 25320 41268 25372 41274
rect 25320 41210 25372 41216
rect 24400 41200 24452 41206
rect 24400 41142 24452 41148
rect 24412 40458 24440 41142
rect 24400 40452 24452 40458
rect 24400 40394 24452 40400
rect 24860 40452 24912 40458
rect 24860 40394 24912 40400
rect 24400 39432 24452 39438
rect 24400 39374 24452 39380
rect 24308 37868 24360 37874
rect 24412 37856 24440 39374
rect 24872 39302 24900 40394
rect 25228 39840 25280 39846
rect 25228 39782 25280 39788
rect 24860 39296 24912 39302
rect 24860 39238 24912 39244
rect 24360 37828 24440 37856
rect 24308 37810 24360 37816
rect 24412 37262 24440 37828
rect 24400 37256 24452 37262
rect 24400 37198 24452 37204
rect 24412 36854 24440 37198
rect 24676 37188 24728 37194
rect 24676 37130 24728 37136
rect 24400 36848 24452 36854
rect 24400 36790 24452 36796
rect 24688 36378 24716 37130
rect 24676 36372 24728 36378
rect 24676 36314 24728 36320
rect 24768 36304 24820 36310
rect 24768 36246 24820 36252
rect 24308 36236 24360 36242
rect 24308 36178 24360 36184
rect 24320 35494 24348 36178
rect 24676 36168 24728 36174
rect 24676 36110 24728 36116
rect 24688 35494 24716 36110
rect 24308 35488 24360 35494
rect 24308 35430 24360 35436
rect 24676 35488 24728 35494
rect 24676 35430 24728 35436
rect 24216 33040 24268 33046
rect 24216 32982 24268 32988
rect 24124 32564 24176 32570
rect 24124 32506 24176 32512
rect 24032 32428 24084 32434
rect 24032 32370 24084 32376
rect 23860 31726 23980 31754
rect 23756 28212 23808 28218
rect 23756 28154 23808 28160
rect 23756 27124 23808 27130
rect 23756 27066 23808 27072
rect 23768 23594 23796 27066
rect 23756 23588 23808 23594
rect 23756 23530 23808 23536
rect 23756 22976 23808 22982
rect 23756 22918 23808 22924
rect 23768 22778 23796 22918
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23676 22630 23796 22658
rect 23572 22568 23624 22574
rect 23572 22510 23624 22516
rect 22560 22432 22612 22438
rect 22560 22374 22612 22380
rect 22572 22030 22600 22374
rect 22652 22160 22704 22166
rect 22652 22102 22704 22108
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 22572 21418 22600 21966
rect 22560 21412 22612 21418
rect 22560 21354 22612 21360
rect 22664 20602 22692 22102
rect 23584 22098 23612 22510
rect 23664 22500 23716 22506
rect 23664 22442 23716 22448
rect 23572 22092 23624 22098
rect 23572 22034 23624 22040
rect 23480 22024 23532 22030
rect 23480 21966 23532 21972
rect 23020 21888 23072 21894
rect 23020 21830 23072 21836
rect 23032 21622 23060 21830
rect 23020 21616 23072 21622
rect 23020 21558 23072 21564
rect 23204 21344 23256 21350
rect 23204 21286 23256 21292
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 22836 20800 22888 20806
rect 22834 20768 22836 20777
rect 22888 20768 22890 20777
rect 22834 20703 22890 20712
rect 23124 20602 23152 20878
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23216 20482 23244 21286
rect 23492 21146 23520 21966
rect 23480 21140 23532 21146
rect 23480 21082 23532 21088
rect 23584 20942 23612 22034
rect 23676 21894 23704 22442
rect 23664 21888 23716 21894
rect 23664 21830 23716 21836
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 23480 20868 23532 20874
rect 23480 20810 23532 20816
rect 23388 20800 23440 20806
rect 23492 20777 23520 20810
rect 23388 20742 23440 20748
rect 23478 20768 23534 20777
rect 23124 20466 23244 20482
rect 23400 20466 23428 20742
rect 23478 20703 23534 20712
rect 23112 20460 23244 20466
rect 23164 20454 23244 20460
rect 23388 20460 23440 20466
rect 23112 20402 23164 20408
rect 23388 20402 23440 20408
rect 23584 20058 23612 20878
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23204 18216 23256 18222
rect 23204 18158 23256 18164
rect 23216 17746 23244 18158
rect 23204 17740 23256 17746
rect 23204 17682 23256 17688
rect 22928 17672 22980 17678
rect 22926 17640 22928 17649
rect 22980 17640 22982 17649
rect 22926 17575 22982 17584
rect 23296 17604 23348 17610
rect 23296 17546 23348 17552
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22572 16590 22600 17138
rect 23308 17134 23336 17546
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23480 17128 23532 17134
rect 23480 17070 23532 17076
rect 23388 16992 23440 16998
rect 23388 16934 23440 16940
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22572 15706 22600 16526
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22664 14498 22692 16594
rect 23204 15972 23256 15978
rect 23204 15914 23256 15920
rect 22744 15360 22796 15366
rect 22744 15302 22796 15308
rect 22756 15026 22784 15302
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 22836 14884 22888 14890
rect 22836 14826 22888 14832
rect 22572 14482 22692 14498
rect 22560 14476 22692 14482
rect 22612 14470 22692 14476
rect 22560 14418 22612 14424
rect 22572 14074 22600 14418
rect 22848 14414 22876 14826
rect 23216 14414 23244 15914
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 23308 15026 23336 15438
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 22652 14408 22704 14414
rect 22652 14350 22704 14356
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 22560 14068 22612 14074
rect 22560 14010 22612 14016
rect 22664 13938 22692 14350
rect 23216 13938 23244 14350
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23308 14006 23336 14282
rect 23296 14000 23348 14006
rect 23296 13942 23348 13948
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 23204 13932 23256 13938
rect 23204 13874 23256 13880
rect 22560 12368 22612 12374
rect 22560 12310 22612 12316
rect 22572 11762 22600 12310
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 23020 11144 23072 11150
rect 22480 11070 22600 11098
rect 23020 11086 23072 11092
rect 22468 11008 22520 11014
rect 22468 10950 22520 10956
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22480 10674 22508 10950
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22480 9722 22508 10610
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22572 9110 22600 11070
rect 23032 10674 23060 11086
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22848 10266 22876 10542
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22652 9580 22704 9586
rect 22928 9580 22980 9586
rect 22704 9540 22928 9568
rect 22652 9522 22704 9528
rect 22928 9522 22980 9528
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22664 6866 22692 9522
rect 23032 8498 23060 10610
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22756 7478 22784 7686
rect 22744 7472 22796 7478
rect 22744 7414 22796 7420
rect 22848 7410 22876 8434
rect 22836 7404 22888 7410
rect 22836 7346 22888 7352
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 22652 6860 22704 6866
rect 22652 6802 22704 6808
rect 22848 6254 22876 7346
rect 22836 6248 22888 6254
rect 22836 6190 22888 6196
rect 22848 5710 22876 6190
rect 22836 5704 22888 5710
rect 22836 5646 22888 5652
rect 22940 5642 22968 7346
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 23124 6118 23152 6258
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 23308 5914 23336 10610
rect 23400 9450 23428 16934
rect 23492 16114 23520 17070
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 23492 15706 23520 16050
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23492 13870 23520 14758
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23676 13977 23704 14010
rect 23662 13968 23718 13977
rect 23662 13903 23718 13912
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23572 13864 23624 13870
rect 23572 13806 23624 13812
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23492 11830 23520 12922
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23492 10742 23520 10950
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 23388 9444 23440 9450
rect 23388 9386 23440 9392
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23400 8498 23428 8774
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23584 8378 23612 13806
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23676 10810 23704 13466
rect 23768 13326 23796 22630
rect 23860 20618 23888 31726
rect 24044 30258 24072 32370
rect 24136 30326 24164 32506
rect 24124 30320 24176 30326
rect 24124 30262 24176 30268
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 24044 29170 24072 30194
rect 24032 29164 24084 29170
rect 24032 29106 24084 29112
rect 24044 27606 24072 29106
rect 24032 27600 24084 27606
rect 24032 27542 24084 27548
rect 24032 27396 24084 27402
rect 24032 27338 24084 27344
rect 24044 26994 24072 27338
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 24124 25832 24176 25838
rect 24124 25774 24176 25780
rect 24136 24070 24164 25774
rect 24124 24064 24176 24070
rect 24124 24006 24176 24012
rect 24124 23588 24176 23594
rect 24124 23530 24176 23536
rect 23940 22704 23992 22710
rect 23940 22646 23992 22652
rect 23952 21622 23980 22646
rect 24136 22642 24164 23530
rect 24124 22636 24176 22642
rect 24124 22578 24176 22584
rect 23940 21616 23992 21622
rect 23940 21558 23992 21564
rect 23860 20590 24072 20618
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 23860 18834 23888 20402
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23940 18828 23992 18834
rect 23940 18770 23992 18776
rect 23952 18358 23980 18770
rect 23940 18352 23992 18358
rect 23940 18294 23992 18300
rect 23940 14272 23992 14278
rect 23940 14214 23992 14220
rect 23952 14074 23980 14214
rect 23940 14068 23992 14074
rect 23940 14010 23992 14016
rect 23756 13320 23808 13326
rect 23756 13262 23808 13268
rect 23768 12986 23796 13262
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 24044 12617 24072 20590
rect 24228 15162 24256 32982
rect 24320 31414 24348 35430
rect 24780 35018 24808 36246
rect 24872 35698 24900 39238
rect 24952 37188 25004 37194
rect 24952 37130 25004 37136
rect 24964 36174 24992 37130
rect 25044 36576 25096 36582
rect 25044 36518 25096 36524
rect 25056 36174 25084 36518
rect 24952 36168 25004 36174
rect 24952 36110 25004 36116
rect 25044 36168 25096 36174
rect 25044 36110 25096 36116
rect 24860 35692 24912 35698
rect 24860 35634 24912 35640
rect 24768 35012 24820 35018
rect 24768 34954 24820 34960
rect 24676 34740 24728 34746
rect 24676 34682 24728 34688
rect 24400 34604 24452 34610
rect 24400 34546 24452 34552
rect 24412 33998 24440 34546
rect 24400 33992 24452 33998
rect 24400 33934 24452 33940
rect 24584 33992 24636 33998
rect 24584 33934 24636 33940
rect 24412 33522 24440 33934
rect 24400 33516 24452 33522
rect 24400 33458 24452 33464
rect 24412 31890 24440 33458
rect 24596 33114 24624 33934
rect 24688 33538 24716 34682
rect 24780 33658 24808 34954
rect 24964 34678 24992 36110
rect 25044 34944 25096 34950
rect 25044 34886 25096 34892
rect 24952 34672 25004 34678
rect 24952 34614 25004 34620
rect 24964 34066 24992 34614
rect 25056 34610 25084 34886
rect 25240 34610 25268 39782
rect 25332 35494 25360 41210
rect 25596 37664 25648 37670
rect 25596 37606 25648 37612
rect 25608 36718 25636 37606
rect 25688 36780 25740 36786
rect 25688 36722 25740 36728
rect 25596 36712 25648 36718
rect 25596 36654 25648 36660
rect 25608 36174 25636 36654
rect 25700 36310 25728 36722
rect 25688 36304 25740 36310
rect 25688 36246 25740 36252
rect 25596 36168 25648 36174
rect 25596 36110 25648 36116
rect 25700 36106 25728 36246
rect 25688 36100 25740 36106
rect 25688 36042 25740 36048
rect 25320 35488 25372 35494
rect 25320 35430 25372 35436
rect 25964 35488 26016 35494
rect 25964 35430 26016 35436
rect 25976 35290 26004 35430
rect 25964 35284 26016 35290
rect 25964 35226 26016 35232
rect 25504 35012 25556 35018
rect 25504 34954 25556 34960
rect 25516 34746 25544 34954
rect 25504 34740 25556 34746
rect 25504 34682 25556 34688
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 25228 34604 25280 34610
rect 25228 34546 25280 34552
rect 24952 34060 25004 34066
rect 24952 34002 25004 34008
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 24964 33590 24992 34002
rect 25044 33856 25096 33862
rect 25044 33798 25096 33804
rect 24952 33584 25004 33590
rect 24688 33522 24808 33538
rect 24952 33526 25004 33532
rect 24688 33516 24820 33522
rect 24688 33510 24768 33516
rect 24768 33458 24820 33464
rect 24584 33108 24636 33114
rect 24584 33050 24636 33056
rect 24400 31884 24452 31890
rect 24400 31826 24452 31832
rect 24676 31884 24728 31890
rect 24676 31826 24728 31832
rect 24400 31476 24452 31482
rect 24400 31418 24452 31424
rect 24308 31408 24360 31414
rect 24308 31350 24360 31356
rect 24412 30870 24440 31418
rect 24400 30864 24452 30870
rect 24400 30806 24452 30812
rect 24688 30734 24716 31826
rect 24676 30728 24728 30734
rect 24676 30670 24728 30676
rect 24688 29646 24716 30670
rect 24676 29640 24728 29646
rect 24676 29582 24728 29588
rect 24780 28762 24808 33458
rect 24860 33108 24912 33114
rect 24860 33050 24912 33056
rect 24872 29782 24900 33050
rect 24964 31890 24992 33526
rect 25056 32502 25084 33798
rect 25136 33448 25188 33454
rect 25136 33390 25188 33396
rect 25148 33114 25176 33390
rect 25136 33108 25188 33114
rect 25136 33050 25188 33056
rect 25044 32496 25096 32502
rect 25044 32438 25096 32444
rect 24952 31884 25004 31890
rect 24952 31826 25004 31832
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25240 30734 25268 31758
rect 25412 31136 25464 31142
rect 25412 31078 25464 31084
rect 25136 30728 25188 30734
rect 25136 30670 25188 30676
rect 25237 30728 25289 30734
rect 25237 30670 25289 30676
rect 24952 30592 25004 30598
rect 24952 30534 25004 30540
rect 24964 30258 24992 30534
rect 25148 30326 25176 30670
rect 25136 30320 25188 30326
rect 25136 30262 25188 30268
rect 24952 30252 25004 30258
rect 24952 30194 25004 30200
rect 24860 29776 24912 29782
rect 24860 29718 24912 29724
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24872 29306 24900 29582
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 24964 29102 24992 30194
rect 25240 29578 25268 30670
rect 25424 30258 25452 31078
rect 25412 30252 25464 30258
rect 25412 30194 25464 30200
rect 25504 30252 25556 30258
rect 25504 30194 25556 30200
rect 25424 29850 25452 30194
rect 25516 30054 25544 30194
rect 25976 30122 26004 35226
rect 26056 34604 26108 34610
rect 26056 34546 26108 34552
rect 25964 30116 26016 30122
rect 25964 30058 26016 30064
rect 25504 30048 25556 30054
rect 25504 29990 25556 29996
rect 25412 29844 25464 29850
rect 25412 29786 25464 29792
rect 25228 29572 25280 29578
rect 25228 29514 25280 29520
rect 25044 29504 25096 29510
rect 25044 29446 25096 29452
rect 24952 29096 25004 29102
rect 24952 29038 25004 29044
rect 25056 28948 25084 29446
rect 25516 29170 25544 29990
rect 25780 29504 25832 29510
rect 25780 29446 25832 29452
rect 25792 29238 25820 29446
rect 26068 29306 26096 34546
rect 26056 29300 26108 29306
rect 26056 29242 26108 29248
rect 25780 29232 25832 29238
rect 25780 29174 25832 29180
rect 25504 29164 25556 29170
rect 25504 29106 25556 29112
rect 24964 28920 25084 28948
rect 24768 28756 24820 28762
rect 24768 28698 24820 28704
rect 24768 27532 24820 27538
rect 24768 27474 24820 27480
rect 24492 27328 24544 27334
rect 24492 27270 24544 27276
rect 24308 26512 24360 26518
rect 24308 26454 24360 26460
rect 24320 23798 24348 26454
rect 24504 26450 24532 27270
rect 24676 26580 24728 26586
rect 24676 26522 24728 26528
rect 24492 26444 24544 26450
rect 24492 26386 24544 26392
rect 24688 26382 24716 26522
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24688 24818 24716 26318
rect 24780 26246 24808 27474
rect 24964 27470 24992 28920
rect 25516 28422 25544 29106
rect 25688 29028 25740 29034
rect 25688 28970 25740 28976
rect 25504 28416 25556 28422
rect 25504 28358 25556 28364
rect 25044 27872 25096 27878
rect 25044 27814 25096 27820
rect 25056 27470 25084 27814
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 25044 27464 25096 27470
rect 25044 27406 25096 27412
rect 25228 27464 25280 27470
rect 25228 27406 25280 27412
rect 25056 26518 25084 27406
rect 25044 26512 25096 26518
rect 25044 26454 25096 26460
rect 24860 26376 24912 26382
rect 24860 26318 24912 26324
rect 24768 26240 24820 26246
rect 24768 26182 24820 26188
rect 24676 24812 24728 24818
rect 24676 24754 24728 24760
rect 24780 24750 24808 26182
rect 24872 25498 24900 26318
rect 25240 26042 25268 27406
rect 25412 27056 25464 27062
rect 25412 26998 25464 27004
rect 25320 26988 25372 26994
rect 25320 26930 25372 26936
rect 25332 26586 25360 26930
rect 25320 26580 25372 26586
rect 25320 26522 25372 26528
rect 25228 26036 25280 26042
rect 25228 25978 25280 25984
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 24952 25288 25004 25294
rect 25424 25276 25452 26998
rect 25516 25770 25544 28358
rect 25700 26382 25728 28970
rect 25688 26376 25740 26382
rect 25688 26318 25740 26324
rect 25700 25974 25728 26318
rect 25688 25968 25740 25974
rect 25688 25910 25740 25916
rect 25504 25764 25556 25770
rect 25504 25706 25556 25712
rect 24952 25230 25004 25236
rect 25332 25248 25452 25276
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24308 23792 24360 23798
rect 24308 23734 24360 23740
rect 24320 22234 24348 23734
rect 24676 23656 24728 23662
rect 24676 23598 24728 23604
rect 24688 22574 24716 23598
rect 24780 23594 24808 24686
rect 24964 24206 24992 25230
rect 25044 24812 25096 24818
rect 25044 24754 25096 24760
rect 25056 24410 25084 24754
rect 25044 24404 25096 24410
rect 25044 24346 25096 24352
rect 25332 24290 25360 25248
rect 25504 24608 25556 24614
rect 25504 24550 25556 24556
rect 25056 24262 25360 24290
rect 24952 24200 25004 24206
rect 24952 24142 25004 24148
rect 24768 23588 24820 23594
rect 24768 23530 24820 23536
rect 24964 22778 24992 24142
rect 24952 22772 25004 22778
rect 24952 22714 25004 22720
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24676 22568 24728 22574
rect 24676 22510 24728 22516
rect 24308 22228 24360 22234
rect 24308 22170 24360 22176
rect 24320 22030 24348 22170
rect 24308 22024 24360 22030
rect 24308 21966 24360 21972
rect 24780 21078 24808 22578
rect 24768 21072 24820 21078
rect 24768 21014 24820 21020
rect 24584 20868 24636 20874
rect 24584 20810 24636 20816
rect 24596 20262 24624 20810
rect 24584 20256 24636 20262
rect 24584 20198 24636 20204
rect 24400 19848 24452 19854
rect 24400 19790 24452 19796
rect 24412 17678 24440 19790
rect 24596 18766 24624 20198
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 24584 18760 24636 18766
rect 24584 18702 24636 18708
rect 24688 18086 24716 19246
rect 24676 18080 24728 18086
rect 24676 18022 24728 18028
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24950 17640 25006 17649
rect 24780 17202 24808 17614
rect 24950 17575 25006 17584
rect 24964 17202 24992 17575
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 24306 15600 24362 15609
rect 24306 15535 24362 15544
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24136 14482 24164 14962
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 24228 14006 24256 15098
rect 24320 14278 24348 15535
rect 25056 15162 25084 24262
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25424 23186 25452 24142
rect 25516 24138 25544 24550
rect 25504 24132 25556 24138
rect 25504 24074 25556 24080
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25412 23180 25464 23186
rect 25412 23122 25464 23128
rect 25608 22778 25636 23666
rect 25872 23520 25924 23526
rect 25872 23462 25924 23468
rect 25884 23118 25912 23462
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25596 22772 25648 22778
rect 25596 22714 25648 22720
rect 25872 22704 25924 22710
rect 25872 22646 25924 22652
rect 25228 20800 25280 20806
rect 25228 20742 25280 20748
rect 25240 20534 25268 20742
rect 25228 20528 25280 20534
rect 25226 20496 25228 20505
rect 25280 20496 25282 20505
rect 25884 20466 25912 22646
rect 25964 22092 26016 22098
rect 26160 22094 26188 55558
rect 26344 42129 26372 55694
rect 26330 42120 26386 42129
rect 26330 42055 26386 42064
rect 26516 37936 26568 37942
rect 26516 37878 26568 37884
rect 26240 37868 26292 37874
rect 26240 37810 26292 37816
rect 26252 37466 26280 37810
rect 26528 37738 26556 37878
rect 26516 37732 26568 37738
rect 26516 37674 26568 37680
rect 26240 37460 26292 37466
rect 26240 37402 26292 37408
rect 26528 37262 26556 37674
rect 26516 37256 26568 37262
rect 26516 37198 26568 37204
rect 26240 37120 26292 37126
rect 26240 37062 26292 37068
rect 26252 36786 26280 37062
rect 26240 36780 26292 36786
rect 26240 36722 26292 36728
rect 26240 33380 26292 33386
rect 26240 33322 26292 33328
rect 26252 32910 26280 33322
rect 26240 32904 26292 32910
rect 26240 32846 26292 32852
rect 26516 32904 26568 32910
rect 26516 32846 26568 32852
rect 26528 32434 26556 32846
rect 26516 32428 26568 32434
rect 26516 32370 26568 32376
rect 26424 28960 26476 28966
rect 26424 28902 26476 28908
rect 26436 28558 26464 28902
rect 26424 28552 26476 28558
rect 26424 28494 26476 28500
rect 26424 26988 26476 26994
rect 26424 26930 26476 26936
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26252 25226 26280 26726
rect 26436 26586 26464 26930
rect 26424 26580 26476 26586
rect 26424 26522 26476 26528
rect 26332 26308 26384 26314
rect 26332 26250 26384 26256
rect 26344 25974 26372 26250
rect 26332 25968 26384 25974
rect 26332 25910 26384 25916
rect 26344 25294 26372 25910
rect 26332 25288 26384 25294
rect 26332 25230 26384 25236
rect 26240 25220 26292 25226
rect 26240 25162 26292 25168
rect 26252 23118 26280 25162
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 25964 22034 26016 22040
rect 26068 22066 26188 22094
rect 25976 21690 26004 22034
rect 25964 21684 26016 21690
rect 25964 21626 26016 21632
rect 25226 20431 25282 20440
rect 25872 20460 25924 20466
rect 25240 20405 25268 20431
rect 25872 20402 25924 20408
rect 25688 19848 25740 19854
rect 25688 19790 25740 19796
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25596 18760 25648 18766
rect 25700 18748 25728 19790
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25792 18970 25820 19110
rect 25780 18964 25832 18970
rect 25780 18906 25832 18912
rect 25648 18720 25728 18748
rect 25596 18702 25648 18708
rect 25424 18630 25452 18702
rect 25504 18692 25556 18698
rect 25504 18634 25556 18640
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25136 17808 25188 17814
rect 25136 17750 25188 17756
rect 25148 16998 25176 17750
rect 25424 17746 25452 18566
rect 25516 18426 25544 18634
rect 25504 18420 25556 18426
rect 25504 18362 25556 18368
rect 25412 17740 25464 17746
rect 25412 17682 25464 17688
rect 25608 17678 25636 18702
rect 25964 18420 26016 18426
rect 25964 18362 26016 18368
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25700 17882 25728 18226
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25596 17672 25648 17678
rect 25596 17614 25648 17620
rect 25872 17604 25924 17610
rect 25872 17546 25924 17552
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25700 17066 25728 17274
rect 25884 17134 25912 17546
rect 25976 17270 26004 18362
rect 25964 17264 26016 17270
rect 25964 17206 26016 17212
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 25688 17060 25740 17066
rect 25688 17002 25740 17008
rect 25136 16992 25188 16998
rect 25136 16934 25188 16940
rect 25884 16794 25912 17070
rect 25872 16788 25924 16794
rect 25872 16730 25924 16736
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 25596 15156 25648 15162
rect 25596 15098 25648 15104
rect 24952 14544 25004 14550
rect 24952 14486 25004 14492
rect 24400 14476 24452 14482
rect 24400 14418 24452 14424
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24216 14000 24268 14006
rect 24216 13942 24268 13948
rect 24030 12608 24086 12617
rect 24030 12543 24086 12552
rect 24412 12434 24440 14418
rect 24768 14408 24820 14414
rect 24768 14350 24820 14356
rect 24584 14068 24636 14074
rect 24584 14010 24636 14016
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 24228 12406 24440 12434
rect 23848 11892 23900 11898
rect 23848 11834 23900 11840
rect 23860 11218 23888 11834
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24136 11218 24164 11494
rect 23848 11212 23900 11218
rect 23848 11154 23900 11160
rect 24124 11212 24176 11218
rect 24124 11154 24176 11160
rect 24228 10826 24256 12406
rect 24504 12186 24532 13874
rect 24596 13841 24624 14010
rect 24582 13832 24638 13841
rect 24582 13767 24638 13776
rect 24780 13462 24808 14350
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24768 13456 24820 13462
rect 24768 13398 24820 13404
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 23664 10804 23716 10810
rect 23664 10746 23716 10752
rect 24136 10798 24256 10826
rect 24320 12158 24532 12186
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23492 8350 23612 8378
rect 23400 6798 23428 8298
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23400 6118 23428 6734
rect 23492 6458 23520 8350
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23584 7886 23612 8230
rect 23952 8090 23980 8434
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 24136 7546 24164 10798
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24228 8566 24256 10610
rect 24320 10198 24348 12158
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24504 11626 24532 11834
rect 24492 11620 24544 11626
rect 24492 11562 24544 11568
rect 24504 10606 24532 11562
rect 24596 11150 24624 13330
rect 24872 11200 24900 13806
rect 24964 13734 24992 14486
rect 25056 14414 25084 15098
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25608 14074 25636 15098
rect 25596 14068 25648 14074
rect 25596 14010 25648 14016
rect 25608 13938 25636 14010
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25872 13796 25924 13802
rect 25872 13738 25924 13744
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 25504 13252 25556 13258
rect 25504 13194 25556 13200
rect 25516 12646 25544 13194
rect 25504 12640 25556 12646
rect 25504 12582 25556 12588
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 25056 11354 25084 12174
rect 25136 12164 25188 12170
rect 25136 12106 25188 12112
rect 25148 11898 25176 12106
rect 25136 11892 25188 11898
rect 25136 11834 25188 11840
rect 25596 11756 25648 11762
rect 25596 11698 25648 11704
rect 25608 11354 25636 11698
rect 25044 11348 25096 11354
rect 25044 11290 25096 11296
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 24780 11172 24900 11200
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24308 10192 24360 10198
rect 24308 10134 24360 10140
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24216 8560 24268 8566
rect 24216 8502 24268 8508
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24228 7478 24256 8502
rect 24216 7472 24268 7478
rect 24216 7414 24268 7420
rect 23664 7200 23716 7206
rect 23664 7142 23716 7148
rect 23676 6798 23704 7142
rect 23940 6928 23992 6934
rect 23940 6870 23992 6876
rect 23952 6798 23980 6870
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23940 6792 23992 6798
rect 23940 6734 23992 6740
rect 24228 6730 24256 7414
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24216 6724 24268 6730
rect 24216 6666 24268 6672
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 23400 5778 23428 6054
rect 23388 5772 23440 5778
rect 23388 5714 23440 5720
rect 22928 5636 22980 5642
rect 22928 5578 22980 5584
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22376 4480 22428 4486
rect 22376 4422 22428 4428
rect 22284 3188 22336 3194
rect 22284 3130 22336 3136
rect 22388 2446 22416 4422
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 22480 2582 22508 4218
rect 22468 2576 22520 2582
rect 22468 2518 22520 2524
rect 22376 2440 22428 2446
rect 22428 2400 22508 2428
rect 22376 2382 22428 2388
rect 22204 2332 22324 2360
rect 22020 2038 22048 2246
rect 22112 2230 22232 2258
rect 22008 2032 22060 2038
rect 22008 1974 22060 1980
rect 21928 1550 22048 1578
rect 21836 1414 21956 1442
rect 21928 800 21956 1414
rect 22020 800 22048 1550
rect 22204 800 22232 2230
rect 22296 800 22324 2332
rect 22480 800 22508 2400
rect 22572 800 22600 4966
rect 22940 4826 22968 5578
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 23020 5024 23072 5030
rect 23020 4966 23072 4972
rect 22928 4820 22980 4826
rect 22928 4762 22980 4768
rect 22928 3936 22980 3942
rect 22928 3878 22980 3884
rect 22836 3392 22888 3398
rect 22836 3334 22888 3340
rect 22848 3058 22876 3334
rect 22836 3052 22888 3058
rect 22836 2994 22888 3000
rect 22848 2938 22876 2994
rect 22756 2910 22876 2938
rect 22756 800 22784 2910
rect 22940 2836 22968 3878
rect 22848 2808 22968 2836
rect 22848 800 22876 2808
rect 23032 2774 23060 4966
rect 23204 4820 23256 4826
rect 23204 4762 23256 4768
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 22940 2746 23060 2774
rect 22940 2582 22968 2746
rect 22928 2576 22980 2582
rect 22928 2518 22980 2524
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 23032 2310 23060 2382
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 23032 800 23060 2246
rect 23124 800 23152 3878
rect 23216 3194 23244 4762
rect 23296 4548 23348 4554
rect 23296 4490 23348 4496
rect 23204 3188 23256 3194
rect 23204 3130 23256 3136
rect 23308 2922 23336 4490
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23296 2916 23348 2922
rect 23296 2858 23348 2864
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23308 800 23336 2382
rect 23400 800 23428 3878
rect 23492 2854 23520 5510
rect 23584 4622 23612 6598
rect 23756 6384 23808 6390
rect 23756 6326 23808 6332
rect 23768 5710 23796 6326
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23768 5370 23796 5646
rect 24412 5642 24440 7346
rect 24504 6780 24532 10066
rect 24596 8498 24624 11086
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24688 10606 24716 10950
rect 24780 10742 24808 11172
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24768 10736 24820 10742
rect 24768 10678 24820 10684
rect 24872 10674 24900 11018
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24688 10062 24716 10542
rect 24964 10266 24992 11086
rect 25056 10674 25084 11290
rect 25412 11008 25464 11014
rect 25412 10950 25464 10956
rect 25424 10742 25452 10950
rect 25412 10736 25464 10742
rect 25412 10678 25464 10684
rect 25044 10668 25096 10674
rect 25044 10610 25096 10616
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 24952 10260 25004 10266
rect 24952 10202 25004 10208
rect 25424 10062 25452 10406
rect 24676 10056 24728 10062
rect 24676 9998 24728 10004
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 24596 7410 24624 8434
rect 24688 7818 24716 9862
rect 25412 9580 25464 9586
rect 25412 9522 25464 9528
rect 25424 9178 25452 9522
rect 25412 9172 25464 9178
rect 25412 9114 25464 9120
rect 25884 7886 25912 13738
rect 26068 12434 26096 22066
rect 26344 21146 26372 22918
rect 26620 22094 26648 56306
rect 27172 44849 27200 56306
rect 28460 55894 28488 57394
rect 30024 56778 30052 57394
rect 30380 57384 30432 57390
rect 30380 57326 30432 57332
rect 30012 56772 30064 56778
rect 30012 56714 30064 56720
rect 30392 56506 30420 57326
rect 33244 56506 33272 57394
rect 34808 56506 34836 57394
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 30380 56500 30432 56506
rect 30380 56442 30432 56448
rect 33232 56500 33284 56506
rect 33232 56442 33284 56448
rect 34796 56500 34848 56506
rect 34796 56442 34848 56448
rect 29644 56364 29696 56370
rect 29644 56306 29696 56312
rect 31668 56364 31720 56370
rect 31668 56306 31720 56312
rect 32128 56364 32180 56370
rect 32128 56306 32180 56312
rect 33968 56364 34020 56370
rect 33968 56306 34020 56312
rect 35808 56364 35860 56370
rect 35808 56306 35860 56312
rect 28448 55888 28500 55894
rect 28448 55830 28500 55836
rect 29656 53145 29684 56306
rect 29642 53136 29698 53145
rect 29642 53071 29698 53080
rect 27158 44840 27214 44849
rect 27158 44775 27214 44784
rect 30840 40452 30892 40458
rect 30840 40394 30892 40400
rect 29184 40180 29236 40186
rect 29184 40122 29236 40128
rect 28356 40044 28408 40050
rect 28356 39986 28408 39992
rect 27620 39840 27672 39846
rect 27620 39782 27672 39788
rect 27632 39370 27660 39782
rect 27252 39364 27304 39370
rect 27252 39306 27304 39312
rect 27620 39364 27672 39370
rect 27620 39306 27672 39312
rect 26976 38752 27028 38758
rect 26976 38694 27028 38700
rect 26700 37256 26752 37262
rect 26700 37198 26752 37204
rect 26884 37256 26936 37262
rect 26884 37198 26936 37204
rect 26712 36378 26740 37198
rect 26700 36372 26752 36378
rect 26700 36314 26752 36320
rect 26896 36242 26924 37198
rect 26884 36236 26936 36242
rect 26884 36178 26936 36184
rect 26988 28762 27016 38694
rect 27264 38554 27292 39306
rect 27632 38758 27660 39306
rect 27620 38752 27672 38758
rect 27620 38694 27672 38700
rect 27252 38548 27304 38554
rect 27252 38490 27304 38496
rect 27068 38208 27120 38214
rect 27068 38150 27120 38156
rect 27080 34354 27108 38150
rect 27436 37732 27488 37738
rect 27436 37674 27488 37680
rect 27160 36032 27212 36038
rect 27160 35974 27212 35980
rect 27172 34474 27200 35974
rect 27160 34468 27212 34474
rect 27160 34410 27212 34416
rect 27080 34326 27200 34354
rect 27172 33522 27200 34326
rect 27160 33516 27212 33522
rect 27160 33458 27212 33464
rect 27172 33318 27200 33458
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 27172 32026 27200 33254
rect 27448 32298 27476 37674
rect 27632 36786 27660 38694
rect 28368 38554 28396 39986
rect 28816 39296 28868 39302
rect 28816 39238 28868 39244
rect 29000 39296 29052 39302
rect 29000 39238 29052 39244
rect 28356 38548 28408 38554
rect 28356 38490 28408 38496
rect 27712 38344 27764 38350
rect 27712 38286 27764 38292
rect 27988 38344 28040 38350
rect 27988 38286 28040 38292
rect 27724 38010 27752 38286
rect 27712 38004 27764 38010
rect 27712 37946 27764 37952
rect 28000 37126 28028 38286
rect 28828 37942 28856 39238
rect 29012 38962 29040 39238
rect 29000 38956 29052 38962
rect 29000 38898 29052 38904
rect 28908 38344 28960 38350
rect 28908 38286 28960 38292
rect 28920 38010 28948 38286
rect 28908 38004 28960 38010
rect 28908 37946 28960 37952
rect 28816 37936 28868 37942
rect 28816 37878 28868 37884
rect 27988 37120 28040 37126
rect 27988 37062 28040 37068
rect 27620 36780 27672 36786
rect 27620 36722 27672 36728
rect 27712 36780 27764 36786
rect 27712 36722 27764 36728
rect 27724 36378 27752 36722
rect 27712 36372 27764 36378
rect 27712 36314 27764 36320
rect 28000 36174 28028 37062
rect 27988 36168 28040 36174
rect 27988 36110 28040 36116
rect 28172 36168 28224 36174
rect 28172 36110 28224 36116
rect 27896 36100 27948 36106
rect 27896 36042 27948 36048
rect 27908 35834 27936 36042
rect 28184 35834 28212 36110
rect 27896 35828 27948 35834
rect 27896 35770 27948 35776
rect 28172 35828 28224 35834
rect 28172 35770 28224 35776
rect 28632 35828 28684 35834
rect 28632 35770 28684 35776
rect 27528 35080 27580 35086
rect 27528 35022 27580 35028
rect 27540 33998 27568 35022
rect 27908 34202 27936 35770
rect 27896 34196 27948 34202
rect 27896 34138 27948 34144
rect 28356 34196 28408 34202
rect 28356 34138 28408 34144
rect 27528 33992 27580 33998
rect 27528 33934 27580 33940
rect 27540 32774 27568 33934
rect 27712 33924 27764 33930
rect 27712 33866 27764 33872
rect 27724 33658 27752 33866
rect 27712 33652 27764 33658
rect 27712 33594 27764 33600
rect 28368 33522 28396 34138
rect 28356 33516 28408 33522
rect 28356 33458 28408 33464
rect 27528 32768 27580 32774
rect 27528 32710 27580 32716
rect 27436 32292 27488 32298
rect 27436 32234 27488 32240
rect 27160 32020 27212 32026
rect 27160 31962 27212 31968
rect 27448 30190 27476 32234
rect 27540 30802 27568 32710
rect 27712 32224 27764 32230
rect 27712 32166 27764 32172
rect 27528 30796 27580 30802
rect 27528 30738 27580 30744
rect 27436 30184 27488 30190
rect 27436 30126 27488 30132
rect 27540 29714 27568 30738
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 27618 29064 27674 29073
rect 27618 28999 27620 29008
rect 27672 28999 27674 29008
rect 27620 28970 27672 28976
rect 26976 28756 27028 28762
rect 26976 28698 27028 28704
rect 26700 28416 26752 28422
rect 26700 28358 26752 28364
rect 26528 22066 26648 22094
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 26240 20800 26292 20806
rect 26292 20760 26464 20788
rect 26240 20742 26292 20748
rect 26332 19984 26384 19990
rect 26332 19926 26384 19932
rect 26240 19236 26292 19242
rect 26240 19178 26292 19184
rect 26148 18964 26200 18970
rect 26148 18906 26200 18912
rect 26160 18630 26188 18906
rect 26252 18834 26280 19178
rect 26240 18828 26292 18834
rect 26240 18770 26292 18776
rect 26148 18624 26200 18630
rect 26148 18566 26200 18572
rect 26148 17672 26200 17678
rect 26148 17614 26200 17620
rect 26160 17338 26188 17614
rect 26148 17332 26200 17338
rect 26148 17274 26200 17280
rect 26252 16182 26280 18770
rect 26344 18766 26372 19926
rect 26332 18760 26384 18766
rect 26332 18702 26384 18708
rect 26332 18420 26384 18426
rect 26332 18362 26384 18368
rect 26344 16250 26372 18362
rect 26332 16244 26384 16250
rect 26332 16186 26384 16192
rect 26240 16176 26292 16182
rect 26240 16118 26292 16124
rect 26148 13932 26200 13938
rect 26148 13874 26200 13880
rect 26160 12918 26188 13874
rect 26148 12912 26200 12918
rect 26148 12854 26200 12860
rect 25976 12406 26096 12434
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25872 7880 25924 7886
rect 25872 7822 25924 7828
rect 24676 7812 24728 7818
rect 24676 7754 24728 7760
rect 24688 7546 24716 7754
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 24596 6934 24624 7346
rect 24688 7342 24716 7482
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 24584 6928 24636 6934
rect 24584 6870 24636 6876
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 24584 6792 24636 6798
rect 24504 6752 24584 6780
rect 24584 6734 24636 6740
rect 24596 6254 24624 6734
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24780 5914 24808 6598
rect 24860 6316 24912 6322
rect 24860 6258 24912 6264
rect 24768 5908 24820 5914
rect 24768 5850 24820 5856
rect 24400 5636 24452 5642
rect 24400 5578 24452 5584
rect 24872 5574 24900 6258
rect 24860 5568 24912 5574
rect 24860 5510 24912 5516
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 24964 5302 24992 6802
rect 24952 5296 25004 5302
rect 24952 5238 25004 5244
rect 25148 5234 25176 7822
rect 25596 7812 25648 7818
rect 25596 7754 25648 7760
rect 25608 7546 25636 7754
rect 25596 7540 25648 7546
rect 25596 7482 25648 7488
rect 25320 7404 25372 7410
rect 25976 7392 26004 12406
rect 26160 12238 26188 12854
rect 26252 12850 26280 16118
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26056 12096 26108 12102
rect 26056 12038 26108 12044
rect 26068 11150 26096 12038
rect 26148 11824 26200 11830
rect 26148 11766 26200 11772
rect 26160 11150 26188 11766
rect 26056 11144 26108 11150
rect 26056 11086 26108 11092
rect 26148 11144 26200 11150
rect 26148 11086 26200 11092
rect 26068 9654 26096 11086
rect 26240 11076 26292 11082
rect 26240 11018 26292 11024
rect 26252 10674 26280 11018
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26056 9648 26108 9654
rect 26056 9590 26108 9596
rect 26332 8492 26384 8498
rect 26332 8434 26384 8440
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26252 7478 26280 8026
rect 26240 7472 26292 7478
rect 26240 7414 26292 7420
rect 25320 7346 25372 7352
rect 25884 7364 26004 7392
rect 25332 7274 25360 7346
rect 25320 7268 25372 7274
rect 25320 7210 25372 7216
rect 25596 6180 25648 6186
rect 25596 6122 25648 6128
rect 25608 5778 25636 6122
rect 25596 5772 25648 5778
rect 25596 5714 25648 5720
rect 25608 5370 25636 5714
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 25148 4690 25176 5170
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 23572 4616 23624 4622
rect 23572 4558 23624 4564
rect 23768 4554 23980 4570
rect 23756 4548 23992 4554
rect 23808 4542 23940 4548
rect 23756 4490 23808 4496
rect 23940 4490 23992 4496
rect 24400 4480 24452 4486
rect 24400 4422 24452 4428
rect 24216 3936 24268 3942
rect 24216 3878 24268 3884
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 23940 3528 23992 3534
rect 23940 3470 23992 3476
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23676 800 23704 3470
rect 23952 800 23980 3470
rect 24228 800 24256 3878
rect 24412 3126 24440 4422
rect 25884 4282 25912 7364
rect 25962 7168 26018 7177
rect 25962 7103 26018 7112
rect 25976 6866 26004 7103
rect 25964 6860 26016 6866
rect 25964 6802 26016 6808
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 26160 5234 26188 6054
rect 26148 5228 26200 5234
rect 26148 5170 26200 5176
rect 25872 4276 25924 4282
rect 25872 4218 25924 4224
rect 25320 3936 25372 3942
rect 25320 3878 25372 3884
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 24400 3120 24452 3126
rect 24400 3062 24452 3068
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24504 800 24532 2926
rect 24780 800 24808 3470
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 25056 800 25084 2790
rect 25332 800 25360 3878
rect 26160 3670 26188 5170
rect 26344 4078 26372 8434
rect 26436 4758 26464 20760
rect 26424 4752 26476 4758
rect 26424 4694 26476 4700
rect 26436 4214 26464 4694
rect 26424 4208 26476 4214
rect 26424 4150 26476 4156
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26148 3664 26200 3670
rect 26148 3606 26200 3612
rect 25596 3528 25648 3534
rect 25596 3470 25648 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 25412 2644 25464 2650
rect 25412 2586 25464 2592
rect 25424 2106 25452 2586
rect 25412 2100 25464 2106
rect 25412 2042 25464 2048
rect 25608 800 25636 3470
rect 25872 2848 25924 2854
rect 25872 2790 25924 2796
rect 25884 800 25912 2790
rect 26160 800 26188 3470
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26240 2508 26292 2514
rect 26240 2450 26292 2456
rect 26252 2106 26280 2450
rect 26240 2100 26292 2106
rect 26240 2042 26292 2048
rect 26436 800 26464 2926
rect 26528 2514 26556 22066
rect 26608 22024 26660 22030
rect 26608 21966 26660 21972
rect 26620 21486 26648 21966
rect 26712 21554 26740 28358
rect 26884 28076 26936 28082
rect 26884 28018 26936 28024
rect 26792 24404 26844 24410
rect 26792 24346 26844 24352
rect 26804 24070 26832 24346
rect 26792 24064 26844 24070
rect 26792 24006 26844 24012
rect 26896 23882 26924 28018
rect 26988 26382 27016 28698
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27620 28552 27672 28558
rect 27620 28494 27672 28500
rect 27068 28484 27120 28490
rect 27068 28426 27120 28432
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 26988 26042 27016 26318
rect 26976 26036 27028 26042
rect 26976 25978 27028 25984
rect 26804 23854 26924 23882
rect 26700 21548 26752 21554
rect 26700 21490 26752 21496
rect 26608 21480 26660 21486
rect 26608 21422 26660 21428
rect 26620 20942 26648 21422
rect 26700 21140 26752 21146
rect 26700 21082 26752 21088
rect 26608 20936 26660 20942
rect 26608 20878 26660 20884
rect 26620 19718 26648 20878
rect 26608 19712 26660 19718
rect 26608 19654 26660 19660
rect 26712 19394 26740 21082
rect 26620 19366 26740 19394
rect 26620 17678 26648 19366
rect 26700 19304 26752 19310
rect 26700 19246 26752 19252
rect 26608 17672 26660 17678
rect 26608 17614 26660 17620
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 26620 10130 26648 14010
rect 26608 10124 26660 10130
rect 26608 10066 26660 10072
rect 26712 9450 26740 19246
rect 26804 18698 26832 23854
rect 27080 22094 27108 28426
rect 26896 22066 27108 22094
rect 26896 21894 26924 22066
rect 26884 21888 26936 21894
rect 26884 21830 26936 21836
rect 26896 20806 26924 21830
rect 27172 21010 27200 28494
rect 27632 27470 27660 28494
rect 27620 27464 27672 27470
rect 27620 27406 27672 27412
rect 27632 26926 27660 27406
rect 27620 26920 27672 26926
rect 27620 26862 27672 26868
rect 27632 25702 27660 26862
rect 27620 25696 27672 25702
rect 27620 25638 27672 25644
rect 27528 24948 27580 24954
rect 27528 24890 27580 24896
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27356 22710 27384 22918
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 27160 21004 27212 21010
rect 27160 20946 27212 20952
rect 27264 20942 27292 21286
rect 27252 20936 27304 20942
rect 27252 20878 27304 20884
rect 26976 20868 27028 20874
rect 26976 20810 27028 20816
rect 26884 20800 26936 20806
rect 26884 20742 26936 20748
rect 26988 20602 27016 20810
rect 27252 20800 27304 20806
rect 27252 20742 27304 20748
rect 26976 20596 27028 20602
rect 26976 20538 27028 20544
rect 27264 20466 27292 20742
rect 27068 20460 27120 20466
rect 27068 20402 27120 20408
rect 27252 20460 27304 20466
rect 27252 20402 27304 20408
rect 26884 20324 26936 20330
rect 26884 20266 26936 20272
rect 26896 19514 26924 20266
rect 26884 19508 26936 19514
rect 26884 19450 26936 19456
rect 26792 18692 26844 18698
rect 26792 18634 26844 18640
rect 27080 18630 27108 20402
rect 27160 19984 27212 19990
rect 27160 19926 27212 19932
rect 27172 19378 27200 19926
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 27068 18624 27120 18630
rect 27068 18566 27120 18572
rect 26976 17808 27028 17814
rect 26976 17750 27028 17756
rect 26988 17649 27016 17750
rect 26974 17640 27030 17649
rect 26974 17575 27030 17584
rect 27068 17604 27120 17610
rect 27068 17546 27120 17552
rect 26884 17536 26936 17542
rect 26884 17478 26936 17484
rect 26896 17338 26924 17478
rect 26884 17332 26936 17338
rect 26884 17274 26936 17280
rect 26976 17196 27028 17202
rect 26976 17138 27028 17144
rect 26988 16250 27016 17138
rect 27080 16436 27108 17546
rect 27264 16658 27292 19654
rect 27356 19378 27384 22646
rect 27436 21480 27488 21486
rect 27436 21422 27488 21428
rect 27448 20330 27476 21422
rect 27436 20324 27488 20330
rect 27436 20266 27488 20272
rect 27436 19780 27488 19786
rect 27436 19722 27488 19728
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27448 19242 27476 19722
rect 27540 19446 27568 24890
rect 27632 24206 27660 25638
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 27632 23798 27660 24142
rect 27620 23792 27672 23798
rect 27620 23734 27672 23740
rect 27724 22094 27752 32166
rect 28540 31952 28592 31958
rect 28540 31894 28592 31900
rect 27896 30252 27948 30258
rect 27896 30194 27948 30200
rect 27908 30054 27936 30194
rect 28264 30116 28316 30122
rect 28264 30058 28316 30064
rect 27896 30048 27948 30054
rect 27896 29990 27948 29996
rect 27908 27946 27936 29990
rect 28276 29646 28304 30058
rect 28448 30048 28500 30054
rect 28448 29990 28500 29996
rect 28356 29844 28408 29850
rect 28356 29786 28408 29792
rect 28264 29640 28316 29646
rect 28264 29582 28316 29588
rect 27896 27940 27948 27946
rect 27896 27882 27948 27888
rect 28264 25152 28316 25158
rect 28264 25094 28316 25100
rect 27988 24880 28040 24886
rect 27988 24822 28040 24828
rect 27804 24268 27856 24274
rect 27804 24210 27856 24216
rect 27816 24138 27844 24210
rect 28000 24138 28028 24822
rect 28276 24614 28304 25094
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 28276 24342 28304 24550
rect 28264 24336 28316 24342
rect 28264 24278 28316 24284
rect 27804 24132 27856 24138
rect 27804 24074 27856 24080
rect 27988 24132 28040 24138
rect 27988 24074 28040 24080
rect 27816 22778 27844 24074
rect 28000 23866 28028 24074
rect 28172 24064 28224 24070
rect 28172 24006 28224 24012
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 27804 22772 27856 22778
rect 27804 22714 27856 22720
rect 28184 22642 28212 24006
rect 28172 22636 28224 22642
rect 28172 22578 28224 22584
rect 28080 22432 28132 22438
rect 28080 22374 28132 22380
rect 27632 22066 27752 22094
rect 27528 19440 27580 19446
rect 27528 19382 27580 19388
rect 27436 19236 27488 19242
rect 27436 19178 27488 19184
rect 27436 18692 27488 18698
rect 27436 18634 27488 18640
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27344 16652 27396 16658
rect 27344 16594 27396 16600
rect 27160 16448 27212 16454
rect 27080 16408 27160 16436
rect 26976 16244 27028 16250
rect 26976 16186 27028 16192
rect 27080 15706 27108 16408
rect 27160 16390 27212 16396
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27172 15978 27200 16050
rect 27160 15972 27212 15978
rect 27160 15914 27212 15920
rect 27068 15700 27120 15706
rect 27068 15642 27120 15648
rect 27172 15502 27200 15914
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 26988 14822 27016 15438
rect 26976 14816 27028 14822
rect 26976 14758 27028 14764
rect 26988 14550 27016 14758
rect 26976 14544 27028 14550
rect 26976 14486 27028 14492
rect 26976 14408 27028 14414
rect 26976 14350 27028 14356
rect 26988 13938 27016 14350
rect 26976 13932 27028 13938
rect 26976 13874 27028 13880
rect 27252 13932 27304 13938
rect 27252 13874 27304 13880
rect 27264 13530 27292 13874
rect 27252 13524 27304 13530
rect 27252 13466 27304 13472
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26700 9444 26752 9450
rect 26700 9386 26752 9392
rect 26804 8362 26832 13126
rect 27068 12844 27120 12850
rect 27068 12786 27120 12792
rect 27080 10538 27108 12786
rect 27356 12782 27384 16594
rect 27344 12776 27396 12782
rect 27344 12718 27396 12724
rect 27448 12434 27476 18634
rect 27528 16040 27580 16046
rect 27528 15982 27580 15988
rect 27540 15473 27568 15982
rect 27526 15464 27582 15473
rect 27526 15399 27582 15408
rect 27632 15162 27660 22066
rect 27712 21956 27764 21962
rect 27712 21898 27764 21904
rect 27724 21690 27752 21898
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 28092 21554 28120 22374
rect 28276 22094 28304 24278
rect 28184 22066 28304 22094
rect 28368 22094 28396 29786
rect 28460 28558 28488 29990
rect 28552 29646 28580 31894
rect 28644 30258 28672 35770
rect 28828 32434 28856 37878
rect 29012 36854 29040 38898
rect 29196 37874 29224 40122
rect 30852 39642 30880 40394
rect 30840 39636 30892 39642
rect 30840 39578 30892 39584
rect 31576 39432 31628 39438
rect 31576 39374 31628 39380
rect 30380 39296 30432 39302
rect 30380 39238 30432 39244
rect 31116 39296 31168 39302
rect 31116 39238 31168 39244
rect 31484 39296 31536 39302
rect 31484 39238 31536 39244
rect 30196 38956 30248 38962
rect 30196 38898 30248 38904
rect 29736 38752 29788 38758
rect 29736 38694 29788 38700
rect 29276 38344 29328 38350
rect 29276 38286 29328 38292
rect 29288 37942 29316 38286
rect 29276 37936 29328 37942
rect 29276 37878 29328 37884
rect 29184 37868 29236 37874
rect 29184 37810 29236 37816
rect 29000 36848 29052 36854
rect 29000 36790 29052 36796
rect 28908 36780 28960 36786
rect 28908 36722 28960 36728
rect 28920 36106 28948 36722
rect 28908 36100 28960 36106
rect 28908 36042 28960 36048
rect 29092 33856 29144 33862
rect 29092 33798 29144 33804
rect 29104 33522 29132 33798
rect 29092 33516 29144 33522
rect 29092 33458 29144 33464
rect 29000 32836 29052 32842
rect 29000 32778 29052 32784
rect 28816 32428 28868 32434
rect 28816 32370 28868 32376
rect 29012 32298 29040 32778
rect 29104 32502 29132 33458
rect 29196 32978 29224 37810
rect 29552 36780 29604 36786
rect 29552 36722 29604 36728
rect 29276 36576 29328 36582
rect 29276 36518 29328 36524
rect 29288 35766 29316 36518
rect 29564 36378 29592 36722
rect 29552 36372 29604 36378
rect 29552 36314 29604 36320
rect 29748 36174 29776 38694
rect 30104 38276 30156 38282
rect 30104 38218 30156 38224
rect 29828 38004 29880 38010
rect 29828 37946 29880 37952
rect 29736 36168 29788 36174
rect 29736 36110 29788 36116
rect 29276 35760 29328 35766
rect 29276 35702 29328 35708
rect 29184 32972 29236 32978
rect 29184 32914 29236 32920
rect 29288 32842 29316 35702
rect 29644 34536 29696 34542
rect 29644 34478 29696 34484
rect 29368 33312 29420 33318
rect 29368 33254 29420 33260
rect 29276 32836 29328 32842
rect 29276 32778 29328 32784
rect 29092 32496 29144 32502
rect 29092 32438 29144 32444
rect 29000 32292 29052 32298
rect 29000 32234 29052 32240
rect 29012 32026 29040 32234
rect 29000 32020 29052 32026
rect 29000 31962 29052 31968
rect 28632 30252 28684 30258
rect 28632 30194 28684 30200
rect 28908 30252 28960 30258
rect 28908 30194 28960 30200
rect 28920 29850 28948 30194
rect 28908 29844 28960 29850
rect 28908 29786 28960 29792
rect 28540 29640 28592 29646
rect 28540 29582 28592 29588
rect 29012 29306 29040 31962
rect 29092 29708 29144 29714
rect 29092 29650 29144 29656
rect 29000 29300 29052 29306
rect 29000 29242 29052 29248
rect 29104 28762 29132 29650
rect 29092 28756 29144 28762
rect 29092 28698 29144 28704
rect 28448 28552 28500 28558
rect 28448 28494 28500 28500
rect 28448 27396 28500 27402
rect 28448 27338 28500 27344
rect 28460 23882 28488 27338
rect 28540 27328 28592 27334
rect 28540 27270 28592 27276
rect 28552 25906 28580 27270
rect 29380 27130 29408 33254
rect 29656 32434 29684 34478
rect 29748 32994 29776 36110
rect 29840 35562 29868 37946
rect 30116 37874 30144 38218
rect 30104 37868 30156 37874
rect 30104 37810 30156 37816
rect 30116 37466 30144 37810
rect 30104 37460 30156 37466
rect 30104 37402 30156 37408
rect 30104 37120 30156 37126
rect 30104 37062 30156 37068
rect 30116 36786 30144 37062
rect 30208 36922 30236 38898
rect 30288 37188 30340 37194
rect 30288 37130 30340 37136
rect 30196 36916 30248 36922
rect 30196 36858 30248 36864
rect 30300 36854 30328 37130
rect 30288 36848 30340 36854
rect 30288 36790 30340 36796
rect 30104 36780 30156 36786
rect 30104 36722 30156 36728
rect 29920 36100 29972 36106
rect 29920 36042 29972 36048
rect 29932 35698 29960 36042
rect 30116 35834 30144 36722
rect 30104 35828 30156 35834
rect 30104 35770 30156 35776
rect 29920 35692 29972 35698
rect 29920 35634 29972 35640
rect 30196 35692 30248 35698
rect 30196 35634 30248 35640
rect 29828 35556 29880 35562
rect 29828 35498 29880 35504
rect 29932 35018 29960 35634
rect 30104 35284 30156 35290
rect 30104 35226 30156 35232
rect 29920 35012 29972 35018
rect 29920 34954 29972 34960
rect 29932 33998 29960 34954
rect 30116 34678 30144 35226
rect 30104 34672 30156 34678
rect 30104 34614 30156 34620
rect 30208 34542 30236 35634
rect 30196 34536 30248 34542
rect 30196 34478 30248 34484
rect 29920 33992 29972 33998
rect 29920 33934 29972 33940
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 30012 33924 30064 33930
rect 30012 33866 30064 33872
rect 29748 32966 29960 32994
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 29748 32570 29776 32846
rect 29932 32722 29960 32966
rect 29840 32694 29960 32722
rect 29736 32564 29788 32570
rect 29736 32506 29788 32512
rect 29644 32428 29696 32434
rect 29644 32370 29696 32376
rect 29552 31476 29604 31482
rect 29552 31418 29604 31424
rect 29460 31136 29512 31142
rect 29460 31078 29512 31084
rect 29472 30394 29500 31078
rect 29564 30938 29592 31418
rect 29552 30932 29604 30938
rect 29552 30874 29604 30880
rect 29460 30388 29512 30394
rect 29460 30330 29512 30336
rect 29552 29504 29604 29510
rect 29552 29446 29604 29452
rect 29460 27872 29512 27878
rect 29460 27814 29512 27820
rect 29472 27674 29500 27814
rect 29460 27668 29512 27674
rect 29460 27610 29512 27616
rect 29368 27124 29420 27130
rect 29368 27066 29420 27072
rect 29564 27062 29592 29446
rect 29552 27056 29604 27062
rect 29552 26998 29604 27004
rect 29656 26994 29684 32370
rect 29748 29646 29776 32506
rect 29840 29646 29868 32694
rect 29920 32564 29972 32570
rect 29920 32506 29972 32512
rect 29932 31482 29960 32506
rect 30024 32026 30052 33866
rect 30116 33590 30144 33934
rect 30104 33584 30156 33590
rect 30104 33526 30156 33532
rect 30012 32020 30064 32026
rect 30012 31962 30064 31968
rect 29920 31476 29972 31482
rect 29920 31418 29972 31424
rect 29920 31340 29972 31346
rect 29920 31282 29972 31288
rect 29736 29640 29788 29646
rect 29736 29582 29788 29588
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 29748 29170 29776 29582
rect 29932 29578 29960 31282
rect 30024 30666 30052 31962
rect 30116 31210 30144 33526
rect 30208 33522 30236 34478
rect 30196 33516 30248 33522
rect 30196 33458 30248 33464
rect 30208 33046 30236 33458
rect 30196 33040 30248 33046
rect 30196 32982 30248 32988
rect 30196 32836 30248 32842
rect 30196 32778 30248 32784
rect 30208 32366 30236 32778
rect 30196 32360 30248 32366
rect 30196 32302 30248 32308
rect 30208 31346 30236 32302
rect 30300 32298 30328 36790
rect 30392 33454 30420 39238
rect 31128 38418 31156 39238
rect 31116 38412 31168 38418
rect 31116 38354 31168 38360
rect 30748 38344 30800 38350
rect 30748 38286 30800 38292
rect 30472 38208 30524 38214
rect 30472 38150 30524 38156
rect 30484 37942 30512 38150
rect 30472 37936 30524 37942
rect 30472 37878 30524 37884
rect 30564 36712 30616 36718
rect 30564 36654 30616 36660
rect 30576 36242 30604 36654
rect 30564 36236 30616 36242
rect 30564 36178 30616 36184
rect 30576 35834 30604 36178
rect 30656 36032 30708 36038
rect 30656 35974 30708 35980
rect 30564 35828 30616 35834
rect 30564 35770 30616 35776
rect 30472 35556 30524 35562
rect 30472 35498 30524 35504
rect 30484 35290 30512 35498
rect 30472 35284 30524 35290
rect 30472 35226 30524 35232
rect 30472 33856 30524 33862
rect 30472 33798 30524 33804
rect 30484 33522 30512 33798
rect 30576 33658 30604 35770
rect 30668 34610 30696 35974
rect 30656 34604 30708 34610
rect 30656 34546 30708 34552
rect 30760 33998 30788 38286
rect 31024 38276 31076 38282
rect 31024 38218 31076 38224
rect 31036 38010 31064 38218
rect 31024 38004 31076 38010
rect 31024 37946 31076 37952
rect 31128 37890 31156 38354
rect 31496 38350 31524 39238
rect 31484 38344 31536 38350
rect 31484 38286 31536 38292
rect 31392 38208 31444 38214
rect 31392 38150 31444 38156
rect 31036 37862 31156 37890
rect 31300 37868 31352 37874
rect 31036 37806 31064 37862
rect 31300 37810 31352 37816
rect 31024 37800 31076 37806
rect 31024 37742 31076 37748
rect 30932 35488 30984 35494
rect 30932 35430 30984 35436
rect 30944 35086 30972 35430
rect 30932 35080 30984 35086
rect 30932 35022 30984 35028
rect 30748 33992 30800 33998
rect 30748 33934 30800 33940
rect 30564 33652 30616 33658
rect 30564 33594 30616 33600
rect 30472 33516 30524 33522
rect 30472 33458 30524 33464
rect 30380 33448 30432 33454
rect 30380 33390 30432 33396
rect 30392 33318 30420 33390
rect 30380 33312 30432 33318
rect 30380 33254 30432 33260
rect 30288 32292 30340 32298
rect 30288 32234 30340 32240
rect 30196 31340 30248 31346
rect 30196 31282 30248 31288
rect 30380 31340 30432 31346
rect 30380 31282 30432 31288
rect 30104 31204 30156 31210
rect 30104 31146 30156 31152
rect 30392 30734 30420 31282
rect 30380 30728 30432 30734
rect 30380 30670 30432 30676
rect 30012 30660 30064 30666
rect 30012 30602 30064 30608
rect 30196 30592 30248 30598
rect 30196 30534 30248 30540
rect 30012 30184 30064 30190
rect 30012 30126 30064 30132
rect 29920 29572 29972 29578
rect 29920 29514 29972 29520
rect 29736 29164 29788 29170
rect 29736 29106 29788 29112
rect 29748 28082 29776 29106
rect 29736 28076 29788 28082
rect 29736 28018 29788 28024
rect 29748 27538 29776 28018
rect 30024 27878 30052 30126
rect 30104 29300 30156 29306
rect 30104 29242 30156 29248
rect 30012 27872 30064 27878
rect 30012 27814 30064 27820
rect 29736 27532 29788 27538
rect 29736 27474 29788 27480
rect 29644 26988 29696 26994
rect 29644 26930 29696 26936
rect 29276 26784 29328 26790
rect 29276 26726 29328 26732
rect 29288 26314 29316 26726
rect 29656 26586 29684 26930
rect 30116 26586 30144 29242
rect 29460 26580 29512 26586
rect 29460 26522 29512 26528
rect 29644 26580 29696 26586
rect 29644 26522 29696 26528
rect 30104 26580 30156 26586
rect 30104 26522 30156 26528
rect 29276 26308 29328 26314
rect 29276 26250 29328 26256
rect 28540 25900 28592 25906
rect 28540 25842 28592 25848
rect 28632 25900 28684 25906
rect 28632 25842 28684 25848
rect 28552 24018 28580 25842
rect 28644 24274 28672 25842
rect 29000 24880 29052 24886
rect 29000 24822 29052 24828
rect 28816 24608 28868 24614
rect 28816 24550 28868 24556
rect 28908 24608 28960 24614
rect 28908 24550 28960 24556
rect 28632 24268 28684 24274
rect 28632 24210 28684 24216
rect 28644 24138 28672 24210
rect 28828 24206 28856 24550
rect 28816 24200 28868 24206
rect 28816 24142 28868 24148
rect 28632 24132 28684 24138
rect 28632 24074 28684 24080
rect 28552 23990 28672 24018
rect 28460 23854 28580 23882
rect 28368 22066 28488 22094
rect 28080 21548 28132 21554
rect 28080 21490 28132 21496
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 27908 20262 27936 20402
rect 27896 20256 27948 20262
rect 27896 20198 27948 20204
rect 27908 19718 27936 20198
rect 27896 19712 27948 19718
rect 27896 19654 27948 19660
rect 27804 16992 27856 16998
rect 27804 16934 27856 16940
rect 27816 16658 27844 16934
rect 27804 16652 27856 16658
rect 27804 16594 27856 16600
rect 27620 15156 27672 15162
rect 27620 15098 27672 15104
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27528 14408 27580 14414
rect 27528 14350 27580 14356
rect 27540 14074 27568 14350
rect 27632 14074 27660 14962
rect 27712 14816 27764 14822
rect 27712 14758 27764 14764
rect 27528 14068 27580 14074
rect 27528 14010 27580 14016
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27724 13326 27752 14758
rect 27804 14340 27856 14346
rect 27804 14282 27856 14288
rect 27816 13394 27844 14282
rect 27804 13388 27856 13394
rect 27804 13330 27856 13336
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27908 12442 27936 19654
rect 28184 17218 28212 22066
rect 28460 21554 28488 22066
rect 28264 21548 28316 21554
rect 28264 21490 28316 21496
rect 28448 21548 28500 21554
rect 28448 21490 28500 21496
rect 28276 20262 28304 21490
rect 28460 20806 28488 21490
rect 28448 20800 28500 20806
rect 28448 20742 28500 20748
rect 28264 20256 28316 20262
rect 28264 20198 28316 20204
rect 28356 19304 28408 19310
rect 28356 19246 28408 19252
rect 28368 18970 28396 19246
rect 28356 18964 28408 18970
rect 28356 18906 28408 18912
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28264 17604 28316 17610
rect 28264 17546 28316 17552
rect 28092 17190 28212 17218
rect 27896 12436 27948 12442
rect 27448 12406 27568 12434
rect 27436 12096 27488 12102
rect 27436 12038 27488 12044
rect 27448 11762 27476 12038
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27068 10532 27120 10538
rect 27068 10474 27120 10480
rect 27436 8492 27488 8498
rect 27436 8434 27488 8440
rect 26792 8356 26844 8362
rect 26792 8298 26844 8304
rect 27448 8090 27476 8434
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 27344 7404 27396 7410
rect 27344 7346 27396 7352
rect 27252 7336 27304 7342
rect 27252 7278 27304 7284
rect 26976 6996 27028 7002
rect 26976 6938 27028 6944
rect 26988 6322 27016 6938
rect 27264 6934 27292 7278
rect 27252 6928 27304 6934
rect 27252 6870 27304 6876
rect 27068 6860 27120 6866
rect 27068 6802 27120 6808
rect 26976 6316 27028 6322
rect 26976 6258 27028 6264
rect 27080 5642 27108 6802
rect 27356 6730 27384 7346
rect 27540 6905 27568 12406
rect 27896 12378 27948 12384
rect 27908 11898 27936 12378
rect 28092 12238 28120 17190
rect 28172 17060 28224 17066
rect 28172 17002 28224 17008
rect 28184 16590 28212 17002
rect 28172 16584 28224 16590
rect 28172 16526 28224 16532
rect 28276 15162 28304 17546
rect 28368 16794 28396 17614
rect 28356 16788 28408 16794
rect 28356 16730 28408 16736
rect 28368 16590 28396 16730
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 28264 15156 28316 15162
rect 28264 15098 28316 15104
rect 28276 14414 28304 15098
rect 28264 14408 28316 14414
rect 28264 14350 28316 14356
rect 28276 13394 28304 14350
rect 28264 13388 28316 13394
rect 28264 13330 28316 13336
rect 28080 12232 28132 12238
rect 28080 12174 28132 12180
rect 28172 12164 28224 12170
rect 28172 12106 28224 12112
rect 27896 11892 27948 11898
rect 27896 11834 27948 11840
rect 27908 11626 27936 11834
rect 28184 11830 28212 12106
rect 28172 11824 28224 11830
rect 28172 11766 28224 11772
rect 27896 11620 27948 11626
rect 27896 11562 27948 11568
rect 28460 11150 28488 20742
rect 28552 18426 28580 23854
rect 28644 20466 28672 23990
rect 28920 23798 28948 24550
rect 29012 24256 29040 24822
rect 29092 24268 29144 24274
rect 29012 24228 29092 24256
rect 28908 23792 28960 23798
rect 28908 23734 28960 23740
rect 28816 23044 28868 23050
rect 28816 22986 28868 22992
rect 28828 21690 28856 22986
rect 28908 22568 28960 22574
rect 28908 22510 28960 22516
rect 28920 22234 28948 22510
rect 28908 22228 28960 22234
rect 28908 22170 28960 22176
rect 28816 21684 28868 21690
rect 28816 21626 28868 21632
rect 29012 21486 29040 24228
rect 29092 24210 29144 24216
rect 29288 22030 29316 26250
rect 29276 22024 29328 22030
rect 29276 21966 29328 21972
rect 29000 21480 29052 21486
rect 29000 21422 29052 21428
rect 29184 21004 29236 21010
rect 29184 20946 29236 20952
rect 29196 20874 29224 20946
rect 29184 20868 29236 20874
rect 29184 20810 29236 20816
rect 29000 20800 29052 20806
rect 29000 20742 29052 20748
rect 28632 20460 28684 20466
rect 28632 20402 28684 20408
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28828 19378 28856 19790
rect 28816 19372 28868 19378
rect 28816 19314 28868 19320
rect 28540 18420 28592 18426
rect 28540 18362 28592 18368
rect 28540 18216 28592 18222
rect 28540 18158 28592 18164
rect 28448 11144 28500 11150
rect 28448 11086 28500 11092
rect 27988 10464 28040 10470
rect 27988 10406 28040 10412
rect 28000 10062 28028 10406
rect 28552 10266 28580 18158
rect 28632 16992 28684 16998
rect 28632 16934 28684 16940
rect 28644 16590 28672 16934
rect 28632 16584 28684 16590
rect 28632 16526 28684 16532
rect 28632 11076 28684 11082
rect 28632 11018 28684 11024
rect 28540 10260 28592 10266
rect 28540 10202 28592 10208
rect 28644 10130 28672 11018
rect 28632 10124 28684 10130
rect 28632 10066 28684 10072
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 28540 10056 28592 10062
rect 28540 9998 28592 10004
rect 27526 6896 27582 6905
rect 27526 6831 27582 6840
rect 27540 6798 27568 6831
rect 27528 6792 27580 6798
rect 27448 6752 27528 6780
rect 27344 6724 27396 6730
rect 27344 6666 27396 6672
rect 27448 6458 27476 6752
rect 27528 6734 27580 6740
rect 27528 6656 27580 6662
rect 27528 6598 27580 6604
rect 27436 6452 27488 6458
rect 27436 6394 27488 6400
rect 27540 6322 27568 6598
rect 27528 6316 27580 6322
rect 27528 6258 27580 6264
rect 27540 5710 27568 6258
rect 27724 5846 27752 9998
rect 28448 9988 28500 9994
rect 28448 9930 28500 9936
rect 28172 9648 28224 9654
rect 28172 9590 28224 9596
rect 28184 8906 28212 9590
rect 28356 8968 28408 8974
rect 28356 8910 28408 8916
rect 28172 8900 28224 8906
rect 28172 8842 28224 8848
rect 28184 8430 28212 8842
rect 28172 8424 28224 8430
rect 28172 8366 28224 8372
rect 28184 7818 28212 8366
rect 28172 7812 28224 7818
rect 28172 7754 28224 7760
rect 28368 7546 28396 8910
rect 28460 8838 28488 9930
rect 28552 9518 28580 9998
rect 28540 9512 28592 9518
rect 28540 9454 28592 9460
rect 28552 9110 28580 9454
rect 28724 9444 28776 9450
rect 28724 9386 28776 9392
rect 28540 9104 28592 9110
rect 28540 9046 28592 9052
rect 28448 8832 28500 8838
rect 28448 8774 28500 8780
rect 28460 8498 28488 8774
rect 28448 8492 28500 8498
rect 28448 8434 28500 8440
rect 28552 8430 28580 9046
rect 28736 8974 28764 9386
rect 28724 8968 28776 8974
rect 28724 8910 28776 8916
rect 28540 8424 28592 8430
rect 28540 8366 28592 8372
rect 28736 7954 28764 8910
rect 29012 8090 29040 20742
rect 29092 13524 29144 13530
rect 29092 13466 29144 13472
rect 29104 11286 29132 13466
rect 29092 11280 29144 11286
rect 29092 11222 29144 11228
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 29000 8084 29052 8090
rect 29000 8026 29052 8032
rect 28724 7948 28776 7954
rect 28724 7890 28776 7896
rect 28448 7880 28500 7886
rect 28448 7822 28500 7828
rect 28356 7540 28408 7546
rect 28356 7482 28408 7488
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 28184 6186 28212 6734
rect 28368 6730 28396 7482
rect 28356 6724 28408 6730
rect 28356 6666 28408 6672
rect 28172 6180 28224 6186
rect 28172 6122 28224 6128
rect 27712 5840 27764 5846
rect 27712 5782 27764 5788
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 27068 5636 27120 5642
rect 27068 5578 27120 5584
rect 27080 4690 27108 5578
rect 27344 5024 27396 5030
rect 27344 4966 27396 4972
rect 27068 4684 27120 4690
rect 27068 4626 27120 4632
rect 27356 4622 27384 4966
rect 27540 4622 27568 5646
rect 27988 5296 28040 5302
rect 27988 5238 28040 5244
rect 27344 4616 27396 4622
rect 27344 4558 27396 4564
rect 27528 4616 27580 4622
rect 27528 4558 27580 4564
rect 26884 4480 26936 4486
rect 26884 4422 26936 4428
rect 26896 3534 26924 4422
rect 28000 3738 28028 5238
rect 28184 5234 28212 6122
rect 28460 5302 28488 7822
rect 28724 6656 28776 6662
rect 28724 6598 28776 6604
rect 28736 6254 28764 6598
rect 29104 6458 29132 11086
rect 29092 6452 29144 6458
rect 29092 6394 29144 6400
rect 29104 6254 29132 6394
rect 28724 6248 28776 6254
rect 28724 6190 28776 6196
rect 28816 6248 28868 6254
rect 28816 6190 28868 6196
rect 29092 6248 29144 6254
rect 29092 6190 29144 6196
rect 28448 5296 28500 5302
rect 28448 5238 28500 5244
rect 28172 5228 28224 5234
rect 28172 5170 28224 5176
rect 27988 3732 28040 3738
rect 27988 3674 28040 3680
rect 26884 3528 26936 3534
rect 26884 3470 26936 3476
rect 28632 3528 28684 3534
rect 28632 3470 28684 3476
rect 26976 2848 27028 2854
rect 26976 2790 27028 2796
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 28080 2848 28132 2854
rect 28080 2790 28132 2796
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 26700 2372 26752 2378
rect 26700 2314 26752 2320
rect 26712 800 26740 2314
rect 26988 800 27016 2790
rect 27252 2576 27304 2582
rect 27252 2518 27304 2524
rect 27264 800 27292 2518
rect 27528 2440 27580 2446
rect 27528 2382 27580 2388
rect 27540 800 27568 2382
rect 27816 800 27844 2790
rect 28092 800 28120 2790
rect 28356 2576 28408 2582
rect 28356 2518 28408 2524
rect 28368 800 28396 2518
rect 28644 800 28672 3470
rect 28828 1970 28856 6190
rect 29196 5914 29224 20810
rect 29368 20460 29420 20466
rect 29368 20402 29420 20408
rect 29380 19310 29408 20402
rect 29368 19304 29420 19310
rect 29368 19246 29420 19252
rect 29276 18624 29328 18630
rect 29276 18566 29328 18572
rect 29288 10266 29316 18566
rect 29472 17134 29500 26522
rect 30116 26042 30144 26522
rect 30104 26036 30156 26042
rect 30104 25978 30156 25984
rect 29828 25424 29880 25430
rect 29828 25366 29880 25372
rect 29840 25294 29868 25366
rect 29828 25288 29880 25294
rect 29828 25230 29880 25236
rect 29736 25220 29788 25226
rect 29736 25162 29788 25168
rect 29644 25152 29696 25158
rect 29644 25094 29696 25100
rect 29656 23730 29684 25094
rect 29748 24886 29776 25162
rect 30012 25152 30064 25158
rect 30012 25094 30064 25100
rect 29736 24880 29788 24886
rect 29736 24822 29788 24828
rect 30024 24410 30052 25094
rect 30104 24812 30156 24818
rect 30104 24754 30156 24760
rect 30116 24410 30144 24754
rect 30012 24404 30064 24410
rect 30012 24346 30064 24352
rect 30104 24404 30156 24410
rect 30104 24346 30156 24352
rect 29920 24064 29972 24070
rect 29920 24006 29972 24012
rect 29644 23724 29696 23730
rect 29644 23666 29696 23672
rect 29932 23322 29960 24006
rect 30012 23588 30064 23594
rect 30012 23530 30064 23536
rect 29644 23316 29696 23322
rect 29644 23258 29696 23264
rect 29920 23316 29972 23322
rect 29920 23258 29972 23264
rect 29656 21690 29684 23258
rect 29920 22094 29972 22098
rect 30024 22094 30052 23530
rect 29920 22092 30052 22094
rect 29972 22066 30052 22092
rect 29920 22034 29972 22040
rect 29644 21684 29696 21690
rect 29644 21626 29696 21632
rect 29656 21486 29684 21626
rect 29644 21480 29696 21486
rect 29644 21422 29696 21428
rect 29828 21480 29880 21486
rect 29828 21422 29880 21428
rect 29736 21344 29788 21350
rect 29736 21286 29788 21292
rect 29748 20602 29776 21286
rect 29840 20806 29868 21422
rect 29828 20800 29880 20806
rect 29828 20742 29880 20748
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 29736 20596 29788 20602
rect 29736 20538 29788 20544
rect 29552 20460 29604 20466
rect 29552 20402 29604 20408
rect 29564 19854 29592 20402
rect 29920 19916 29972 19922
rect 29920 19858 29972 19864
rect 29552 19848 29604 19854
rect 29552 19790 29604 19796
rect 29736 19304 29788 19310
rect 29736 19246 29788 19252
rect 29552 19236 29604 19242
rect 29552 19178 29604 19184
rect 29460 17128 29512 17134
rect 29460 17070 29512 17076
rect 29564 15706 29592 19178
rect 29748 18766 29776 19246
rect 29932 18766 29960 19858
rect 29736 18760 29788 18766
rect 29736 18702 29788 18708
rect 29920 18760 29972 18766
rect 29920 18702 29972 18708
rect 29828 18692 29880 18698
rect 29828 18634 29880 18640
rect 29840 16454 29868 18634
rect 29828 16448 29880 16454
rect 29828 16390 29880 16396
rect 29840 16114 29868 16390
rect 29828 16108 29880 16114
rect 29828 16050 29880 16056
rect 29920 16040 29972 16046
rect 29920 15982 29972 15988
rect 29828 15972 29880 15978
rect 29828 15914 29880 15920
rect 29552 15700 29604 15706
rect 29552 15642 29604 15648
rect 29368 14408 29420 14414
rect 29368 14350 29420 14356
rect 29380 12918 29408 14350
rect 29564 14346 29592 15642
rect 29644 15020 29696 15026
rect 29644 14962 29696 14968
rect 29656 14822 29684 14962
rect 29840 14958 29868 15914
rect 29932 14958 29960 15982
rect 29828 14952 29880 14958
rect 29828 14894 29880 14900
rect 29920 14952 29972 14958
rect 29920 14894 29972 14900
rect 29644 14816 29696 14822
rect 29644 14758 29696 14764
rect 29552 14340 29604 14346
rect 29552 14282 29604 14288
rect 29552 13796 29604 13802
rect 29552 13738 29604 13744
rect 29564 12918 29592 13738
rect 29368 12912 29420 12918
rect 29368 12854 29420 12860
rect 29552 12912 29604 12918
rect 29552 12854 29604 12860
rect 29368 11280 29420 11286
rect 29368 11222 29420 11228
rect 29276 10260 29328 10266
rect 29276 10202 29328 10208
rect 29288 10062 29316 10202
rect 29276 10056 29328 10062
rect 29276 9998 29328 10004
rect 29380 6361 29408 11222
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29564 9654 29592 10406
rect 29552 9648 29604 9654
rect 29552 9590 29604 9596
rect 29656 8022 29684 14758
rect 29840 14414 29868 14894
rect 29828 14408 29880 14414
rect 29828 14350 29880 14356
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29748 12986 29776 13262
rect 29932 13190 29960 14894
rect 30012 13524 30064 13530
rect 30012 13466 30064 13472
rect 30024 13326 30052 13466
rect 30012 13320 30064 13326
rect 30012 13262 30064 13268
rect 29920 13184 29972 13190
rect 29920 13126 29972 13132
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 30116 12306 30144 20742
rect 30208 18358 30236 30534
rect 30576 30258 30604 33594
rect 30656 32768 30708 32774
rect 30656 32710 30708 32716
rect 30668 30326 30696 32710
rect 30760 32026 30788 33934
rect 30840 33312 30892 33318
rect 30840 33254 30892 33260
rect 30748 32020 30800 32026
rect 30748 31962 30800 31968
rect 30852 31822 30880 33254
rect 31036 32910 31064 37742
rect 31312 37466 31340 37810
rect 31300 37460 31352 37466
rect 31300 37402 31352 37408
rect 31312 36786 31340 37402
rect 31300 36780 31352 36786
rect 31300 36722 31352 36728
rect 31116 34944 31168 34950
rect 31116 34886 31168 34892
rect 31024 32904 31076 32910
rect 31024 32846 31076 32852
rect 30932 32768 30984 32774
rect 30932 32710 30984 32716
rect 30840 31816 30892 31822
rect 30840 31758 30892 31764
rect 30944 31414 30972 32710
rect 31128 31414 31156 34886
rect 31300 32836 31352 32842
rect 31300 32778 31352 32784
rect 31208 32224 31260 32230
rect 31208 32166 31260 32172
rect 31220 32026 31248 32166
rect 31208 32020 31260 32026
rect 31208 31962 31260 31968
rect 30932 31408 30984 31414
rect 30932 31350 30984 31356
rect 31116 31408 31168 31414
rect 31116 31350 31168 31356
rect 30944 30938 30972 31350
rect 31208 31340 31260 31346
rect 31208 31282 31260 31288
rect 31024 31136 31076 31142
rect 31024 31078 31076 31084
rect 31116 31136 31168 31142
rect 31116 31078 31168 31084
rect 30932 30932 30984 30938
rect 30932 30874 30984 30880
rect 30840 30388 30892 30394
rect 30840 30330 30892 30336
rect 30656 30320 30708 30326
rect 30656 30262 30708 30268
rect 30288 30252 30340 30258
rect 30288 30194 30340 30200
rect 30564 30252 30616 30258
rect 30564 30194 30616 30200
rect 30300 29034 30328 30194
rect 30748 29640 30800 29646
rect 30748 29582 30800 29588
rect 30380 29572 30432 29578
rect 30380 29514 30432 29520
rect 30288 29028 30340 29034
rect 30288 28970 30340 28976
rect 30392 28626 30420 29514
rect 30380 28620 30432 28626
rect 30380 28562 30432 28568
rect 30760 28082 30788 29582
rect 30852 29102 30880 30330
rect 30840 29096 30892 29102
rect 30840 29038 30892 29044
rect 30852 28762 30880 29038
rect 30840 28756 30892 28762
rect 30840 28698 30892 28704
rect 30748 28076 30800 28082
rect 30748 28018 30800 28024
rect 30288 27872 30340 27878
rect 30288 27814 30340 27820
rect 30300 26926 30328 27814
rect 30932 27464 30984 27470
rect 30932 27406 30984 27412
rect 30944 27130 30972 27406
rect 30932 27124 30984 27130
rect 30932 27066 30984 27072
rect 30288 26920 30340 26926
rect 30288 26862 30340 26868
rect 30748 25696 30800 25702
rect 30748 25638 30800 25644
rect 30380 25424 30432 25430
rect 30380 25366 30432 25372
rect 30392 20806 30420 25366
rect 30656 25288 30708 25294
rect 30656 25230 30708 25236
rect 30668 24818 30696 25230
rect 30760 24818 30788 25638
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 30748 24812 30800 24818
rect 30748 24754 30800 24760
rect 30668 24342 30696 24754
rect 30656 24336 30708 24342
rect 30656 24278 30708 24284
rect 30656 23792 30708 23798
rect 30656 23734 30708 23740
rect 30380 20800 30432 20806
rect 30380 20742 30432 20748
rect 30668 20534 30696 23734
rect 30656 20528 30708 20534
rect 30656 20470 30708 20476
rect 30472 20392 30524 20398
rect 30472 20334 30524 20340
rect 30380 20256 30432 20262
rect 30380 20198 30432 20204
rect 30392 19514 30420 20198
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30196 18352 30248 18358
rect 30196 18294 30248 18300
rect 30380 17128 30432 17134
rect 30380 17070 30432 17076
rect 30392 16522 30420 17070
rect 30380 16516 30432 16522
rect 30380 16458 30432 16464
rect 30392 16114 30420 16458
rect 30380 16108 30432 16114
rect 30380 16050 30432 16056
rect 30380 15904 30432 15910
rect 30380 15846 30432 15852
rect 30392 15026 30420 15846
rect 30380 15020 30432 15026
rect 30380 14962 30432 14968
rect 30380 13932 30432 13938
rect 30380 13874 30432 13880
rect 30392 13530 30420 13874
rect 30380 13524 30432 13530
rect 30380 13466 30432 13472
rect 30104 12300 30156 12306
rect 30104 12242 30156 12248
rect 30196 12096 30248 12102
rect 30196 12038 30248 12044
rect 30208 11694 30236 12038
rect 30288 11756 30340 11762
rect 30288 11698 30340 11704
rect 30196 11688 30248 11694
rect 30196 11630 30248 11636
rect 30208 10656 30236 11630
rect 30300 11354 30328 11698
rect 30288 11348 30340 11354
rect 30288 11290 30340 11296
rect 30288 10668 30340 10674
rect 30208 10628 30288 10656
rect 30288 10610 30340 10616
rect 29920 10464 29972 10470
rect 29920 10406 29972 10412
rect 29736 9580 29788 9586
rect 29736 9522 29788 9528
rect 29748 8906 29776 9522
rect 29932 9518 29960 10406
rect 30012 10056 30064 10062
rect 30012 9998 30064 10004
rect 30024 9722 30052 9998
rect 30012 9716 30064 9722
rect 30012 9658 30064 9664
rect 30300 9654 30328 10610
rect 30380 10532 30432 10538
rect 30380 10474 30432 10480
rect 30392 10198 30420 10474
rect 30380 10192 30432 10198
rect 30380 10134 30432 10140
rect 30288 9648 30340 9654
rect 30288 9590 30340 9596
rect 29920 9512 29972 9518
rect 29920 9454 29972 9460
rect 29932 8906 29960 9454
rect 29736 8900 29788 8906
rect 29736 8842 29788 8848
rect 29920 8900 29972 8906
rect 29920 8842 29972 8848
rect 29748 8634 29776 8842
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 29644 8016 29696 8022
rect 29644 7958 29696 7964
rect 29656 7478 29684 7958
rect 29644 7472 29696 7478
rect 29644 7414 29696 7420
rect 29644 7200 29696 7206
rect 29644 7142 29696 7148
rect 29366 6352 29422 6361
rect 29656 6322 29684 7142
rect 29366 6287 29422 6296
rect 29552 6316 29604 6322
rect 29380 6118 29408 6287
rect 29552 6258 29604 6264
rect 29644 6316 29696 6322
rect 29644 6258 29696 6264
rect 29368 6112 29420 6118
rect 29368 6054 29420 6060
rect 29184 5908 29236 5914
rect 29236 5868 29316 5896
rect 29184 5850 29236 5856
rect 29000 5568 29052 5574
rect 29000 5510 29052 5516
rect 29012 5302 29040 5510
rect 29000 5296 29052 5302
rect 29000 5238 29052 5244
rect 29184 2848 29236 2854
rect 29184 2790 29236 2796
rect 28908 2440 28960 2446
rect 28908 2382 28960 2388
rect 28816 1964 28868 1970
rect 28816 1906 28868 1912
rect 28920 800 28948 2382
rect 29196 800 29224 2790
rect 29288 2650 29316 5868
rect 29564 5710 29592 6258
rect 29828 6180 29880 6186
rect 29828 6122 29880 6128
rect 29552 5704 29604 5710
rect 29552 5646 29604 5652
rect 29840 5642 29868 6122
rect 29828 5636 29880 5642
rect 29828 5578 29880 5584
rect 29932 5302 29960 8842
rect 30300 7750 30328 9590
rect 30484 9178 30512 20334
rect 30840 19916 30892 19922
rect 30840 19858 30892 19864
rect 30852 19378 30880 19858
rect 30840 19372 30892 19378
rect 30840 19314 30892 19320
rect 30748 19304 30800 19310
rect 30800 19252 30880 19258
rect 30748 19246 30880 19252
rect 30760 19230 30880 19246
rect 30852 19174 30880 19230
rect 30748 19168 30800 19174
rect 30748 19110 30800 19116
rect 30840 19168 30892 19174
rect 30840 19110 30892 19116
rect 30562 18728 30618 18737
rect 30562 18663 30618 18672
rect 30576 18630 30604 18663
rect 30564 18624 30616 18630
rect 30564 18566 30616 18572
rect 30760 18086 30788 19110
rect 30930 18864 30986 18873
rect 30930 18799 30932 18808
rect 30984 18799 30986 18808
rect 30932 18770 30984 18776
rect 31036 18766 31064 31078
rect 31128 30734 31156 31078
rect 31116 30728 31168 30734
rect 31116 30670 31168 30676
rect 31220 30598 31248 31282
rect 31312 30802 31340 32778
rect 31404 31346 31432 38150
rect 31588 37874 31616 39374
rect 31576 37868 31628 37874
rect 31576 37810 31628 37816
rect 31576 36712 31628 36718
rect 31576 36654 31628 36660
rect 31588 36038 31616 36654
rect 31576 36032 31628 36038
rect 31576 35974 31628 35980
rect 31484 32904 31536 32910
rect 31484 32846 31536 32852
rect 31496 32774 31524 32846
rect 31484 32768 31536 32774
rect 31484 32710 31536 32716
rect 31392 31340 31444 31346
rect 31392 31282 31444 31288
rect 31300 30796 31352 30802
rect 31300 30738 31352 30744
rect 31208 30592 31260 30598
rect 31208 30534 31260 30540
rect 31220 30394 31248 30534
rect 31208 30388 31260 30394
rect 31208 30330 31260 30336
rect 31312 29850 31340 30738
rect 31576 30728 31628 30734
rect 31576 30670 31628 30676
rect 31588 30122 31616 30670
rect 31576 30116 31628 30122
rect 31576 30058 31628 30064
rect 31300 29844 31352 29850
rect 31300 29786 31352 29792
rect 31576 28552 31628 28558
rect 31576 28494 31628 28500
rect 31588 28014 31616 28494
rect 31576 28008 31628 28014
rect 31576 27950 31628 27956
rect 31576 26036 31628 26042
rect 31576 25978 31628 25984
rect 31300 25832 31352 25838
rect 31300 25774 31352 25780
rect 31208 25764 31260 25770
rect 31208 25706 31260 25712
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 31024 18760 31076 18766
rect 31024 18702 31076 18708
rect 30748 18080 30800 18086
rect 30748 18022 30800 18028
rect 30564 16516 30616 16522
rect 30564 16458 30616 16464
rect 30576 15162 30604 16458
rect 30656 16040 30708 16046
rect 30656 15982 30708 15988
rect 30668 15706 30696 15982
rect 30656 15700 30708 15706
rect 30656 15642 30708 15648
rect 30564 15156 30616 15162
rect 30564 15098 30616 15104
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 30576 13394 30604 14962
rect 30852 14634 30880 18702
rect 30932 17196 30984 17202
rect 30932 17138 30984 17144
rect 30944 16590 30972 17138
rect 30932 16584 30984 16590
rect 30932 16526 30984 16532
rect 30944 16046 30972 16526
rect 30932 16040 30984 16046
rect 30932 15982 30984 15988
rect 30944 15638 30972 15982
rect 30932 15632 30984 15638
rect 30932 15574 30984 15580
rect 30760 14606 30880 14634
rect 30564 13388 30616 13394
rect 30564 13330 30616 13336
rect 30656 13320 30708 13326
rect 30656 13262 30708 13268
rect 30668 12986 30696 13262
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30760 12434 30788 14606
rect 30944 13938 30972 15574
rect 31024 15496 31076 15502
rect 31024 15438 31076 15444
rect 31036 14822 31064 15438
rect 31024 14816 31076 14822
rect 31024 14758 31076 14764
rect 30932 13932 30984 13938
rect 30932 13874 30984 13880
rect 30840 12980 30892 12986
rect 30840 12922 30892 12928
rect 30668 12406 30788 12434
rect 30564 12232 30616 12238
rect 30564 12174 30616 12180
rect 30576 11762 30604 12174
rect 30564 11756 30616 11762
rect 30564 11698 30616 11704
rect 30668 10010 30696 12406
rect 30748 12232 30800 12238
rect 30748 12174 30800 12180
rect 30760 11898 30788 12174
rect 30748 11892 30800 11898
rect 30748 11834 30800 11840
rect 30576 9982 30696 10010
rect 30472 9172 30524 9178
rect 30472 9114 30524 9120
rect 30576 8566 30604 9982
rect 30656 9920 30708 9926
rect 30656 9862 30708 9868
rect 30668 8566 30696 9862
rect 30564 8560 30616 8566
rect 30564 8502 30616 8508
rect 30656 8560 30708 8566
rect 30656 8502 30708 8508
rect 30288 7744 30340 7750
rect 30288 7686 30340 7692
rect 30196 6724 30248 6730
rect 30196 6666 30248 6672
rect 30208 6458 30236 6666
rect 30012 6452 30064 6458
rect 30012 6394 30064 6400
rect 30196 6452 30248 6458
rect 30196 6394 30248 6400
rect 30024 6322 30052 6394
rect 30012 6316 30064 6322
rect 30012 6258 30064 6264
rect 30196 6112 30248 6118
rect 30196 6054 30248 6060
rect 30208 5778 30236 6054
rect 30564 5908 30616 5914
rect 30564 5850 30616 5856
rect 30196 5772 30248 5778
rect 30196 5714 30248 5720
rect 30576 5710 30604 5850
rect 30564 5704 30616 5710
rect 30564 5646 30616 5652
rect 30288 5568 30340 5574
rect 30288 5510 30340 5516
rect 29920 5296 29972 5302
rect 29920 5238 29972 5244
rect 30300 4622 30328 5510
rect 30852 4622 30880 12922
rect 31036 12306 31064 14758
rect 31220 13326 31248 25706
rect 31312 25498 31340 25774
rect 31300 25492 31352 25498
rect 31300 25434 31352 25440
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31404 22098 31432 22578
rect 31392 22092 31444 22098
rect 31392 22034 31444 22040
rect 31404 19922 31432 22034
rect 31392 19916 31444 19922
rect 31392 19858 31444 19864
rect 31300 19372 31352 19378
rect 31300 19314 31352 19320
rect 31312 18902 31340 19314
rect 31300 18896 31352 18902
rect 31300 18838 31352 18844
rect 31392 17672 31444 17678
rect 31392 17614 31444 17620
rect 31404 16250 31432 17614
rect 31588 17270 31616 25978
rect 31576 17264 31628 17270
rect 31576 17206 31628 17212
rect 31484 16516 31536 16522
rect 31484 16458 31536 16464
rect 31496 16250 31524 16458
rect 31392 16244 31444 16250
rect 31392 16186 31444 16192
rect 31484 16244 31536 16250
rect 31484 16186 31536 16192
rect 31404 16114 31432 16186
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31484 15428 31536 15434
rect 31484 15370 31536 15376
rect 31496 14618 31524 15370
rect 31484 14612 31536 14618
rect 31484 14554 31536 14560
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 31680 12434 31708 56306
rect 32140 50289 32168 56306
rect 32126 50280 32182 50289
rect 32126 50215 32182 50224
rect 33980 47598 34008 56306
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 33968 47592 34020 47598
rect 33968 47534 34020 47540
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 32220 40520 32272 40526
rect 32220 40462 32272 40468
rect 32036 40384 32088 40390
rect 32036 40326 32088 40332
rect 32048 39370 32076 40326
rect 32036 39364 32088 39370
rect 32036 39306 32088 39312
rect 32048 37856 32076 39306
rect 32232 38418 32260 40462
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 32220 38412 32272 38418
rect 32220 38354 32272 38360
rect 32680 38412 32732 38418
rect 32680 38354 32732 38360
rect 31956 37828 32076 37856
rect 32588 37868 32640 37874
rect 31760 34604 31812 34610
rect 31760 34546 31812 34552
rect 31772 33998 31800 34546
rect 31760 33992 31812 33998
rect 31760 33934 31812 33940
rect 31772 32434 31800 33934
rect 31852 33448 31904 33454
rect 31852 33390 31904 33396
rect 31864 32842 31892 33390
rect 31852 32836 31904 32842
rect 31852 32778 31904 32784
rect 31760 32428 31812 32434
rect 31760 32370 31812 32376
rect 31956 31142 31984 37828
rect 32588 37810 32640 37816
rect 32600 36922 32628 37810
rect 32692 37466 32720 38354
rect 33048 38276 33100 38282
rect 33048 38218 33100 38224
rect 33060 38010 33088 38218
rect 33876 38208 33928 38214
rect 33876 38150 33928 38156
rect 33048 38004 33100 38010
rect 33048 37946 33100 37952
rect 32680 37460 32732 37466
rect 32680 37402 32732 37408
rect 32588 36916 32640 36922
rect 32588 36858 32640 36864
rect 32692 35154 32720 37402
rect 33888 36854 33916 38150
rect 34612 38004 34664 38010
rect 34612 37946 34664 37952
rect 34244 37868 34296 37874
rect 34244 37810 34296 37816
rect 34520 37868 34572 37874
rect 34520 37810 34572 37816
rect 34152 37664 34204 37670
rect 34152 37606 34204 37612
rect 33876 36848 33928 36854
rect 33230 36816 33286 36825
rect 33230 36751 33232 36760
rect 33284 36751 33286 36760
rect 33782 36816 33838 36825
rect 33876 36790 33928 36796
rect 34060 36848 34112 36854
rect 34060 36790 34112 36796
rect 33782 36751 33838 36760
rect 33232 36722 33284 36728
rect 33600 36712 33652 36718
rect 33600 36654 33652 36660
rect 33612 36174 33640 36654
rect 33692 36576 33744 36582
rect 33692 36518 33744 36524
rect 33600 36168 33652 36174
rect 33600 36110 33652 36116
rect 32680 35148 32732 35154
rect 32680 35090 32732 35096
rect 32036 35080 32088 35086
rect 32036 35022 32088 35028
rect 32048 33998 32076 35022
rect 33612 34066 33640 36110
rect 33600 34060 33652 34066
rect 33600 34002 33652 34008
rect 32036 33992 32088 33998
rect 32036 33934 32088 33940
rect 32220 33924 32272 33930
rect 32220 33866 32272 33872
rect 32232 33114 32260 33866
rect 33324 33856 33376 33862
rect 33324 33798 33376 33804
rect 32220 33108 32272 33114
rect 32220 33050 32272 33056
rect 32496 32904 32548 32910
rect 32496 32846 32548 32852
rect 32312 32564 32364 32570
rect 32312 32506 32364 32512
rect 32220 32428 32272 32434
rect 32220 32370 32272 32376
rect 32232 31482 32260 32370
rect 32324 31822 32352 32506
rect 32508 32502 32536 32846
rect 32496 32496 32548 32502
rect 32496 32438 32548 32444
rect 33336 32434 33364 33798
rect 33612 33522 33640 34002
rect 33600 33516 33652 33522
rect 33600 33458 33652 33464
rect 33612 32910 33640 33458
rect 33600 32904 33652 32910
rect 33600 32846 33652 32852
rect 33324 32428 33376 32434
rect 33324 32370 33376 32376
rect 32312 31816 32364 31822
rect 32312 31758 32364 31764
rect 32220 31476 32272 31482
rect 32220 31418 32272 31424
rect 31944 31136 31996 31142
rect 31944 31078 31996 31084
rect 32232 30326 32260 31418
rect 32324 30802 32352 31758
rect 33140 31340 33192 31346
rect 33140 31282 33192 31288
rect 32312 30796 32364 30802
rect 32312 30738 32364 30744
rect 32312 30592 32364 30598
rect 32312 30534 32364 30540
rect 32404 30592 32456 30598
rect 32404 30534 32456 30540
rect 32956 30592 33008 30598
rect 32956 30534 33008 30540
rect 32324 30326 32352 30534
rect 32220 30320 32272 30326
rect 32220 30262 32272 30268
rect 32312 30320 32364 30326
rect 32312 30262 32364 30268
rect 32416 30258 32444 30534
rect 32404 30252 32456 30258
rect 32404 30194 32456 30200
rect 32220 30116 32272 30122
rect 32220 30058 32272 30064
rect 31760 29028 31812 29034
rect 31760 28970 31812 28976
rect 31772 27062 31800 28970
rect 31760 27056 31812 27062
rect 31760 26998 31812 27004
rect 32232 26518 32260 30058
rect 32772 28076 32824 28082
rect 32772 28018 32824 28024
rect 32784 27674 32812 28018
rect 32772 27668 32824 27674
rect 32772 27610 32824 27616
rect 32784 27402 32812 27610
rect 32968 27470 32996 30534
rect 33152 29782 33180 31282
rect 33140 29776 33192 29782
rect 33140 29718 33192 29724
rect 33152 29306 33180 29718
rect 33140 29300 33192 29306
rect 33140 29242 33192 29248
rect 33152 27690 33180 29242
rect 33152 27662 33272 27690
rect 33140 27600 33192 27606
rect 33140 27542 33192 27548
rect 32956 27464 33008 27470
rect 32956 27406 33008 27412
rect 32772 27396 32824 27402
rect 32772 27338 32824 27344
rect 32404 27328 32456 27334
rect 32404 27270 32456 27276
rect 32588 27328 32640 27334
rect 32588 27270 32640 27276
rect 32220 26512 32272 26518
rect 32220 26454 32272 26460
rect 32036 25220 32088 25226
rect 32036 25162 32088 25168
rect 32048 24750 32076 25162
rect 32416 24954 32444 27270
rect 32600 26994 32628 27270
rect 32588 26988 32640 26994
rect 32588 26930 32640 26936
rect 32772 26988 32824 26994
rect 32772 26930 32824 26936
rect 32784 26518 32812 26930
rect 32772 26512 32824 26518
rect 32772 26454 32824 26460
rect 32956 26376 33008 26382
rect 33152 26330 33180 27542
rect 33244 27470 33272 27662
rect 33232 27464 33284 27470
rect 33232 27406 33284 27412
rect 33232 26784 33284 26790
rect 33232 26726 33284 26732
rect 33008 26324 33180 26330
rect 32956 26318 33180 26324
rect 32968 26302 33180 26318
rect 32772 26240 32824 26246
rect 32772 26182 32824 26188
rect 32784 26042 32812 26182
rect 32772 26036 32824 26042
rect 32772 25978 32824 25984
rect 33244 25974 33272 26726
rect 33336 26382 33364 32370
rect 33600 31408 33652 31414
rect 33600 31350 33652 31356
rect 33508 31272 33560 31278
rect 33508 31214 33560 31220
rect 33520 30297 33548 31214
rect 33612 30326 33640 31350
rect 33600 30320 33652 30326
rect 33506 30288 33562 30297
rect 33600 30262 33652 30268
rect 33506 30223 33508 30232
rect 33560 30223 33562 30232
rect 33508 30194 33560 30200
rect 33520 29646 33548 30194
rect 33600 30048 33652 30054
rect 33600 29990 33652 29996
rect 33508 29640 33560 29646
rect 33508 29582 33560 29588
rect 33416 29504 33468 29510
rect 33416 29446 33468 29452
rect 33324 26376 33376 26382
rect 33324 26318 33376 26324
rect 33232 25968 33284 25974
rect 33232 25910 33284 25916
rect 33140 25696 33192 25702
rect 33140 25638 33192 25644
rect 33152 25294 33180 25638
rect 33140 25288 33192 25294
rect 33140 25230 33192 25236
rect 32496 25152 32548 25158
rect 32496 25094 32548 25100
rect 32508 24954 32536 25094
rect 32404 24948 32456 24954
rect 32404 24890 32456 24896
rect 32496 24948 32548 24954
rect 32496 24890 32548 24896
rect 32036 24744 32088 24750
rect 32036 24686 32088 24692
rect 32508 23866 32536 24890
rect 32496 23860 32548 23866
rect 32496 23802 32548 23808
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 31944 23044 31996 23050
rect 31944 22986 31996 22992
rect 32036 23044 32088 23050
rect 32036 22986 32088 22992
rect 31852 21480 31904 21486
rect 31852 21422 31904 21428
rect 31588 12406 31708 12434
rect 31024 12300 31076 12306
rect 31024 12242 31076 12248
rect 31036 11218 31064 12242
rect 31208 12232 31260 12238
rect 31208 12174 31260 12180
rect 31220 11762 31248 12174
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31116 11756 31168 11762
rect 31116 11698 31168 11704
rect 31208 11756 31260 11762
rect 31208 11698 31260 11704
rect 31024 11212 31076 11218
rect 31024 11154 31076 11160
rect 30932 11144 30984 11150
rect 30932 11086 30984 11092
rect 30944 8838 30972 11086
rect 31128 10810 31156 11698
rect 31116 10804 31168 10810
rect 31116 10746 31168 10752
rect 31220 10130 31248 11698
rect 31404 11082 31432 12038
rect 31484 11756 31536 11762
rect 31484 11698 31536 11704
rect 31392 11076 31444 11082
rect 31392 11018 31444 11024
rect 31496 11014 31524 11698
rect 31484 11008 31536 11014
rect 31484 10950 31536 10956
rect 31208 10124 31260 10130
rect 31208 10066 31260 10072
rect 31300 8968 31352 8974
rect 31300 8910 31352 8916
rect 30932 8832 30984 8838
rect 30932 8774 30984 8780
rect 30944 8430 30972 8774
rect 30932 8424 30984 8430
rect 30932 8366 30984 8372
rect 30944 7002 30972 8366
rect 31312 7478 31340 8910
rect 31392 7880 31444 7886
rect 31392 7822 31444 7828
rect 31404 7546 31432 7822
rect 31392 7540 31444 7546
rect 31392 7482 31444 7488
rect 31300 7472 31352 7478
rect 31300 7414 31352 7420
rect 31116 7404 31168 7410
rect 31116 7346 31168 7352
rect 30932 6996 30984 7002
rect 30932 6938 30984 6944
rect 31128 6798 31156 7346
rect 31312 7002 31340 7414
rect 31300 6996 31352 7002
rect 31300 6938 31352 6944
rect 31116 6792 31168 6798
rect 31116 6734 31168 6740
rect 31128 6322 31156 6734
rect 31116 6316 31168 6322
rect 31116 6258 31168 6264
rect 31024 5704 31076 5710
rect 31024 5646 31076 5652
rect 30288 4616 30340 4622
rect 30288 4558 30340 4564
rect 30840 4616 30892 4622
rect 30840 4558 30892 4564
rect 30656 4480 30708 4486
rect 30656 4422 30708 4428
rect 29920 4276 29972 4282
rect 29920 4218 29972 4224
rect 29932 3641 29960 4218
rect 29918 3632 29974 3641
rect 29918 3567 29974 3576
rect 30668 3534 30696 4422
rect 30852 4282 30880 4558
rect 30840 4276 30892 4282
rect 30840 4218 30892 4224
rect 31036 3602 31064 5646
rect 31128 4622 31156 6258
rect 31588 5098 31616 12406
rect 31668 11620 31720 11626
rect 31668 11562 31720 11568
rect 31680 11014 31708 11562
rect 31668 11008 31720 11014
rect 31668 10950 31720 10956
rect 31864 9178 31892 21422
rect 31956 19854 31984 22986
rect 32048 22030 32076 22986
rect 32220 22976 32272 22982
rect 32220 22918 32272 22924
rect 32232 22710 32260 22918
rect 33048 22772 33100 22778
rect 33048 22714 33100 22720
rect 32128 22704 32180 22710
rect 32126 22672 32128 22681
rect 32220 22704 32272 22710
rect 32180 22672 32182 22681
rect 32220 22646 32272 22652
rect 32126 22607 32182 22616
rect 32312 22636 32364 22642
rect 32036 22024 32088 22030
rect 32036 21966 32088 21972
rect 32140 21962 32168 22607
rect 32864 22636 32916 22642
rect 32312 22578 32364 22584
rect 32692 22596 32864 22624
rect 32128 21956 32180 21962
rect 32128 21898 32180 21904
rect 32036 21684 32088 21690
rect 32036 21626 32088 21632
rect 32048 21146 32076 21626
rect 32036 21140 32088 21146
rect 32036 21082 32088 21088
rect 31944 19848 31996 19854
rect 31944 19790 31996 19796
rect 31956 18358 31984 19790
rect 31944 18352 31996 18358
rect 31944 18294 31996 18300
rect 31956 17882 31984 18294
rect 31944 17876 31996 17882
rect 31944 17818 31996 17824
rect 31944 17536 31996 17542
rect 32048 17524 32076 21082
rect 32140 19378 32168 21898
rect 32220 20800 32272 20806
rect 32220 20742 32272 20748
rect 32232 20505 32260 20742
rect 32218 20496 32274 20505
rect 32324 20466 32352 22578
rect 32692 20466 32720 22596
rect 32864 22578 32916 22584
rect 32956 22432 33008 22438
rect 32956 22374 33008 22380
rect 32968 21350 32996 22374
rect 33060 22030 33088 22714
rect 33152 22642 33180 23802
rect 33324 23588 33376 23594
rect 33324 23530 33376 23536
rect 33232 23044 33284 23050
rect 33232 22986 33284 22992
rect 33244 22778 33272 22986
rect 33232 22772 33284 22778
rect 33232 22714 33284 22720
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 33140 22432 33192 22438
rect 33140 22374 33192 22380
rect 33048 22024 33100 22030
rect 33048 21966 33100 21972
rect 33152 21554 33180 22374
rect 33336 22098 33364 23530
rect 33324 22092 33376 22098
rect 33324 22034 33376 22040
rect 33428 22030 33456 29446
rect 33520 29170 33548 29582
rect 33508 29164 33560 29170
rect 33508 29106 33560 29112
rect 33508 27872 33560 27878
rect 33508 27814 33560 27820
rect 33520 23798 33548 27814
rect 33508 23792 33560 23798
rect 33508 23734 33560 23740
rect 33508 23656 33560 23662
rect 33508 23598 33560 23604
rect 33416 22024 33468 22030
rect 33416 21966 33468 21972
rect 33140 21548 33192 21554
rect 33140 21490 33192 21496
rect 32956 21344 33008 21350
rect 32956 21286 33008 21292
rect 32862 20496 32918 20505
rect 32218 20431 32274 20440
rect 32312 20460 32364 20466
rect 32232 19718 32260 20431
rect 32312 20402 32364 20408
rect 32680 20460 32732 20466
rect 32862 20431 32864 20440
rect 32680 20402 32732 20408
rect 32916 20431 32918 20440
rect 32864 20402 32916 20408
rect 32220 19712 32272 19718
rect 32220 19654 32272 19660
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 31996 17496 32076 17524
rect 31944 17478 31996 17484
rect 31956 11762 31984 17478
rect 32036 16584 32088 16590
rect 32036 16526 32088 16532
rect 32048 15502 32076 16526
rect 32036 15496 32088 15502
rect 32036 15438 32088 15444
rect 32048 15026 32076 15438
rect 32036 15020 32088 15026
rect 32036 14962 32088 14968
rect 32048 14482 32076 14962
rect 32036 14476 32088 14482
rect 32036 14418 32088 14424
rect 31944 11756 31996 11762
rect 31944 11698 31996 11704
rect 32128 11688 32180 11694
rect 32128 11630 32180 11636
rect 31944 10668 31996 10674
rect 31944 10610 31996 10616
rect 31956 10470 31984 10610
rect 31944 10464 31996 10470
rect 31944 10406 31996 10412
rect 32140 10062 32168 11630
rect 32232 11054 32260 19654
rect 32324 18766 32352 20402
rect 32404 19440 32456 19446
rect 32404 19382 32456 19388
rect 32312 18760 32364 18766
rect 32312 18702 32364 18708
rect 32324 16794 32352 18702
rect 32416 18358 32444 19382
rect 32692 18630 32720 20402
rect 33048 20324 33100 20330
rect 33048 20266 33100 20272
rect 32864 20256 32916 20262
rect 32864 20198 32916 20204
rect 32876 19854 32904 20198
rect 33060 20058 33088 20266
rect 33048 20052 33100 20058
rect 33048 19994 33100 20000
rect 32864 19848 32916 19854
rect 32864 19790 32916 19796
rect 33232 19372 33284 19378
rect 33232 19314 33284 19320
rect 33244 18970 33272 19314
rect 33232 18964 33284 18970
rect 33232 18906 33284 18912
rect 32588 18624 32640 18630
rect 32588 18566 32640 18572
rect 32680 18624 32732 18630
rect 32680 18566 32732 18572
rect 32600 18426 32628 18566
rect 32588 18420 32640 18426
rect 32588 18362 32640 18368
rect 32404 18352 32456 18358
rect 32404 18294 32456 18300
rect 32496 17672 32548 17678
rect 32496 17614 32548 17620
rect 32586 17640 32642 17649
rect 32312 16788 32364 16794
rect 32312 16730 32364 16736
rect 32508 16590 32536 17614
rect 32586 17575 32588 17584
rect 32640 17575 32642 17584
rect 32692 17626 32720 18566
rect 32956 18148 33008 18154
rect 32956 18090 33008 18096
rect 32772 17648 32824 17654
rect 32692 17598 32772 17626
rect 32588 17546 32640 17552
rect 32692 17134 32720 17598
rect 32772 17590 32824 17596
rect 32772 17332 32824 17338
rect 32772 17274 32824 17280
rect 32680 17128 32732 17134
rect 32680 17070 32732 17076
rect 32692 16658 32720 17070
rect 32680 16652 32732 16658
rect 32680 16594 32732 16600
rect 32496 16584 32548 16590
rect 32496 16526 32548 16532
rect 32312 16516 32364 16522
rect 32312 16458 32364 16464
rect 32324 13258 32352 16458
rect 32588 15904 32640 15910
rect 32588 15846 32640 15852
rect 32600 15706 32628 15846
rect 32588 15700 32640 15706
rect 32588 15642 32640 15648
rect 32312 13252 32364 13258
rect 32312 13194 32364 13200
rect 32324 12986 32352 13194
rect 32588 13184 32640 13190
rect 32588 13126 32640 13132
rect 32312 12980 32364 12986
rect 32312 12922 32364 12928
rect 32600 12170 32628 13126
rect 32680 12844 32732 12850
rect 32680 12786 32732 12792
rect 32588 12164 32640 12170
rect 32588 12106 32640 12112
rect 32232 11026 32352 11054
rect 32324 10554 32352 11026
rect 32324 10526 32536 10554
rect 32404 10464 32456 10470
rect 32404 10406 32456 10412
rect 32128 10056 32180 10062
rect 32128 9998 32180 10004
rect 32140 9586 32168 9998
rect 32128 9580 32180 9586
rect 32128 9522 32180 9528
rect 32312 9580 32364 9586
rect 32312 9522 32364 9528
rect 31852 9172 31904 9178
rect 31852 9114 31904 9120
rect 32324 8090 32352 9522
rect 32416 8974 32444 10406
rect 32508 9586 32536 10526
rect 32496 9580 32548 9586
rect 32496 9522 32548 9528
rect 32404 8968 32456 8974
rect 32404 8910 32456 8916
rect 32496 8832 32548 8838
rect 32496 8774 32548 8780
rect 32508 8498 32536 8774
rect 32600 8566 32628 12106
rect 32692 11694 32720 12786
rect 32680 11688 32732 11694
rect 32680 11630 32732 11636
rect 32680 8968 32732 8974
rect 32680 8910 32732 8916
rect 32588 8560 32640 8566
rect 32588 8502 32640 8508
rect 32692 8498 32720 8910
rect 32784 8634 32812 17274
rect 32968 16590 32996 18090
rect 33048 18080 33100 18086
rect 33048 18022 33100 18028
rect 33060 17746 33088 18022
rect 33048 17740 33100 17746
rect 33048 17682 33100 17688
rect 33140 17536 33192 17542
rect 33140 17478 33192 17484
rect 33152 17270 33180 17478
rect 33520 17338 33548 23598
rect 33612 21622 33640 29990
rect 33704 28218 33732 36518
rect 33796 36174 33824 36751
rect 33784 36168 33836 36174
rect 33784 36110 33836 36116
rect 33796 34746 33824 36110
rect 33784 34740 33836 34746
rect 33784 34682 33836 34688
rect 33796 33998 33824 34682
rect 33784 33992 33836 33998
rect 33784 33934 33836 33940
rect 33796 32910 33824 33934
rect 33784 32904 33836 32910
rect 33784 32846 33836 32852
rect 33784 30932 33836 30938
rect 33784 30874 33836 30880
rect 33692 28212 33744 28218
rect 33692 28154 33744 28160
rect 33796 27996 33824 30874
rect 33888 30258 33916 36790
rect 34072 36378 34100 36790
rect 34060 36372 34112 36378
rect 34060 36314 34112 36320
rect 34164 33658 34192 37606
rect 34256 36786 34284 37810
rect 34532 36922 34560 37810
rect 34520 36916 34572 36922
rect 34520 36858 34572 36864
rect 34624 36802 34652 37946
rect 35348 37664 35400 37670
rect 35348 37606 35400 37612
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35360 37262 35388 37606
rect 34796 37256 34848 37262
rect 34796 37198 34848 37204
rect 35348 37256 35400 37262
rect 35348 37198 35400 37204
rect 34244 36780 34296 36786
rect 34244 36722 34296 36728
rect 34532 36774 34652 36802
rect 34532 36666 34560 36774
rect 34440 36650 34560 36666
rect 34428 36644 34560 36650
rect 34480 36638 34560 36644
rect 34428 36586 34480 36592
rect 34152 33652 34204 33658
rect 34152 33594 34204 33600
rect 34060 33516 34112 33522
rect 34060 33458 34112 33464
rect 34072 33114 34100 33458
rect 34060 33108 34112 33114
rect 34060 33050 34112 33056
rect 33968 30320 34020 30326
rect 33968 30262 34020 30268
rect 33876 30252 33928 30258
rect 33876 30194 33928 30200
rect 33980 30138 34008 30262
rect 34060 30184 34112 30190
rect 33980 30132 34060 30138
rect 33980 30126 34112 30132
rect 33980 30110 34100 30126
rect 33980 29646 34008 30110
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 33980 28626 34008 29582
rect 34164 29510 34192 33594
rect 34428 33516 34480 33522
rect 34428 33458 34480 33464
rect 34440 32978 34468 33458
rect 34532 33454 34560 36638
rect 34704 36576 34756 36582
rect 34704 36518 34756 36524
rect 34716 36174 34744 36518
rect 34808 36242 34836 37198
rect 35532 37120 35584 37126
rect 35532 37062 35584 37068
rect 35346 36816 35402 36825
rect 35544 36786 35572 37062
rect 35346 36751 35348 36760
rect 35400 36751 35402 36760
rect 35532 36780 35584 36786
rect 35348 36722 35400 36728
rect 35532 36722 35584 36728
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34796 36236 34848 36242
rect 34796 36178 34848 36184
rect 34704 36168 34756 36174
rect 34704 36110 34756 36116
rect 34704 36032 34756 36038
rect 34704 35974 34756 35980
rect 34612 33992 34664 33998
rect 34612 33934 34664 33940
rect 34520 33448 34572 33454
rect 34520 33390 34572 33396
rect 34520 33312 34572 33318
rect 34520 33254 34572 33260
rect 34428 32972 34480 32978
rect 34428 32914 34480 32920
rect 34440 30394 34468 32914
rect 34532 32910 34560 33254
rect 34624 33114 34652 33934
rect 34612 33108 34664 33114
rect 34612 33050 34664 33056
rect 34520 32904 34572 32910
rect 34520 32846 34572 32852
rect 34428 30388 34480 30394
rect 34428 30330 34480 30336
rect 34334 30288 34390 30297
rect 34334 30223 34336 30232
rect 34388 30223 34390 30232
rect 34336 30194 34388 30200
rect 34336 30048 34388 30054
rect 34336 29990 34388 29996
rect 34244 29844 34296 29850
rect 34244 29786 34296 29792
rect 34152 29504 34204 29510
rect 34152 29446 34204 29452
rect 34152 29096 34204 29102
rect 34152 29038 34204 29044
rect 33968 28620 34020 28626
rect 33968 28562 34020 28568
rect 34164 28558 34192 29038
rect 34152 28552 34204 28558
rect 34152 28494 34204 28500
rect 34164 28082 34192 28494
rect 34152 28076 34204 28082
rect 34152 28018 34204 28024
rect 33796 27968 33916 27996
rect 33784 27668 33836 27674
rect 33784 27610 33836 27616
rect 33692 27396 33744 27402
rect 33692 27338 33744 27344
rect 33704 26042 33732 27338
rect 33796 26450 33824 27610
rect 33888 26450 33916 27968
rect 34164 27606 34192 28018
rect 34152 27600 34204 27606
rect 34152 27542 34204 27548
rect 34256 27010 34284 29786
rect 34164 26994 34284 27010
rect 34152 26988 34284 26994
rect 34204 26982 34284 26988
rect 34152 26930 34204 26936
rect 33968 26920 34020 26926
rect 33968 26862 34020 26868
rect 33980 26586 34008 26862
rect 34164 26858 34192 26930
rect 34152 26852 34204 26858
rect 34152 26794 34204 26800
rect 33968 26580 34020 26586
rect 33968 26522 34020 26528
rect 33784 26444 33836 26450
rect 33784 26386 33836 26392
rect 33876 26444 33928 26450
rect 33876 26386 33928 26392
rect 33692 26036 33744 26042
rect 33692 25978 33744 25984
rect 33980 24818 34008 26522
rect 34060 25288 34112 25294
rect 34060 25230 34112 25236
rect 33968 24812 34020 24818
rect 33968 24754 34020 24760
rect 33876 24608 33928 24614
rect 33876 24550 33928 24556
rect 33692 23520 33744 23526
rect 33692 23462 33744 23468
rect 33704 22778 33732 23462
rect 33888 23322 33916 24550
rect 33876 23316 33928 23322
rect 33876 23258 33928 23264
rect 33692 22772 33744 22778
rect 33692 22714 33744 22720
rect 33784 22500 33836 22506
rect 33784 22442 33836 22448
rect 33692 21956 33744 21962
rect 33692 21898 33744 21904
rect 33600 21616 33652 21622
rect 33600 21558 33652 21564
rect 33508 17332 33560 17338
rect 33508 17274 33560 17280
rect 33140 17264 33192 17270
rect 33140 17206 33192 17212
rect 32956 16584 33008 16590
rect 32956 16526 33008 16532
rect 33232 15496 33284 15502
rect 33232 15438 33284 15444
rect 33600 15496 33652 15502
rect 33600 15438 33652 15444
rect 33244 14822 33272 15438
rect 33232 14816 33284 14822
rect 33232 14758 33284 14764
rect 32864 12844 32916 12850
rect 32864 12786 32916 12792
rect 32956 12844 33008 12850
rect 32956 12786 33008 12792
rect 32876 12442 32904 12786
rect 32864 12436 32916 12442
rect 32864 12378 32916 12384
rect 32968 12238 32996 12786
rect 33244 12646 33272 14758
rect 33612 14482 33640 15438
rect 33600 14476 33652 14482
rect 33600 14418 33652 14424
rect 33416 14408 33468 14414
rect 33416 14350 33468 14356
rect 33428 13938 33456 14350
rect 33416 13932 33468 13938
rect 33416 13874 33468 13880
rect 33612 13870 33640 14418
rect 33600 13864 33652 13870
rect 33600 13806 33652 13812
rect 33324 13252 33376 13258
rect 33324 13194 33376 13200
rect 33336 12986 33364 13194
rect 33324 12980 33376 12986
rect 33324 12922 33376 12928
rect 33232 12640 33284 12646
rect 33232 12582 33284 12588
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32968 9518 32996 12174
rect 33048 11552 33100 11558
rect 33048 11494 33100 11500
rect 33060 10742 33088 11494
rect 33416 11348 33468 11354
rect 33416 11290 33468 11296
rect 33048 10736 33100 10742
rect 33048 10678 33100 10684
rect 32956 9512 33008 9518
rect 32956 9454 33008 9460
rect 33428 8974 33456 11290
rect 33600 9376 33652 9382
rect 33600 9318 33652 9324
rect 33140 8968 33192 8974
rect 33140 8910 33192 8916
rect 33416 8968 33468 8974
rect 33416 8910 33468 8916
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 32404 8492 32456 8498
rect 32404 8434 32456 8440
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 32312 8084 32364 8090
rect 32312 8026 32364 8032
rect 31576 5092 31628 5098
rect 31576 5034 31628 5040
rect 32416 4622 32444 8434
rect 33152 6390 33180 8910
rect 33612 7478 33640 9318
rect 33704 9178 33732 21898
rect 33796 19666 33824 22442
rect 33888 20482 33916 23258
rect 34072 23186 34100 25230
rect 34348 23798 34376 29990
rect 34440 29238 34468 30330
rect 34532 29646 34560 32846
rect 34612 30728 34664 30734
rect 34612 30670 34664 30676
rect 34624 30326 34652 30670
rect 34612 30320 34664 30326
rect 34612 30262 34664 30268
rect 34520 29640 34572 29646
rect 34520 29582 34572 29588
rect 34428 29232 34480 29238
rect 34428 29174 34480 29180
rect 34428 28484 34480 28490
rect 34428 28426 34480 28432
rect 34440 28082 34468 28426
rect 34612 28416 34664 28422
rect 34612 28358 34664 28364
rect 34428 28076 34480 28082
rect 34428 28018 34480 28024
rect 34440 27674 34468 28018
rect 34428 27668 34480 27674
rect 34428 27610 34480 27616
rect 34428 27464 34480 27470
rect 34428 27406 34480 27412
rect 34440 27146 34468 27406
rect 34440 27118 34560 27146
rect 34532 26994 34560 27118
rect 34428 26988 34480 26994
rect 34428 26930 34480 26936
rect 34520 26988 34572 26994
rect 34520 26930 34572 26936
rect 34440 26450 34468 26930
rect 34520 26784 34572 26790
rect 34520 26726 34572 26732
rect 34428 26444 34480 26450
rect 34428 26386 34480 26392
rect 34532 26382 34560 26726
rect 34520 26376 34572 26382
rect 34520 26318 34572 26324
rect 34336 23792 34388 23798
rect 34336 23734 34388 23740
rect 34060 23180 34112 23186
rect 34060 23122 34112 23128
rect 34244 23112 34296 23118
rect 34244 23054 34296 23060
rect 34060 22704 34112 22710
rect 34058 22672 34060 22681
rect 34112 22672 34114 22681
rect 33968 22636 34020 22642
rect 34256 22642 34284 23054
rect 34058 22607 34114 22616
rect 34244 22636 34296 22642
rect 33968 22578 34020 22584
rect 34244 22578 34296 22584
rect 33980 20618 34008 22578
rect 34624 21690 34652 28358
rect 34716 28082 34744 35974
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34980 33856 35032 33862
rect 34980 33798 35032 33804
rect 34992 33454 35020 33798
rect 34980 33448 35032 33454
rect 34980 33390 35032 33396
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34796 33108 34848 33114
rect 34796 33050 34848 33056
rect 34808 30258 34836 33050
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35348 31340 35400 31346
rect 35348 31282 35400 31288
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35360 30666 35388 31282
rect 35348 30660 35400 30666
rect 35400 30620 35480 30648
rect 35348 30602 35400 30608
rect 34796 30252 34848 30258
rect 34796 30194 34848 30200
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35452 29866 35480 30620
rect 35360 29850 35480 29866
rect 35348 29844 35480 29850
rect 35400 29838 35480 29844
rect 35348 29786 35400 29792
rect 35360 29170 35388 29786
rect 35440 29776 35492 29782
rect 35440 29718 35492 29724
rect 35452 29238 35480 29718
rect 35440 29232 35492 29238
rect 35440 29174 35492 29180
rect 35348 29164 35400 29170
rect 35348 29106 35400 29112
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35360 28082 35388 29106
rect 35452 28626 35480 29174
rect 35440 28620 35492 28626
rect 35440 28562 35492 28568
rect 35544 28558 35572 36722
rect 35716 34672 35768 34678
rect 35716 34614 35768 34620
rect 35728 33998 35756 34614
rect 35716 33992 35768 33998
rect 35716 33934 35768 33940
rect 35728 30802 35756 33934
rect 35716 30796 35768 30802
rect 35716 30738 35768 30744
rect 35532 28552 35584 28558
rect 35532 28494 35584 28500
rect 34704 28076 34756 28082
rect 34704 28018 34756 28024
rect 35348 28076 35400 28082
rect 35348 28018 35400 28024
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35440 26988 35492 26994
rect 35440 26930 35492 26936
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35452 26586 35480 26930
rect 35440 26580 35492 26586
rect 35440 26522 35492 26528
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35624 25152 35676 25158
rect 35624 25094 35676 25100
rect 35636 24682 35664 25094
rect 35716 24744 35768 24750
rect 35716 24686 35768 24692
rect 35624 24676 35676 24682
rect 35624 24618 35676 24624
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35532 23724 35584 23730
rect 35532 23666 35584 23672
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35544 21894 35572 23666
rect 35636 22642 35664 24618
rect 35728 23186 35756 24686
rect 35716 23180 35768 23186
rect 35716 23122 35768 23128
rect 35624 22636 35676 22642
rect 35624 22578 35676 22584
rect 35532 21888 35584 21894
rect 35532 21830 35584 21836
rect 34612 21684 34664 21690
rect 34612 21626 34664 21632
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 33980 20590 34192 20618
rect 33888 20454 34008 20482
rect 33796 19638 33916 19666
rect 33784 19508 33836 19514
rect 33784 19450 33836 19456
rect 33796 18222 33824 19450
rect 33888 18426 33916 19638
rect 33876 18420 33928 18426
rect 33876 18362 33928 18368
rect 33784 18216 33836 18222
rect 33784 18158 33836 18164
rect 33888 17066 33916 18362
rect 33876 17060 33928 17066
rect 33876 17002 33928 17008
rect 33980 16590 34008 20454
rect 34164 18358 34192 20590
rect 34244 20256 34296 20262
rect 34244 20198 34296 20204
rect 34256 19378 34284 20198
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34152 18352 34204 18358
rect 34152 18294 34204 18300
rect 34164 17338 34192 18294
rect 35624 18080 35676 18086
rect 35624 18022 35676 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34612 17808 34664 17814
rect 34612 17750 34664 17756
rect 34152 17332 34204 17338
rect 34152 17274 34204 17280
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 33968 16584 34020 16590
rect 33968 16526 34020 16532
rect 34532 16522 34560 17138
rect 34520 16516 34572 16522
rect 34520 16458 34572 16464
rect 34428 13320 34480 13326
rect 34428 13262 34480 13268
rect 34336 12776 34388 12782
rect 34336 12718 34388 12724
rect 33876 12640 33928 12646
rect 33876 12582 33928 12588
rect 33888 12442 33916 12582
rect 33876 12436 33928 12442
rect 33876 12378 33928 12384
rect 34348 12238 34376 12718
rect 34336 12232 34388 12238
rect 34336 12174 34388 12180
rect 34348 11762 34376 12174
rect 34440 11898 34468 13262
rect 34428 11892 34480 11898
rect 34428 11834 34480 11840
rect 34336 11756 34388 11762
rect 34336 11698 34388 11704
rect 34520 10464 34572 10470
rect 34520 10406 34572 10412
rect 33692 9172 33744 9178
rect 33692 9114 33744 9120
rect 34532 7546 34560 10406
rect 34520 7540 34572 7546
rect 34520 7482 34572 7488
rect 33600 7472 33652 7478
rect 33600 7414 33652 7420
rect 34152 6724 34204 6730
rect 34152 6666 34204 6672
rect 34164 6458 34192 6666
rect 34520 6656 34572 6662
rect 34520 6598 34572 6604
rect 34152 6452 34204 6458
rect 34152 6394 34204 6400
rect 33140 6384 33192 6390
rect 34428 6384 34480 6390
rect 33140 6326 33192 6332
rect 34426 6352 34428 6361
rect 34480 6352 34482 6361
rect 33152 5914 33180 6326
rect 34426 6287 34482 6296
rect 34532 5914 34560 6598
rect 33140 5908 33192 5914
rect 33140 5850 33192 5856
rect 34520 5908 34572 5914
rect 34520 5850 34572 5856
rect 31116 4616 31168 4622
rect 31116 4558 31168 4564
rect 32404 4616 32456 4622
rect 32404 4558 32456 4564
rect 32416 3738 32444 4558
rect 32404 3732 32456 3738
rect 32404 3674 32456 3680
rect 31024 3596 31076 3602
rect 31024 3538 31076 3544
rect 30656 3528 30708 3534
rect 30656 3470 30708 3476
rect 32772 2984 32824 2990
rect 32772 2926 32824 2932
rect 29736 2848 29788 2854
rect 29736 2790 29788 2796
rect 30012 2848 30064 2854
rect 30012 2790 30064 2796
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 31668 2848 31720 2854
rect 31668 2790 31720 2796
rect 32220 2848 32272 2854
rect 32220 2790 32272 2796
rect 29276 2644 29328 2650
rect 29276 2586 29328 2592
rect 29460 2440 29512 2446
rect 29460 2382 29512 2388
rect 29472 800 29500 2382
rect 29748 800 29776 2790
rect 30024 800 30052 2790
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 30300 800 30328 2382
rect 30576 800 30604 2790
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 31116 2440 31168 2446
rect 31116 2382 31168 2388
rect 31392 2440 31444 2446
rect 31392 2382 31444 2388
rect 30852 800 30880 2382
rect 31128 800 31156 2382
rect 31404 800 31432 2382
rect 31680 800 31708 2790
rect 31944 2508 31996 2514
rect 31944 2450 31996 2456
rect 31956 800 31984 2450
rect 32232 800 32260 2790
rect 32496 2440 32548 2446
rect 32496 2382 32548 2388
rect 32508 800 32536 2382
rect 32784 800 32812 2926
rect 33324 2916 33376 2922
rect 33324 2858 33376 2864
rect 34428 2916 34480 2922
rect 34428 2858 34480 2864
rect 33048 2508 33100 2514
rect 33048 2450 33100 2456
rect 33060 800 33088 2450
rect 33336 800 33364 2858
rect 33876 2848 33928 2854
rect 33876 2790 33928 2796
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 33612 800 33640 2382
rect 33888 800 33916 2790
rect 34152 2576 34204 2582
rect 34152 2518 34204 2524
rect 34164 800 34192 2518
rect 34440 800 34468 2858
rect 34624 2106 34652 17750
rect 35636 17678 35664 18022
rect 35820 17814 35848 56306
rect 37844 55962 37872 57394
rect 37936 56506 37964 57394
rect 37924 56500 37976 56506
rect 37924 56442 37976 56448
rect 40972 56234 41000 57394
rect 42352 56710 42380 57394
rect 42340 56704 42392 56710
rect 42340 56646 42392 56652
rect 42352 56438 42380 56646
rect 42340 56432 42392 56438
rect 42340 56374 42392 56380
rect 44100 56234 44128 57394
rect 45664 56506 45692 57394
rect 47596 56506 47624 57394
rect 54956 57390 54984 59200
rect 56520 57882 56548 59200
rect 57518 57896 57574 57905
rect 56520 57854 56640 57882
rect 56612 57458 56640 57854
rect 57518 57831 57574 57840
rect 56600 57452 56652 57458
rect 56600 57394 56652 57400
rect 54944 57384 54996 57390
rect 54944 57326 54996 57332
rect 57532 57050 57560 57831
rect 58084 57458 58112 59200
rect 58438 59191 58494 59200
rect 58072 57452 58124 57458
rect 58072 57394 58124 57400
rect 57520 57044 57572 57050
rect 57520 56986 57572 56992
rect 57888 56840 57940 56846
rect 57888 56782 57940 56788
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 57900 56545 57928 56782
rect 57886 56536 57942 56545
rect 45652 56500 45704 56506
rect 45652 56442 45704 56448
rect 47584 56500 47636 56506
rect 57886 56471 57942 56480
rect 47584 56442 47636 56448
rect 58452 56370 58480 59191
rect 45560 56364 45612 56370
rect 45560 56306 45612 56312
rect 58440 56364 58492 56370
rect 58440 56306 58492 56312
rect 40960 56228 41012 56234
rect 40960 56170 41012 56176
rect 44088 56228 44140 56234
rect 44088 56170 44140 56176
rect 42064 56160 42116 56166
rect 42064 56102 42116 56108
rect 37832 55956 37884 55962
rect 37832 55898 37884 55904
rect 35992 33856 36044 33862
rect 35992 33798 36044 33804
rect 35900 33108 35952 33114
rect 35900 33050 35952 33056
rect 35912 31754 35940 33050
rect 36004 32910 36032 33798
rect 36268 33516 36320 33522
rect 36268 33458 36320 33464
rect 36280 32910 36308 33458
rect 35992 32904 36044 32910
rect 35992 32846 36044 32852
rect 36268 32904 36320 32910
rect 36268 32846 36320 32852
rect 36280 32570 36308 32846
rect 36268 32564 36320 32570
rect 36268 32506 36320 32512
rect 36280 31958 36308 32506
rect 36452 32020 36504 32026
rect 36452 31962 36504 31968
rect 36268 31952 36320 31958
rect 36268 31894 36320 31900
rect 36464 31822 36492 31962
rect 37556 31884 37608 31890
rect 37556 31826 37608 31832
rect 36268 31816 36320 31822
rect 36268 31758 36320 31764
rect 36452 31816 36504 31822
rect 36452 31758 36504 31764
rect 35912 31748 36044 31754
rect 35912 31726 35992 31748
rect 35912 30734 35940 31726
rect 35992 31690 36044 31696
rect 36176 31748 36228 31754
rect 36176 31690 36228 31696
rect 35900 30728 35952 30734
rect 35900 30670 35952 30676
rect 35912 30258 35940 30670
rect 36188 30598 36216 31690
rect 36280 31482 36308 31758
rect 36268 31476 36320 31482
rect 36268 31418 36320 31424
rect 37280 31340 37332 31346
rect 37280 31282 37332 31288
rect 36176 30592 36228 30598
rect 36176 30534 36228 30540
rect 36188 30258 36216 30534
rect 37292 30326 37320 31282
rect 37568 30802 37596 31826
rect 38936 31680 38988 31686
rect 38936 31622 38988 31628
rect 38948 31414 38976 31622
rect 38936 31408 38988 31414
rect 38936 31350 38988 31356
rect 37556 30796 37608 30802
rect 37556 30738 37608 30744
rect 37280 30320 37332 30326
rect 37280 30262 37332 30268
rect 35900 30252 35952 30258
rect 35900 30194 35952 30200
rect 36176 30252 36228 30258
rect 36176 30194 36228 30200
rect 36360 30252 36412 30258
rect 36360 30194 36412 30200
rect 37464 30252 37516 30258
rect 37464 30194 37516 30200
rect 36188 29714 36216 30194
rect 36372 30054 36400 30194
rect 36360 30048 36412 30054
rect 36360 29990 36412 29996
rect 36176 29708 36228 29714
rect 36176 29650 36228 29656
rect 36084 29164 36136 29170
rect 36084 29106 36136 29112
rect 36096 28558 36124 29106
rect 36188 29102 36216 29650
rect 37476 29646 37504 30194
rect 39672 30048 39724 30054
rect 39672 29990 39724 29996
rect 37464 29640 37516 29646
rect 37464 29582 37516 29588
rect 39304 29640 39356 29646
rect 39304 29582 39356 29588
rect 36728 29572 36780 29578
rect 36728 29514 36780 29520
rect 36636 29504 36688 29510
rect 36636 29446 36688 29452
rect 36648 29170 36676 29446
rect 36740 29306 36768 29514
rect 37476 29306 37504 29582
rect 36728 29300 36780 29306
rect 36728 29242 36780 29248
rect 37464 29300 37516 29306
rect 37464 29242 37516 29248
rect 36636 29164 36688 29170
rect 36636 29106 36688 29112
rect 36176 29096 36228 29102
rect 36176 29038 36228 29044
rect 36188 28694 36216 29038
rect 39316 28966 39344 29582
rect 39684 29238 39712 29990
rect 39672 29232 39724 29238
rect 39672 29174 39724 29180
rect 38752 28960 38804 28966
rect 38752 28902 38804 28908
rect 39304 28960 39356 28966
rect 39304 28902 39356 28908
rect 36176 28688 36228 28694
rect 36176 28630 36228 28636
rect 38764 28558 38792 28902
rect 36084 28552 36136 28558
rect 36084 28494 36136 28500
rect 36360 28552 36412 28558
rect 36360 28494 36412 28500
rect 38752 28552 38804 28558
rect 38752 28494 38804 28500
rect 35992 28484 36044 28490
rect 35992 28426 36044 28432
rect 36004 28218 36032 28426
rect 35992 28212 36044 28218
rect 35992 28154 36044 28160
rect 36004 27674 36032 28154
rect 35992 27668 36044 27674
rect 35992 27610 36044 27616
rect 36096 27130 36124 28494
rect 36176 28416 36228 28422
rect 36176 28358 36228 28364
rect 36188 28150 36216 28358
rect 36372 28218 36400 28494
rect 36360 28212 36412 28218
rect 36360 28154 36412 28160
rect 36176 28144 36228 28150
rect 36176 28086 36228 28092
rect 36084 27124 36136 27130
rect 36084 27066 36136 27072
rect 36912 26512 36964 26518
rect 36912 26454 36964 26460
rect 36360 25696 36412 25702
rect 36360 25638 36412 25644
rect 36084 24608 36136 24614
rect 36084 24550 36136 24556
rect 35992 23724 36044 23730
rect 35992 23666 36044 23672
rect 36004 22438 36032 23666
rect 35992 22432 36044 22438
rect 35992 22374 36044 22380
rect 36004 22030 36032 22374
rect 36096 22030 36124 24550
rect 36268 23724 36320 23730
rect 36268 23666 36320 23672
rect 36176 23044 36228 23050
rect 36176 22986 36228 22992
rect 36188 22778 36216 22986
rect 36176 22772 36228 22778
rect 36176 22714 36228 22720
rect 36280 22506 36308 23666
rect 36372 22642 36400 25638
rect 36924 23730 36952 26454
rect 38764 26382 38792 28494
rect 39948 26784 40000 26790
rect 39948 26726 40000 26732
rect 39960 26382 39988 26726
rect 37096 26376 37148 26382
rect 37096 26318 37148 26324
rect 38752 26376 38804 26382
rect 38752 26318 38804 26324
rect 39948 26376 40000 26382
rect 39948 26318 40000 26324
rect 37108 25362 37136 26318
rect 39764 26308 39816 26314
rect 39764 26250 39816 26256
rect 39856 26308 39908 26314
rect 39856 26250 39908 26256
rect 37280 25764 37332 25770
rect 37280 25706 37332 25712
rect 38568 25764 38620 25770
rect 38568 25706 38620 25712
rect 37096 25356 37148 25362
rect 37096 25298 37148 25304
rect 36912 23724 36964 23730
rect 36912 23666 36964 23672
rect 37292 23474 37320 25706
rect 37372 25696 37424 25702
rect 37372 25638 37424 25644
rect 37384 25294 37412 25638
rect 37372 25288 37424 25294
rect 37372 25230 37424 25236
rect 38580 25226 38608 25706
rect 39304 25696 39356 25702
rect 39304 25638 39356 25644
rect 39316 25498 39344 25638
rect 39776 25498 39804 26250
rect 39304 25492 39356 25498
rect 39304 25434 39356 25440
rect 39764 25492 39816 25498
rect 39764 25434 39816 25440
rect 39868 25294 39896 26250
rect 39960 25838 39988 26318
rect 40408 26240 40460 26246
rect 40408 26182 40460 26188
rect 40776 26240 40828 26246
rect 40776 26182 40828 26188
rect 39948 25832 40000 25838
rect 39948 25774 40000 25780
rect 38936 25288 38988 25294
rect 38936 25230 38988 25236
rect 39856 25288 39908 25294
rect 39856 25230 39908 25236
rect 37648 25220 37700 25226
rect 37648 25162 37700 25168
rect 38568 25220 38620 25226
rect 38568 25162 38620 25168
rect 37660 24750 37688 25162
rect 38948 24818 38976 25230
rect 39960 24818 39988 25774
rect 40224 25764 40276 25770
rect 40224 25706 40276 25712
rect 40236 25498 40264 25706
rect 40224 25492 40276 25498
rect 40224 25434 40276 25440
rect 40132 25288 40184 25294
rect 40132 25230 40184 25236
rect 40144 24954 40172 25230
rect 40132 24948 40184 24954
rect 40132 24890 40184 24896
rect 38936 24812 38988 24818
rect 38936 24754 38988 24760
rect 39764 24812 39816 24818
rect 39764 24754 39816 24760
rect 39948 24812 40000 24818
rect 39948 24754 40000 24760
rect 37648 24744 37700 24750
rect 37648 24686 37700 24692
rect 38660 24608 38712 24614
rect 38660 24550 38712 24556
rect 38672 24274 38700 24550
rect 38660 24268 38712 24274
rect 38660 24210 38712 24216
rect 37108 23446 37320 23474
rect 36728 22976 36780 22982
rect 36728 22918 36780 22924
rect 36740 22642 36768 22918
rect 36360 22636 36412 22642
rect 36360 22578 36412 22584
rect 36728 22636 36780 22642
rect 36728 22578 36780 22584
rect 37004 22636 37056 22642
rect 37004 22578 37056 22584
rect 36268 22500 36320 22506
rect 36268 22442 36320 22448
rect 35992 22024 36044 22030
rect 35992 21966 36044 21972
rect 36084 22024 36136 22030
rect 36084 21966 36136 21972
rect 35900 21344 35952 21350
rect 35900 21286 35952 21292
rect 35912 21146 35940 21286
rect 35900 21140 35952 21146
rect 35900 21082 35952 21088
rect 36004 19922 36032 21966
rect 36280 21962 36308 22442
rect 36268 21956 36320 21962
rect 36268 21898 36320 21904
rect 36280 20466 36308 21898
rect 36372 21350 36400 22578
rect 36360 21344 36412 21350
rect 36360 21286 36412 21292
rect 36912 20596 36964 20602
rect 36912 20538 36964 20544
rect 36268 20460 36320 20466
rect 36268 20402 36320 20408
rect 35992 19916 36044 19922
rect 35992 19858 36044 19864
rect 36004 19378 36032 19858
rect 36280 19514 36308 20402
rect 36924 20058 36952 20538
rect 36912 20052 36964 20058
rect 36912 19994 36964 20000
rect 36728 19984 36780 19990
rect 36728 19926 36780 19932
rect 36268 19508 36320 19514
rect 36320 19468 36492 19496
rect 36268 19450 36320 19456
rect 35992 19372 36044 19378
rect 35992 19314 36044 19320
rect 36004 18766 36032 19314
rect 36084 18896 36136 18902
rect 36082 18864 36084 18873
rect 36136 18864 36138 18873
rect 36082 18799 36138 18808
rect 36464 18766 36492 19468
rect 35992 18760 36044 18766
rect 35992 18702 36044 18708
rect 36452 18760 36504 18766
rect 36452 18702 36504 18708
rect 36636 18760 36688 18766
rect 36636 18702 36688 18708
rect 36360 18692 36412 18698
rect 36360 18634 36412 18640
rect 35808 17808 35860 17814
rect 35808 17750 35860 17756
rect 35624 17672 35676 17678
rect 35622 17640 35624 17649
rect 35808 17672 35860 17678
rect 35676 17640 35678 17649
rect 35808 17614 35860 17620
rect 35992 17672 36044 17678
rect 35992 17614 36044 17620
rect 35622 17575 35678 17584
rect 35072 17536 35124 17542
rect 35072 17478 35124 17484
rect 35532 17536 35584 17542
rect 35532 17478 35584 17484
rect 35084 17270 35112 17478
rect 35072 17264 35124 17270
rect 35072 17206 35124 17212
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35348 16040 35400 16046
rect 35348 15982 35400 15988
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34704 15496 34756 15502
rect 34704 15438 34756 15444
rect 34716 14890 34744 15438
rect 35360 15026 35388 15982
rect 35348 15020 35400 15026
rect 35348 14962 35400 14968
rect 34704 14884 34756 14890
rect 34704 14826 34756 14832
rect 34716 14482 34744 14826
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34704 14476 34756 14482
rect 34704 14418 34756 14424
rect 34796 14408 34848 14414
rect 34796 14350 34848 14356
rect 34808 13938 34836 14350
rect 34796 13932 34848 13938
rect 34796 13874 34848 13880
rect 34808 11762 34836 13874
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35440 13252 35492 13258
rect 35440 13194 35492 13200
rect 35452 12986 35480 13194
rect 35544 12986 35572 17478
rect 35820 17338 35848 17614
rect 36004 17542 36032 17614
rect 35992 17536 36044 17542
rect 35992 17478 36044 17484
rect 36268 17536 36320 17542
rect 36268 17478 36320 17484
rect 35808 17332 35860 17338
rect 35808 17274 35860 17280
rect 36280 16590 36308 17478
rect 36268 16584 36320 16590
rect 36268 16526 36320 16532
rect 35806 15464 35862 15473
rect 35806 15399 35862 15408
rect 35716 15020 35768 15026
rect 35716 14962 35768 14968
rect 35624 14952 35676 14958
rect 35624 14894 35676 14900
rect 35636 14226 35664 14894
rect 35728 14414 35756 14962
rect 35820 14958 35848 15399
rect 35808 14952 35860 14958
rect 35808 14894 35860 14900
rect 35820 14482 35848 14894
rect 35808 14476 35860 14482
rect 35808 14418 35860 14424
rect 35716 14408 35768 14414
rect 35716 14350 35768 14356
rect 35716 14272 35768 14278
rect 35636 14220 35716 14226
rect 35636 14214 35768 14220
rect 35636 14198 35756 14214
rect 35624 13864 35676 13870
rect 35624 13806 35676 13812
rect 35440 12980 35492 12986
rect 35440 12922 35492 12928
rect 35532 12980 35584 12986
rect 35532 12922 35584 12928
rect 35636 12918 35664 13806
rect 35624 12912 35676 12918
rect 35544 12860 35624 12866
rect 35544 12854 35676 12860
rect 35544 12838 35664 12854
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34796 11756 34848 11762
rect 34796 11698 34848 11704
rect 34704 10600 34756 10606
rect 34704 10542 34756 10548
rect 34716 9042 34744 10542
rect 34704 9036 34756 9042
rect 34704 8978 34756 8984
rect 34808 7886 34836 11698
rect 35440 11620 35492 11626
rect 35440 11562 35492 11568
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35348 11008 35400 11014
rect 35348 10950 35400 10956
rect 35360 10674 35388 10950
rect 35348 10668 35400 10674
rect 35348 10610 35400 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35348 9376 35400 9382
rect 35348 9318 35400 9324
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34980 8900 35032 8906
rect 34980 8842 35032 8848
rect 34992 8634 35020 8842
rect 34980 8628 35032 8634
rect 34980 8570 35032 8576
rect 35360 8498 35388 9318
rect 35348 8492 35400 8498
rect 35348 8434 35400 8440
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34796 7880 34848 7886
rect 34796 7822 34848 7828
rect 35256 7880 35308 7886
rect 35256 7822 35308 7828
rect 35268 7410 35296 7822
rect 35452 7818 35480 11562
rect 35544 8498 35572 12838
rect 35624 12776 35676 12782
rect 35624 12718 35676 12724
rect 35636 12442 35664 12718
rect 35624 12436 35676 12442
rect 35624 12378 35676 12384
rect 35728 11694 35756 14198
rect 35820 13530 35848 14418
rect 35992 13796 36044 13802
rect 35992 13738 36044 13744
rect 35900 13728 35952 13734
rect 35900 13670 35952 13676
rect 35808 13524 35860 13530
rect 35808 13466 35860 13472
rect 35912 12850 35940 13670
rect 35900 12844 35952 12850
rect 35900 12786 35952 12792
rect 36004 12782 36032 13738
rect 35992 12776 36044 12782
rect 35992 12718 36044 12724
rect 35808 11756 35860 11762
rect 35808 11698 35860 11704
rect 35716 11688 35768 11694
rect 35716 11630 35768 11636
rect 35624 11144 35676 11150
rect 35624 11086 35676 11092
rect 35636 10470 35664 11086
rect 35624 10464 35676 10470
rect 35624 10406 35676 10412
rect 35532 8492 35584 8498
rect 35532 8434 35584 8440
rect 35440 7812 35492 7818
rect 35440 7754 35492 7760
rect 35452 7478 35480 7754
rect 35440 7472 35492 7478
rect 35440 7414 35492 7420
rect 35256 7404 35308 7410
rect 35256 7346 35308 7352
rect 34796 7336 34848 7342
rect 34796 7278 34848 7284
rect 34704 6112 34756 6118
rect 34704 6054 34756 6060
rect 34716 5642 34744 6054
rect 34808 5710 34836 7278
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35544 6798 35572 8434
rect 35636 8430 35664 10406
rect 35820 9654 35848 11698
rect 36372 9654 36400 18634
rect 36544 17604 36596 17610
rect 36544 17546 36596 17552
rect 36556 14006 36584 17546
rect 36544 14000 36596 14006
rect 36544 13942 36596 13948
rect 36556 13530 36584 13942
rect 36544 13524 36596 13530
rect 36544 13466 36596 13472
rect 36452 12640 36504 12646
rect 36452 12582 36504 12588
rect 35808 9648 35860 9654
rect 35808 9590 35860 9596
rect 36360 9648 36412 9654
rect 36360 9590 36412 9596
rect 35820 9178 35848 9590
rect 36464 9586 36492 12582
rect 36648 11914 36676 18702
rect 36740 17882 36768 19926
rect 36912 19304 36964 19310
rect 36912 19246 36964 19252
rect 36728 17876 36780 17882
rect 36728 17818 36780 17824
rect 36924 15910 36952 19246
rect 36912 15904 36964 15910
rect 36912 15846 36964 15852
rect 36924 15706 36952 15846
rect 36912 15700 36964 15706
rect 36912 15642 36964 15648
rect 36728 14816 36780 14822
rect 36728 14758 36780 14764
rect 36740 13938 36768 14758
rect 36924 14414 36952 15642
rect 36912 14408 36964 14414
rect 36912 14350 36964 14356
rect 36728 13932 36780 13938
rect 36728 13874 36780 13880
rect 37016 12374 37044 22578
rect 37108 22094 37136 23446
rect 37280 22976 37332 22982
rect 37280 22918 37332 22924
rect 37292 22710 37320 22918
rect 37280 22704 37332 22710
rect 37280 22646 37332 22652
rect 38568 22704 38620 22710
rect 38568 22646 38620 22652
rect 38476 22636 38528 22642
rect 38476 22578 38528 22584
rect 37108 22066 37228 22094
rect 37200 22030 37228 22066
rect 37188 22024 37240 22030
rect 37188 21966 37240 21972
rect 37280 21412 37332 21418
rect 37280 21354 37332 21360
rect 37292 20602 37320 21354
rect 37832 21344 37884 21350
rect 37832 21286 37884 21292
rect 37280 20596 37332 20602
rect 37280 20538 37332 20544
rect 37844 20466 37872 21286
rect 37188 20460 37240 20466
rect 37188 20402 37240 20408
rect 37832 20460 37884 20466
rect 37832 20402 37884 20408
rect 37096 20392 37148 20398
rect 37096 20334 37148 20340
rect 37108 19786 37136 20334
rect 37200 19854 37228 20402
rect 37188 19848 37240 19854
rect 37188 19790 37240 19796
rect 37096 19780 37148 19786
rect 37096 19722 37148 19728
rect 37108 17610 37136 19722
rect 37200 17678 37228 19790
rect 37280 19372 37332 19378
rect 37280 19314 37332 19320
rect 37188 17672 37240 17678
rect 37188 17614 37240 17620
rect 37096 17604 37148 17610
rect 37096 17546 37148 17552
rect 37108 16182 37136 17546
rect 37096 16176 37148 16182
rect 37096 16118 37148 16124
rect 37200 16114 37228 17614
rect 37188 16108 37240 16114
rect 37188 16050 37240 16056
rect 37200 15570 37228 16050
rect 37188 15564 37240 15570
rect 37188 15506 37240 15512
rect 37188 14408 37240 14414
rect 37188 14350 37240 14356
rect 37096 13252 37148 13258
rect 37096 13194 37148 13200
rect 37108 12646 37136 13194
rect 37096 12640 37148 12646
rect 37096 12582 37148 12588
rect 37004 12368 37056 12374
rect 37004 12310 37056 12316
rect 36648 11886 36768 11914
rect 36636 11824 36688 11830
rect 36636 11766 36688 11772
rect 36648 11150 36676 11766
rect 36636 11144 36688 11150
rect 36636 11086 36688 11092
rect 36648 10810 36676 11086
rect 36636 10804 36688 10810
rect 36636 10746 36688 10752
rect 36452 9580 36504 9586
rect 36452 9522 36504 9528
rect 35808 9172 35860 9178
rect 35808 9114 35860 9120
rect 36464 8906 36492 9522
rect 36452 8900 36504 8906
rect 36452 8842 36504 8848
rect 35808 8560 35860 8566
rect 35808 8502 35860 8508
rect 35624 8424 35676 8430
rect 35624 8366 35676 8372
rect 35624 7404 35676 7410
rect 35624 7346 35676 7352
rect 35532 6792 35584 6798
rect 35532 6734 35584 6740
rect 35440 6656 35492 6662
rect 35440 6598 35492 6604
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34796 5704 34848 5710
rect 34796 5646 34848 5652
rect 34704 5636 34756 5642
rect 34704 5578 34756 5584
rect 34808 5370 34836 5646
rect 34796 5364 34848 5370
rect 34796 5306 34848 5312
rect 34808 4146 34836 5306
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 35452 4146 35480 6598
rect 35544 6322 35572 6734
rect 35532 6316 35584 6322
rect 35532 6258 35584 6264
rect 35532 5908 35584 5914
rect 35636 5896 35664 7346
rect 35820 6934 35848 8502
rect 36268 7880 36320 7886
rect 36268 7822 36320 7828
rect 35808 6928 35860 6934
rect 35808 6870 35860 6876
rect 35820 6390 35848 6870
rect 36280 6390 36308 7822
rect 36464 6390 36492 8842
rect 36740 8838 36768 11886
rect 37016 11354 37044 12310
rect 37004 11348 37056 11354
rect 37004 11290 37056 11296
rect 37200 10062 37228 14350
rect 37292 13190 37320 19314
rect 38488 18290 38516 22578
rect 38580 21350 38608 22646
rect 38948 22642 38976 24754
rect 39776 23322 39804 24754
rect 39856 24132 39908 24138
rect 39856 24074 39908 24080
rect 39764 23316 39816 23322
rect 39764 23258 39816 23264
rect 39868 23202 39896 24074
rect 39960 23866 39988 24754
rect 39948 23860 40000 23866
rect 39948 23802 40000 23808
rect 39776 23174 39896 23202
rect 38936 22636 38988 22642
rect 38936 22578 38988 22584
rect 39776 22574 39804 23174
rect 39764 22568 39816 22574
rect 39764 22510 39816 22516
rect 38568 21344 38620 21350
rect 38568 21286 38620 21292
rect 39776 20466 39804 22510
rect 40040 22024 40092 22030
rect 40040 21966 40092 21972
rect 39856 21888 39908 21894
rect 39856 21830 39908 21836
rect 39868 21622 39896 21830
rect 39856 21616 39908 21622
rect 39856 21558 39908 21564
rect 39948 21480 40000 21486
rect 39948 21422 40000 21428
rect 39580 20460 39632 20466
rect 39580 20402 39632 20408
rect 39764 20460 39816 20466
rect 39764 20402 39816 20408
rect 39592 20058 39620 20402
rect 39580 20052 39632 20058
rect 39580 19994 39632 20000
rect 38752 19848 38804 19854
rect 38752 19790 38804 19796
rect 38764 18426 38792 19790
rect 39672 19508 39724 19514
rect 39672 19450 39724 19456
rect 38752 18420 38804 18426
rect 38752 18362 38804 18368
rect 38476 18284 38528 18290
rect 38476 18226 38528 18232
rect 37648 18216 37700 18222
rect 37648 18158 37700 18164
rect 37372 17808 37424 17814
rect 37372 17750 37424 17756
rect 37384 16250 37412 17750
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37476 17202 37504 17614
rect 37660 17202 37688 18158
rect 38488 17610 38516 18226
rect 38764 17678 38792 18362
rect 38936 18284 38988 18290
rect 38936 18226 38988 18232
rect 38948 18086 38976 18226
rect 38936 18080 38988 18086
rect 38936 18022 38988 18028
rect 38752 17672 38804 17678
rect 38752 17614 38804 17620
rect 37832 17604 37884 17610
rect 37832 17546 37884 17552
rect 38476 17604 38528 17610
rect 38476 17546 38528 17552
rect 37464 17196 37516 17202
rect 37464 17138 37516 17144
rect 37648 17196 37700 17202
rect 37648 17138 37700 17144
rect 37476 16726 37504 17138
rect 37464 16720 37516 16726
rect 37464 16662 37516 16668
rect 37372 16244 37424 16250
rect 37372 16186 37424 16192
rect 37660 15502 37688 17138
rect 37844 15570 37872 17546
rect 38948 16794 38976 18022
rect 38108 16788 38160 16794
rect 38108 16730 38160 16736
rect 38200 16788 38252 16794
rect 38200 16730 38252 16736
rect 38936 16788 38988 16794
rect 38936 16730 38988 16736
rect 37832 15564 37884 15570
rect 37832 15506 37884 15512
rect 37648 15496 37700 15502
rect 37648 15438 37700 15444
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 37476 14074 37504 14962
rect 37660 14278 37688 15438
rect 37844 15162 37872 15506
rect 37832 15156 37884 15162
rect 37832 15098 37884 15104
rect 38120 14958 38148 16730
rect 38212 15502 38240 16730
rect 38660 16108 38712 16114
rect 38660 16050 38712 16056
rect 38200 15496 38252 15502
rect 38200 15438 38252 15444
rect 38672 15366 38700 16050
rect 38752 15972 38804 15978
rect 38752 15914 38804 15920
rect 38764 15502 38792 15914
rect 38936 15904 38988 15910
rect 38936 15846 38988 15852
rect 38752 15496 38804 15502
rect 38752 15438 38804 15444
rect 38660 15360 38712 15366
rect 38660 15302 38712 15308
rect 38672 15162 38700 15302
rect 38568 15156 38620 15162
rect 38568 15098 38620 15104
rect 38660 15156 38712 15162
rect 38660 15098 38712 15104
rect 38108 14952 38160 14958
rect 38108 14894 38160 14900
rect 38120 14278 38148 14894
rect 37648 14272 37700 14278
rect 37648 14214 37700 14220
rect 38108 14272 38160 14278
rect 38108 14214 38160 14220
rect 37464 14068 37516 14074
rect 37464 14010 37516 14016
rect 37280 13184 37332 13190
rect 37280 13126 37332 13132
rect 37292 12986 37320 13126
rect 37280 12980 37332 12986
rect 37280 12922 37332 12928
rect 37660 12850 37688 14214
rect 38120 13326 38148 14214
rect 38580 13938 38608 15098
rect 38764 15026 38792 15438
rect 38844 15360 38896 15366
rect 38844 15302 38896 15308
rect 38856 15094 38884 15302
rect 38844 15088 38896 15094
rect 38844 15030 38896 15036
rect 38752 15020 38804 15026
rect 38752 14962 38804 14968
rect 38948 14414 38976 15846
rect 39580 15632 39632 15638
rect 39580 15574 39632 15580
rect 38936 14408 38988 14414
rect 38936 14350 38988 14356
rect 39488 14340 39540 14346
rect 39488 14282 39540 14288
rect 38568 13932 38620 13938
rect 38568 13874 38620 13880
rect 39500 13870 39528 14282
rect 38384 13864 38436 13870
rect 38384 13806 38436 13812
rect 39488 13864 39540 13870
rect 39488 13806 39540 13812
rect 38396 13462 38424 13806
rect 39304 13728 39356 13734
rect 39304 13670 39356 13676
rect 38384 13456 38436 13462
rect 38384 13398 38436 13404
rect 38108 13320 38160 13326
rect 38108 13262 38160 13268
rect 38120 12850 38148 13262
rect 37648 12844 37700 12850
rect 37648 12786 37700 12792
rect 38108 12844 38160 12850
rect 38108 12786 38160 12792
rect 38292 12232 38344 12238
rect 38292 12174 38344 12180
rect 38304 11830 38332 12174
rect 38292 11824 38344 11830
rect 38292 11766 38344 11772
rect 38108 11348 38160 11354
rect 38108 11290 38160 11296
rect 37556 11076 37608 11082
rect 37556 11018 37608 11024
rect 37188 10056 37240 10062
rect 37188 9998 37240 10004
rect 37568 9654 37596 11018
rect 38120 11014 38148 11290
rect 38304 11082 38332 11766
rect 38292 11076 38344 11082
rect 38292 11018 38344 11024
rect 38108 11008 38160 11014
rect 38108 10950 38160 10956
rect 38120 10810 38148 10950
rect 38108 10804 38160 10810
rect 38108 10746 38160 10752
rect 37740 10668 37792 10674
rect 37740 10610 37792 10616
rect 37556 9648 37608 9654
rect 37556 9590 37608 9596
rect 37568 8922 37596 9590
rect 37568 8894 37688 8922
rect 36728 8832 36780 8838
rect 36728 8774 36780 8780
rect 37556 8832 37608 8838
rect 37556 8774 37608 8780
rect 37568 8498 37596 8774
rect 37556 8492 37608 8498
rect 37556 8434 37608 8440
rect 37096 7744 37148 7750
rect 37096 7686 37148 7692
rect 37108 6914 37136 7686
rect 37660 7478 37688 8894
rect 37752 8498 37780 10610
rect 37924 9512 37976 9518
rect 37924 9454 37976 9460
rect 37936 8974 37964 9454
rect 37924 8968 37976 8974
rect 37924 8910 37976 8916
rect 37740 8492 37792 8498
rect 37740 8434 37792 8440
rect 37752 8090 37780 8434
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 37648 7472 37700 7478
rect 37648 7414 37700 7420
rect 37108 6886 37228 6914
rect 36820 6792 36872 6798
rect 36820 6734 36872 6740
rect 37004 6792 37056 6798
rect 37004 6734 37056 6740
rect 36832 6458 36860 6734
rect 36820 6452 36872 6458
rect 36820 6394 36872 6400
rect 35808 6384 35860 6390
rect 35808 6326 35860 6332
rect 36268 6384 36320 6390
rect 36268 6326 36320 6332
rect 36452 6384 36504 6390
rect 36452 6326 36504 6332
rect 36280 5914 36308 6326
rect 37016 6186 37044 6734
rect 37200 6322 37228 6886
rect 37556 6656 37608 6662
rect 37556 6598 37608 6604
rect 37188 6316 37240 6322
rect 37188 6258 37240 6264
rect 37004 6180 37056 6186
rect 37004 6122 37056 6128
rect 37200 5914 37228 6258
rect 35584 5868 35664 5896
rect 35532 5850 35584 5856
rect 34796 4140 34848 4146
rect 34796 4082 34848 4088
rect 35440 4140 35492 4146
rect 35440 4082 35492 4088
rect 35636 3942 35664 5868
rect 36268 5908 36320 5914
rect 36268 5850 36320 5856
rect 37188 5908 37240 5914
rect 37188 5850 37240 5856
rect 37568 5710 37596 6598
rect 37660 6390 37688 7414
rect 37648 6384 37700 6390
rect 37648 6326 37700 6332
rect 37936 6322 37964 8910
rect 38016 8900 38068 8906
rect 38016 8842 38068 8848
rect 38028 8634 38056 8842
rect 38016 8628 38068 8634
rect 38016 8570 38068 8576
rect 38120 7546 38148 10746
rect 38396 8566 38424 13398
rect 38568 13320 38620 13326
rect 38568 13262 38620 13268
rect 38580 12374 38608 13262
rect 39316 13258 39344 13670
rect 39304 13252 39356 13258
rect 39304 13194 39356 13200
rect 38844 13184 38896 13190
rect 38844 13126 38896 13132
rect 38856 12918 38884 13126
rect 38844 12912 38896 12918
rect 38844 12854 38896 12860
rect 38568 12368 38620 12374
rect 38568 12310 38620 12316
rect 38580 11778 38608 12310
rect 39028 12300 39080 12306
rect 39028 12242 39080 12248
rect 38488 11750 38608 11778
rect 38660 11756 38712 11762
rect 38488 11150 38516 11750
rect 38660 11698 38712 11704
rect 38568 11688 38620 11694
rect 38568 11630 38620 11636
rect 38476 11144 38528 11150
rect 38476 11086 38528 11092
rect 38580 10742 38608 11630
rect 38672 11354 38700 11698
rect 38660 11348 38712 11354
rect 38660 11290 38712 11296
rect 39040 11286 39068 12242
rect 39500 12238 39528 13806
rect 39592 12850 39620 15574
rect 39684 14226 39712 19450
rect 39776 18698 39804 20402
rect 39960 20398 39988 21422
rect 39948 20392 40000 20398
rect 39948 20334 40000 20340
rect 39960 19310 39988 20334
rect 40052 19854 40080 21966
rect 40236 21894 40264 25434
rect 40420 25226 40448 26182
rect 40788 25906 40816 26182
rect 40592 25900 40644 25906
rect 40592 25842 40644 25848
rect 40776 25900 40828 25906
rect 40776 25842 40828 25848
rect 40500 25832 40552 25838
rect 40500 25774 40552 25780
rect 40408 25220 40460 25226
rect 40408 25162 40460 25168
rect 40512 25158 40540 25774
rect 40604 25702 40632 25842
rect 40592 25696 40644 25702
rect 40592 25638 40644 25644
rect 40500 25152 40552 25158
rect 40500 25094 40552 25100
rect 40408 24064 40460 24070
rect 40408 24006 40460 24012
rect 40420 23118 40448 24006
rect 40408 23112 40460 23118
rect 40408 23054 40460 23060
rect 40408 22976 40460 22982
rect 40408 22918 40460 22924
rect 40420 22506 40448 22918
rect 40408 22500 40460 22506
rect 40408 22442 40460 22448
rect 40316 22432 40368 22438
rect 40316 22374 40368 22380
rect 40328 22027 40356 22374
rect 40316 22021 40368 22027
rect 40316 21963 40368 21969
rect 40224 21888 40276 21894
rect 40224 21830 40276 21836
rect 40420 19922 40448 22442
rect 40512 22030 40540 25094
rect 40684 23656 40736 23662
rect 40684 23598 40736 23604
rect 40696 23050 40724 23598
rect 40788 23254 40816 25842
rect 40868 25152 40920 25158
rect 40868 25094 40920 25100
rect 40880 24954 40908 25094
rect 40868 24948 40920 24954
rect 40868 24890 40920 24896
rect 40880 23730 40908 24890
rect 41052 24200 41104 24206
rect 41052 24142 41104 24148
rect 40868 23724 40920 23730
rect 40868 23666 40920 23672
rect 40880 23322 40908 23666
rect 41064 23526 41092 24142
rect 41144 24064 41196 24070
rect 41144 24006 41196 24012
rect 41156 23730 41184 24006
rect 41144 23724 41196 23730
rect 41144 23666 41196 23672
rect 41236 23724 41288 23730
rect 41236 23666 41288 23672
rect 41052 23520 41104 23526
rect 41052 23462 41104 23468
rect 40868 23316 40920 23322
rect 40868 23258 40920 23264
rect 40776 23248 40828 23254
rect 41248 23202 41276 23666
rect 40776 23190 40828 23196
rect 41156 23174 41276 23202
rect 41156 23118 41184 23174
rect 41144 23112 41196 23118
rect 41144 23054 41196 23060
rect 40684 23044 40736 23050
rect 40684 22986 40736 22992
rect 40500 22024 40552 22030
rect 40500 21966 40552 21972
rect 40408 19916 40460 19922
rect 40408 19858 40460 19864
rect 40040 19848 40092 19854
rect 40040 19790 40092 19796
rect 40052 19718 40080 19790
rect 40040 19712 40092 19718
rect 40040 19654 40092 19660
rect 40408 19372 40460 19378
rect 40408 19314 40460 19320
rect 39948 19304 40000 19310
rect 39948 19246 40000 19252
rect 39764 18692 39816 18698
rect 39764 18634 39816 18640
rect 39776 17202 39804 18634
rect 39960 18086 39988 19246
rect 40420 18970 40448 19314
rect 40408 18964 40460 18970
rect 40408 18906 40460 18912
rect 40512 18850 40540 21966
rect 40960 21888 41012 21894
rect 40960 21830 41012 21836
rect 40684 20256 40736 20262
rect 40684 20198 40736 20204
rect 40696 19854 40724 20198
rect 40776 19916 40828 19922
rect 40776 19858 40828 19864
rect 40684 19848 40736 19854
rect 40684 19790 40736 19796
rect 40420 18822 40540 18850
rect 39948 18080 40000 18086
rect 39948 18022 40000 18028
rect 39960 17270 39988 18022
rect 39948 17264 40000 17270
rect 39948 17206 40000 17212
rect 39764 17196 39816 17202
rect 39764 17138 39816 17144
rect 39856 17128 39908 17134
rect 39856 17070 39908 17076
rect 39868 14346 39896 17070
rect 39960 16250 39988 17206
rect 39948 16244 40000 16250
rect 39948 16186 40000 16192
rect 40132 16108 40184 16114
rect 40132 16050 40184 16056
rect 40144 15706 40172 16050
rect 40132 15700 40184 15706
rect 40132 15642 40184 15648
rect 39856 14340 39908 14346
rect 39856 14282 39908 14288
rect 39684 14198 39896 14226
rect 39580 12844 39632 12850
rect 39580 12786 39632 12792
rect 39592 12434 39620 12786
rect 39592 12406 39804 12434
rect 39776 12238 39804 12406
rect 39488 12232 39540 12238
rect 39488 12174 39540 12180
rect 39764 12232 39816 12238
rect 39764 12174 39816 12180
rect 39868 11898 39896 14198
rect 40420 13870 40448 18822
rect 40788 18766 40816 19858
rect 40500 18760 40552 18766
rect 40500 18702 40552 18708
rect 40776 18760 40828 18766
rect 40776 18702 40828 18708
rect 40512 18290 40540 18702
rect 40500 18284 40552 18290
rect 40500 18226 40552 18232
rect 40512 17746 40540 18226
rect 40500 17740 40552 17746
rect 40500 17682 40552 17688
rect 40788 16794 40816 18702
rect 40972 18290 41000 21830
rect 41156 19854 41184 23054
rect 41144 19848 41196 19854
rect 41144 19790 41196 19796
rect 41156 18766 41184 19790
rect 41696 19780 41748 19786
rect 41696 19722 41748 19728
rect 41708 19514 41736 19722
rect 41696 19508 41748 19514
rect 41696 19450 41748 19456
rect 41708 18766 41736 19450
rect 41144 18760 41196 18766
rect 41144 18702 41196 18708
rect 41696 18760 41748 18766
rect 41696 18702 41748 18708
rect 40960 18284 41012 18290
rect 40960 18226 41012 18232
rect 41052 18284 41104 18290
rect 41052 18226 41104 18232
rect 40868 18148 40920 18154
rect 40868 18090 40920 18096
rect 40776 16788 40828 16794
rect 40776 16730 40828 16736
rect 40500 16516 40552 16522
rect 40500 16458 40552 16464
rect 40512 15638 40540 16458
rect 40500 15632 40552 15638
rect 40500 15574 40552 15580
rect 40684 15496 40736 15502
rect 40684 15438 40736 15444
rect 40696 14414 40724 15438
rect 40880 14550 40908 18090
rect 40972 17814 41000 18226
rect 41064 17882 41092 18226
rect 41052 17876 41104 17882
rect 41052 17818 41104 17824
rect 40960 17808 41012 17814
rect 40960 17750 41012 17756
rect 41156 15502 41184 18702
rect 41144 15496 41196 15502
rect 41144 15438 41196 15444
rect 41328 15496 41380 15502
rect 41328 15438 41380 15444
rect 41512 15496 41564 15502
rect 41512 15438 41564 15444
rect 41340 14618 41368 15438
rect 41524 15026 41552 15438
rect 41512 15020 41564 15026
rect 41512 14962 41564 14968
rect 41328 14612 41380 14618
rect 41328 14554 41380 14560
rect 40868 14544 40920 14550
rect 40868 14486 40920 14492
rect 40684 14408 40736 14414
rect 40684 14350 40736 14356
rect 40696 14006 40724 14350
rect 40684 14000 40736 14006
rect 40684 13942 40736 13948
rect 40408 13864 40460 13870
rect 40408 13806 40460 13812
rect 39856 11892 39908 11898
rect 39856 11834 39908 11840
rect 40776 11552 40828 11558
rect 40776 11494 40828 11500
rect 39028 11280 39080 11286
rect 39028 11222 39080 11228
rect 38568 10736 38620 10742
rect 38568 10678 38620 10684
rect 38580 10266 38608 10678
rect 39040 10606 39068 11222
rect 40788 11218 40816 11494
rect 40776 11212 40828 11218
rect 40776 11154 40828 11160
rect 39396 10668 39448 10674
rect 39396 10610 39448 10616
rect 39028 10600 39080 10606
rect 39028 10542 39080 10548
rect 38936 10464 38988 10470
rect 38936 10406 38988 10412
rect 38568 10260 38620 10266
rect 38568 10202 38620 10208
rect 38948 9654 38976 10406
rect 38936 9648 38988 9654
rect 38936 9590 38988 9596
rect 38384 8560 38436 8566
rect 38384 8502 38436 8508
rect 38108 7540 38160 7546
rect 38108 7482 38160 7488
rect 38120 6730 38148 7482
rect 38844 7200 38896 7206
rect 38844 7142 38896 7148
rect 38568 6996 38620 7002
rect 38568 6938 38620 6944
rect 38752 6996 38804 7002
rect 38752 6938 38804 6944
rect 38580 6798 38608 6938
rect 38568 6792 38620 6798
rect 38764 6746 38792 6938
rect 38856 6798 38884 7142
rect 39040 6934 39068 10542
rect 39408 9722 39436 10610
rect 39396 9716 39448 9722
rect 39396 9658 39448 9664
rect 39672 7336 39724 7342
rect 39672 7278 39724 7284
rect 39028 6928 39080 6934
rect 39028 6870 39080 6876
rect 38620 6740 38792 6746
rect 38568 6734 38792 6740
rect 38844 6792 38896 6798
rect 39040 6746 39068 6870
rect 38844 6734 38896 6740
rect 38108 6724 38160 6730
rect 38108 6666 38160 6672
rect 38580 6718 38792 6734
rect 38948 6730 39068 6746
rect 38936 6724 39068 6730
rect 38580 6669 38608 6718
rect 38988 6718 39068 6724
rect 38936 6666 38988 6672
rect 38384 6656 38436 6662
rect 38384 6598 38436 6604
rect 38396 6390 38424 6598
rect 39684 6458 39712 7278
rect 39672 6452 39724 6458
rect 39672 6394 39724 6400
rect 38384 6384 38436 6390
rect 38384 6326 38436 6332
rect 37924 6316 37976 6322
rect 37924 6258 37976 6264
rect 37556 5704 37608 5710
rect 37556 5646 37608 5652
rect 42076 4826 42104 56102
rect 42064 4820 42116 4826
rect 42064 4762 42116 4768
rect 35624 3936 35676 3942
rect 35624 3878 35676 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 35348 3528 35400 3534
rect 35348 3470 35400 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 36636 3528 36688 3534
rect 36636 3470 36688 3476
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 38568 3528 38620 3534
rect 38568 3470 38620 3476
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 40500 3528 40552 3534
rect 40500 3470 40552 3476
rect 41052 3528 41104 3534
rect 41052 3470 41104 3476
rect 42432 3528 42484 3534
rect 42432 3470 42484 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 44364 3528 44416 3534
rect 44364 3470 44416 3476
rect 45192 3528 45244 3534
rect 45192 3470 45244 3476
rect 34612 2100 34664 2106
rect 34612 2042 34664 2048
rect 34716 800 34744 3470
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 1850 35388 3470
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 34992 1822 35388 1850
rect 34992 800 35020 1822
rect 35452 1442 35480 2790
rect 35532 2508 35584 2514
rect 35532 2450 35584 2456
rect 35268 1414 35480 1442
rect 35268 800 35296 1414
rect 35544 800 35572 2450
rect 35820 800 35848 3470
rect 36360 2848 36412 2854
rect 36360 2790 36412 2796
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 36096 800 36124 2382
rect 36372 800 36400 2790
rect 36648 800 36676 3470
rect 37188 2916 37240 2922
rect 37188 2858 37240 2864
rect 36912 2372 36964 2378
rect 36912 2314 36964 2320
rect 36924 800 36952 2314
rect 37200 800 37228 2858
rect 37476 800 37504 3470
rect 38292 2984 38344 2990
rect 38292 2926 38344 2932
rect 37740 2848 37792 2854
rect 37740 2790 37792 2796
rect 37752 800 37780 2790
rect 38016 2576 38068 2582
rect 38016 2518 38068 2524
rect 38028 800 38056 2518
rect 38304 800 38332 2926
rect 38580 800 38608 3470
rect 39120 2916 39172 2922
rect 39120 2858 39172 2864
rect 38844 2508 38896 2514
rect 38844 2450 38896 2456
rect 38856 800 38884 2450
rect 39132 800 39160 2858
rect 39672 2848 39724 2854
rect 39672 2790 39724 2796
rect 39396 2440 39448 2446
rect 39396 2382 39448 2388
rect 39408 800 39436 2382
rect 39684 800 39712 2790
rect 39960 800 39988 3470
rect 40224 2916 40276 2922
rect 40224 2858 40276 2864
rect 40236 800 40264 2858
rect 40512 800 40540 3470
rect 40776 2508 40828 2514
rect 40776 2450 40828 2456
rect 40788 800 40816 2450
rect 41064 800 41092 3470
rect 42156 2984 42208 2990
rect 42156 2926 42208 2932
rect 41604 2848 41656 2854
rect 41604 2790 41656 2796
rect 41328 2440 41380 2446
rect 41328 2382 41380 2388
rect 41340 800 41368 2382
rect 41616 800 41644 2790
rect 41880 2576 41932 2582
rect 41880 2518 41932 2524
rect 41892 800 41920 2518
rect 42168 800 42196 2926
rect 42444 800 42472 3470
rect 42720 800 42748 3470
rect 42984 2916 43036 2922
rect 42984 2858 43036 2864
rect 44088 2916 44140 2922
rect 44088 2858 44140 2864
rect 42996 800 43024 2858
rect 43536 2848 43588 2854
rect 43536 2790 43588 2796
rect 43260 2508 43312 2514
rect 43260 2450 43312 2456
rect 43272 800 43300 2450
rect 43548 800 43576 2790
rect 43812 2440 43864 2446
rect 43812 2382 43864 2388
rect 43824 800 43852 2382
rect 44100 800 44128 2858
rect 44376 800 44404 3470
rect 44916 2848 44968 2854
rect 44916 2790 44968 2796
rect 44640 2372 44692 2378
rect 44640 2314 44692 2320
rect 44652 800 44680 2314
rect 44928 800 44956 2790
rect 45204 800 45232 3470
rect 45468 2848 45520 2854
rect 45468 2790 45520 2796
rect 45480 800 45508 2790
rect 45572 2038 45600 56306
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 58162 55176 58218 55185
rect 58162 55111 58164 55120
rect 58216 55111 58218 55120
rect 58164 55082 58216 55088
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 57888 53984 57940 53990
rect 57888 53926 57940 53932
rect 57900 53825 57928 53926
rect 57886 53816 57942 53825
rect 57886 53751 57942 53760
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 57888 52488 57940 52494
rect 57886 52456 57888 52465
rect 57940 52456 57942 52465
rect 57886 52391 57942 52400
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 58164 51400 58216 51406
rect 58164 51342 58216 51348
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 58176 51105 58204 51342
rect 58162 51096 58218 51105
rect 58162 51031 58218 51040
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 58164 49768 58216 49774
rect 58162 49736 58164 49745
rect 58216 49736 58218 49745
rect 58162 49671 58218 49680
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 58164 48544 58216 48550
rect 58164 48486 58216 48492
rect 58176 48385 58204 48486
rect 58162 48376 58218 48385
rect 58162 48311 58218 48320
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 58164 47048 58216 47054
rect 58162 47016 58164 47025
rect 58216 47016 58218 47025
rect 58162 46951 58218 46960
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 58164 45960 58216 45966
rect 58164 45902 58216 45908
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 58176 45665 58204 45902
rect 58162 45656 58218 45665
rect 58162 45591 58218 45600
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 58162 44296 58218 44305
rect 58162 44231 58164 44240
rect 58216 44231 58218 44240
rect 58164 44202 58216 44208
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 58164 43104 58216 43110
rect 58164 43046 58216 43052
rect 58176 42945 58204 43046
rect 58162 42936 58218 42945
rect 58162 42871 58218 42880
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 58164 41608 58216 41614
rect 58162 41576 58164 41585
rect 58216 41576 58218 41585
rect 58162 41511 58218 41520
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 58164 40520 58216 40526
rect 58164 40462 58216 40468
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 58176 40225 58204 40462
rect 58162 40216 58218 40225
rect 58162 40151 58218 40160
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 58162 38856 58218 38865
rect 58162 38791 58164 38800
rect 58216 38791 58218 38800
rect 58164 38762 58216 38768
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 58164 37664 58216 37670
rect 58164 37606 58216 37612
rect 58176 37505 58204 37606
rect 58162 37496 58218 37505
rect 58162 37431 58218 37440
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 58164 36168 58216 36174
rect 58162 36136 58164 36145
rect 58216 36136 58218 36145
rect 58162 36071 58218 36080
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 58164 35080 58216 35086
rect 58164 35022 58216 35028
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 58176 34785 58204 35022
rect 58162 34776 58218 34785
rect 58162 34711 58218 34720
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 58162 33416 58218 33425
rect 58162 33351 58164 33360
rect 58216 33351 58218 33360
rect 58164 33322 58216 33328
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 58164 32224 58216 32230
rect 58164 32166 58216 32172
rect 58176 32065 58204 32166
rect 58162 32056 58218 32065
rect 58162 31991 58218 32000
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 58164 30728 58216 30734
rect 58162 30696 58164 30705
rect 58216 30696 58218 30705
rect 58162 30631 58218 30640
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 58164 29640 58216 29646
rect 58164 29582 58216 29588
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 58176 29345 58204 29582
rect 58162 29336 58218 29345
rect 58162 29271 58218 29280
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 58162 27976 58218 27985
rect 58162 27911 58164 27920
rect 58216 27911 58218 27920
rect 58164 27882 58216 27888
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 58164 26784 58216 26790
rect 58164 26726 58216 26732
rect 58176 26625 58204 26726
rect 58162 26616 58218 26625
rect 58162 26551 58218 26560
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 58164 25288 58216 25294
rect 58162 25256 58164 25265
rect 58216 25256 58218 25265
rect 58162 25191 58218 25200
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 58164 24200 58216 24206
rect 58164 24142 58216 24148
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 58176 23905 58204 24142
rect 58162 23896 58218 23905
rect 58162 23831 58218 23840
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 58162 22536 58218 22545
rect 58162 22471 58164 22480
rect 58216 22471 58218 22480
rect 58164 22442 58216 22448
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 58164 21344 58216 21350
rect 58164 21286 58216 21292
rect 58176 21185 58204 21286
rect 58162 21176 58218 21185
rect 58162 21111 58218 21120
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 58164 19848 58216 19854
rect 58162 19816 58164 19825
rect 58216 19816 58218 19825
rect 58162 19751 58218 19760
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 58164 18760 58216 18766
rect 58164 18702 58216 18708
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 58176 18465 58204 18702
rect 58162 18456 58218 18465
rect 58162 18391 58218 18400
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 58162 17096 58218 17105
rect 58162 17031 58164 17040
rect 58216 17031 58218 17040
rect 58164 17002 58216 17008
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 58164 15904 58216 15910
rect 58164 15846 58216 15852
rect 58176 15745 58204 15846
rect 58162 15736 58218 15745
rect 58162 15671 58218 15680
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 58164 14408 58216 14414
rect 58162 14376 58164 14385
rect 58216 14376 58218 14385
rect 58162 14311 58218 14320
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 58164 13320 58216 13326
rect 58164 13262 58216 13268
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 58176 13025 58204 13262
rect 58162 13016 58218 13025
rect 58162 12951 58218 12960
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 58162 11656 58218 11665
rect 58162 11591 58164 11600
rect 58216 11591 58218 11600
rect 58164 11562 58216 11568
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 58164 10464 58216 10470
rect 58164 10406 58216 10412
rect 58176 10305 58204 10406
rect 58162 10296 58218 10305
rect 58162 10231 58218 10240
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 58164 8968 58216 8974
rect 58162 8936 58164 8945
rect 58216 8936 58218 8945
rect 58162 8871 58218 8880
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 58164 7880 58216 7886
rect 58164 7822 58216 7828
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 58176 7585 58204 7822
rect 58162 7576 58218 7585
rect 58162 7511 58218 7520
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 58162 6216 58218 6225
rect 58162 6151 58164 6160
rect 58216 6151 58218 6160
rect 58164 6122 58216 6128
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 53748 5160 53800 5166
rect 53748 5102 53800 5108
rect 53656 5024 53708 5030
rect 53656 4966 53708 4972
rect 52184 4752 52236 4758
rect 52184 4694 52236 4700
rect 52092 4616 52144 4622
rect 52092 4558 52144 4564
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 51816 4072 51868 4078
rect 51816 4014 51868 4020
rect 51080 3936 51132 3942
rect 51080 3878 51132 3884
rect 51356 3936 51408 3942
rect 51356 3878 51408 3884
rect 46296 3664 46348 3670
rect 46296 3606 46348 3612
rect 46020 3528 46072 3534
rect 46020 3470 46072 3476
rect 45744 2576 45796 2582
rect 45744 2518 45796 2524
rect 45560 2032 45612 2038
rect 45560 1974 45612 1980
rect 45756 800 45784 2518
rect 46032 800 46060 3470
rect 46308 800 46336 3606
rect 50804 3596 50856 3602
rect 50804 3538 50856 3544
rect 47676 3528 47728 3534
rect 47676 3470 47728 3476
rect 48228 3528 48280 3534
rect 48228 3470 48280 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50620 3528 50672 3534
rect 50620 3470 50672 3476
rect 47400 2916 47452 2922
rect 47400 2858 47452 2864
rect 46848 2848 46900 2854
rect 46848 2790 46900 2796
rect 46572 2508 46624 2514
rect 46572 2450 46624 2456
rect 46584 800 46612 2450
rect 46860 800 46888 2790
rect 47124 2440 47176 2446
rect 47124 2382 47176 2388
rect 47136 800 47164 2382
rect 47412 800 47440 2858
rect 47688 800 47716 3470
rect 47952 2848 48004 2854
rect 47952 2790 48004 2796
rect 47964 800 47992 2790
rect 48240 800 48268 3470
rect 48780 2916 48832 2922
rect 48780 2858 48832 2864
rect 49884 2916 49936 2922
rect 49884 2858 49936 2864
rect 48504 2508 48556 2514
rect 48504 2450 48556 2456
rect 48516 800 48544 2450
rect 48792 800 48820 2858
rect 49332 2848 49384 2854
rect 49332 2790 49384 2796
rect 49056 2440 49108 2446
rect 49056 2382 49108 2388
rect 49068 800 49096 2382
rect 49344 800 49372 2790
rect 49608 2576 49660 2582
rect 49608 2518 49660 2524
rect 49620 800 49648 2518
rect 49896 800 49924 2858
rect 50172 800 50200 3470
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50632 1850 50660 3470
rect 50712 2848 50764 2854
rect 50712 2790 50764 2796
rect 50448 1822 50660 1850
rect 50448 800 50476 1822
rect 50724 1442 50752 2790
rect 50632 1414 50752 1442
rect 50632 800 50660 1414
rect 50816 1306 50844 3538
rect 50988 2916 51040 2922
rect 50988 2858 51040 2864
rect 50896 2440 50948 2446
rect 50896 2382 50948 2388
rect 50724 1278 50844 1306
rect 50724 800 50752 1278
rect 50908 1170 50936 2382
rect 50816 1142 50936 1170
rect 50816 800 50844 1142
rect 51000 1034 51028 2858
rect 50908 1006 51028 1034
rect 50908 800 50936 1006
rect 50988 944 51040 950
rect 50988 886 51040 892
rect 51000 800 51028 886
rect 51092 800 51120 3878
rect 51172 3528 51224 3534
rect 51172 3470 51224 3476
rect 51184 800 51212 3470
rect 51264 2304 51316 2310
rect 51264 2246 51316 2252
rect 51276 800 51304 2246
rect 51368 800 51396 3878
rect 51448 3664 51500 3670
rect 51448 3606 51500 3612
rect 51460 800 51488 3606
rect 51632 3596 51684 3602
rect 51632 3538 51684 3544
rect 51540 2848 51592 2854
rect 51540 2790 51592 2796
rect 51552 800 51580 2790
rect 51644 800 51672 3538
rect 51724 3052 51776 3058
rect 51724 2994 51776 3000
rect 51736 800 51764 2994
rect 51828 800 51856 4014
rect 51908 3120 51960 3126
rect 51908 3062 51960 3068
rect 51920 800 51948 3062
rect 52000 2644 52052 2650
rect 52000 2586 52052 2592
rect 52012 800 52040 2586
rect 52104 800 52132 4558
rect 52196 800 52224 4694
rect 53196 4684 53248 4690
rect 53196 4626 53248 4632
rect 52644 4616 52696 4622
rect 52644 4558 52696 4564
rect 52460 3936 52512 3942
rect 52460 3878 52512 3884
rect 52276 3528 52328 3534
rect 52276 3470 52328 3476
rect 52288 800 52316 3470
rect 52368 2100 52420 2106
rect 52368 2042 52420 2048
rect 52380 800 52408 2042
rect 52472 800 52500 3878
rect 52552 2440 52604 2446
rect 52552 2382 52604 2388
rect 52564 1154 52592 2382
rect 52552 1148 52604 1154
rect 52552 1090 52604 1096
rect 52552 944 52604 950
rect 52552 886 52604 892
rect 52564 800 52592 886
rect 52656 800 52684 4558
rect 53012 4140 53064 4146
rect 53012 4082 53064 4088
rect 52828 4004 52880 4010
rect 52828 3946 52880 3952
rect 52736 3732 52788 3738
rect 52736 3674 52788 3680
rect 52748 1426 52776 3674
rect 52736 1420 52788 1426
rect 52736 1362 52788 1368
rect 52840 1170 52868 3946
rect 53024 2774 53052 4082
rect 53104 2984 53156 2990
rect 53104 2926 53156 2932
rect 52748 1142 52868 1170
rect 52932 2746 53052 2774
rect 52748 800 52776 1142
rect 52932 1034 52960 2746
rect 53012 1420 53064 1426
rect 53012 1362 53064 1368
rect 52840 1006 52960 1034
rect 52840 800 52868 1006
rect 52920 944 52972 950
rect 52920 886 52972 892
rect 52932 800 52960 886
rect 53024 800 53052 1362
rect 53116 800 53144 2926
rect 53208 800 53236 4626
rect 53288 3460 53340 3466
rect 53288 3402 53340 3408
rect 53300 800 53328 3402
rect 53378 2952 53434 2961
rect 53378 2887 53434 2896
rect 53392 800 53420 2887
rect 53470 2816 53526 2825
rect 53470 2751 53526 2760
rect 53484 800 53512 2751
rect 53564 2032 53616 2038
rect 53564 1974 53616 1980
rect 53576 800 53604 1974
rect 53668 800 53696 4966
rect 53760 800 53788 5102
rect 54116 5092 54168 5098
rect 54116 5034 54168 5040
rect 53932 4752 53984 4758
rect 53932 4694 53984 4700
rect 53840 3596 53892 3602
rect 53840 3538 53892 3544
rect 53852 800 53880 3538
rect 53944 800 53972 4694
rect 54024 4072 54076 4078
rect 54024 4014 54076 4020
rect 54036 800 54064 4014
rect 54128 800 54156 5034
rect 58164 5024 58216 5030
rect 58164 4966 58216 4972
rect 58176 4865 58204 4966
rect 58162 4856 58218 4865
rect 58162 4791 58218 4800
rect 54300 4684 54352 4690
rect 54300 4626 54352 4632
rect 54208 2916 54260 2922
rect 54208 2858 54260 2864
rect 54220 800 54248 2858
rect 54312 800 54340 4626
rect 55312 3936 55364 3942
rect 55312 3878 55364 3884
rect 58440 3936 58492 3942
rect 58440 3878 58492 3884
rect 54760 3052 54812 3058
rect 54760 2994 54812 3000
rect 54772 882 54800 2994
rect 55324 2825 55352 3878
rect 57520 3528 57572 3534
rect 58164 3528 58216 3534
rect 57520 3470 57572 3476
rect 58162 3496 58164 3505
rect 58216 3496 58218 3505
rect 56600 2984 56652 2990
rect 56598 2952 56600 2961
rect 56652 2952 56654 2961
rect 56598 2887 56654 2896
rect 55310 2816 55366 2825
rect 55310 2751 55366 2760
rect 55956 2440 56008 2446
rect 55956 2382 56008 2388
rect 56600 2440 56652 2446
rect 56600 2382 56652 2388
rect 55968 2106 55996 2382
rect 55956 2100 56008 2106
rect 55956 2042 56008 2048
rect 56612 1426 56640 2382
rect 57532 2145 57560 3470
rect 58162 3431 58218 3440
rect 57888 2508 57940 2514
rect 57888 2450 57940 2456
rect 57518 2136 57574 2145
rect 57518 2071 57574 2080
rect 57900 2038 57928 2450
rect 57888 2032 57940 2038
rect 57888 1974 57940 1980
rect 56600 1420 56652 1426
rect 56600 1362 56652 1368
rect 54760 876 54812 882
rect 54760 818 54812 824
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5814 0 5870 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6090 0 6146 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6366 0 6422 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6734 0 6790 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7010 0 7066 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53194 0 53250 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 58452 785 58480 3878
rect 58438 776 58494 785
rect 58438 711 58494 720
<< via2 >>
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 58438 59200 58494 59256
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 18510 56788 18512 56808
rect 18512 56788 18564 56808
rect 18564 56788 18566 56808
rect 18510 56752 18566 56788
rect 16210 55564 16212 55584
rect 16212 55564 16264 55584
rect 16264 55564 16266 55584
rect 16210 55528 16266 55564
rect 17130 55292 17132 55312
rect 17132 55292 17184 55312
rect 17184 55292 17186 55312
rect 17130 55256 17186 55292
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 5262 31320 5318 31376
rect 4618 26288 4674 26344
rect 5078 26288 5134 26344
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 2042 3168 2098 3224
rect 1766 2896 1822 2952
rect 2962 7928 3018 7984
rect 3238 3576 3294 3632
rect 3146 3032 3202 3088
rect 3606 4120 3662 4176
rect 3790 3984 3846 4040
rect 3238 2624 3294 2680
rect 3974 7928 4030 7984
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4526 5108 4528 5128
rect 4528 5108 4580 5128
rect 4580 5108 4582 5128
rect 4526 5072 4582 5108
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4894 11600 4950 11656
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4986 4664 5042 4720
rect 4894 2760 4950 2816
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 5814 14220 5816 14240
rect 5816 14220 5868 14240
rect 5868 14220 5870 14240
rect 5814 14184 5870 14220
rect 7470 31340 7526 31376
rect 7470 31320 7472 31340
rect 7472 31320 7524 31340
rect 7524 31320 7526 31340
rect 7930 26324 7932 26344
rect 7932 26324 7984 26344
rect 7984 26324 7986 26344
rect 7930 26288 7986 26324
rect 8482 28464 8538 28520
rect 8114 18672 8170 18728
rect 9402 28500 9404 28520
rect 9404 28500 9456 28520
rect 9456 28500 9458 28520
rect 9402 28464 9458 28500
rect 7746 14728 7802 14784
rect 7654 13912 7710 13968
rect 7562 13776 7618 13832
rect 7654 12552 7710 12608
rect 5538 3440 5594 3496
rect 5906 4256 5962 4312
rect 5814 3984 5870 4040
rect 5906 3340 5908 3360
rect 5908 3340 5960 3360
rect 5960 3340 5962 3360
rect 5906 3304 5962 3340
rect 5814 2760 5870 2816
rect 6090 2896 6146 2952
rect 6090 1264 6146 1320
rect 6366 4156 6368 4176
rect 6368 4156 6420 4176
rect 6420 4156 6422 4176
rect 6366 4120 6422 4156
rect 6918 7520 6974 7576
rect 6734 3884 6736 3904
rect 6736 3884 6788 3904
rect 6788 3884 6790 3904
rect 6734 3848 6790 3884
rect 6274 1264 6330 1320
rect 6734 3168 6790 3224
rect 6734 2252 6736 2272
rect 6736 2252 6788 2272
rect 6788 2252 6790 2272
rect 6734 2216 6790 2252
rect 7286 4700 7288 4720
rect 7288 4700 7340 4720
rect 7340 4700 7342 4720
rect 7286 4664 7342 4700
rect 7194 4256 7250 4312
rect 7654 3712 7710 3768
rect 8022 5072 8078 5128
rect 7838 3032 7894 3088
rect 10230 31184 10286 31240
rect 9402 15544 9458 15600
rect 9678 14220 9680 14240
rect 9680 14220 9732 14240
rect 9732 14220 9734 14240
rect 9678 14184 9734 14220
rect 10690 23840 10746 23896
rect 10966 17992 11022 18048
rect 12438 29008 12494 29064
rect 18050 55564 18052 55584
rect 18052 55564 18104 55584
rect 18104 55564 18106 55584
rect 18050 55528 18106 55564
rect 15014 31220 15016 31240
rect 15016 31220 15068 31240
rect 15068 31220 15070 31240
rect 15014 31184 15070 31220
rect 11702 16632 11758 16688
rect 8482 5092 8538 5128
rect 8482 5072 8484 5092
rect 8484 5072 8536 5092
rect 8536 5072 8538 5092
rect 8298 3732 8354 3768
rect 8298 3712 8300 3732
rect 8300 3712 8352 3732
rect 8352 3712 8354 3732
rect 8482 3576 8538 3632
rect 8942 3984 8998 4040
rect 9770 7928 9826 7984
rect 10322 9868 10324 9888
rect 10324 9868 10376 9888
rect 10376 9868 10378 9888
rect 10322 9832 10378 9868
rect 10138 6840 10194 6896
rect 10046 3984 10102 4040
rect 10414 2644 10470 2680
rect 10414 2624 10416 2644
rect 10416 2624 10468 2644
rect 10468 2624 10470 2644
rect 10874 3168 10930 3224
rect 12530 8200 12586 8256
rect 12898 3848 12954 3904
rect 13450 2644 13506 2680
rect 13450 2624 13452 2644
rect 13452 2624 13504 2644
rect 13504 2624 13506 2644
rect 14646 23860 14702 23896
rect 14646 23840 14648 23860
rect 14648 23840 14700 23860
rect 14700 23840 14702 23860
rect 13726 8200 13782 8256
rect 13910 6704 13966 6760
rect 15382 27396 15438 27432
rect 15382 27376 15384 27396
rect 15384 27376 15436 27396
rect 15436 27376 15438 27396
rect 14554 7284 14556 7304
rect 14556 7284 14608 7304
rect 14608 7284 14610 7304
rect 14554 7248 14610 7284
rect 14830 6840 14886 6896
rect 14830 5616 14886 5672
rect 14094 3340 14096 3360
rect 14096 3340 14148 3360
rect 14148 3340 14150 3360
rect 14094 3304 14150 3340
rect 14554 3188 14610 3224
rect 14554 3168 14556 3188
rect 14556 3168 14608 3188
rect 14608 3168 14610 3188
rect 14554 2644 14610 2680
rect 14554 2624 14556 2644
rect 14556 2624 14608 2644
rect 14608 2624 14610 2644
rect 15842 21936 15898 21992
rect 15474 6704 15530 6760
rect 15474 5652 15476 5672
rect 15476 5652 15528 5672
rect 15528 5652 15530 5672
rect 15474 5616 15530 5652
rect 16118 3732 16174 3768
rect 16118 3712 16120 3732
rect 16120 3712 16172 3732
rect 16172 3712 16174 3732
rect 16118 3188 16174 3224
rect 16118 3168 16120 3188
rect 16120 3168 16172 3188
rect 16172 3168 16174 3188
rect 16946 21972 16948 21992
rect 16948 21972 17000 21992
rect 17000 21972 17002 21992
rect 16946 21936 17002 21972
rect 16762 16668 16764 16688
rect 16764 16668 16816 16688
rect 16816 16668 16818 16688
rect 16762 16632 16818 16668
rect 16854 6840 16910 6896
rect 16394 3984 16450 4040
rect 17130 3984 17186 4040
rect 20074 57196 20076 57216
rect 20076 57196 20128 57216
rect 20128 57196 20130 57216
rect 20074 57160 20130 57196
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 25134 56652 25136 56672
rect 25136 56652 25188 56672
rect 25188 56652 25190 56672
rect 25134 56616 25190 56652
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 18970 55292 18972 55312
rect 18972 55292 19024 55312
rect 19024 55292 19026 55312
rect 18970 55256 19026 55292
rect 18786 37304 18842 37360
rect 18602 17992 18658 18048
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19338 41420 19340 41440
rect 19340 41420 19392 41440
rect 19392 41420 19394 41440
rect 19338 41384 19394 41420
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19338 41112 19394 41168
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 18602 12280 18658 12336
rect 18142 7284 18144 7304
rect 18144 7284 18196 7304
rect 18196 7284 18198 7304
rect 18142 7248 18198 7284
rect 19246 20460 19302 20496
rect 19246 20440 19248 20460
rect 19248 20440 19300 20460
rect 19300 20440 19302 20460
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19246 12280 19302 12336
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 20350 55564 20352 55584
rect 20352 55564 20404 55584
rect 20404 55564 20406 55584
rect 20350 55528 20406 55564
rect 17590 5072 17646 5128
rect 17682 4120 17738 4176
rect 17774 3732 17830 3768
rect 17774 3712 17776 3732
rect 17776 3712 17828 3732
rect 17828 3712 17830 3732
rect 18142 3984 18198 4040
rect 18050 2624 18106 2680
rect 18602 3984 18658 4040
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 18786 3168 18842 3224
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19430 3188 19486 3224
rect 19430 3168 19432 3188
rect 19432 3168 19484 3188
rect 19484 3168 19486 3188
rect 19522 3032 19578 3088
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 20534 13640 20590 13696
rect 20810 17604 20866 17640
rect 20810 17584 20812 17604
rect 20812 17584 20864 17604
rect 20864 17584 20866 17604
rect 22558 55564 22560 55584
rect 22560 55564 22612 55584
rect 22612 55564 22614 55584
rect 22558 55528 22614 55564
rect 22742 35944 22798 36000
rect 22006 22228 22062 22264
rect 22006 22208 22008 22228
rect 22008 22208 22060 22228
rect 22060 22208 22062 22228
rect 20350 3712 20406 3768
rect 20258 3440 20314 3496
rect 20350 3304 20406 3360
rect 20166 2624 20222 2680
rect 20534 3168 20590 3224
rect 20994 3984 21050 4040
rect 21914 7148 21916 7168
rect 21916 7148 21968 7168
rect 21968 7148 21970 7168
rect 21914 7112 21970 7148
rect 22558 24792 22614 24848
rect 23570 27376 23626 27432
rect 24950 44920 25006 44976
rect 22834 20748 22836 20768
rect 22836 20748 22888 20768
rect 22888 20748 22890 20768
rect 22834 20712 22890 20748
rect 23478 20712 23534 20768
rect 22926 17620 22928 17640
rect 22928 17620 22980 17640
rect 22980 17620 22982 17640
rect 22926 17584 22982 17620
rect 23662 13912 23718 13968
rect 24950 17584 25006 17640
rect 24306 15544 24362 15600
rect 25226 20476 25228 20496
rect 25228 20476 25280 20496
rect 25280 20476 25282 20496
rect 25226 20440 25282 20476
rect 26330 42064 26386 42120
rect 24030 12552 24086 12608
rect 24582 13776 24638 13832
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 29642 53080 29698 53136
rect 27158 44784 27214 44840
rect 27618 29028 27674 29064
rect 27618 29008 27620 29028
rect 27620 29008 27672 29028
rect 27672 29008 27674 29028
rect 25962 7112 26018 7168
rect 26974 17584 27030 17640
rect 27526 15408 27582 15464
rect 27526 6840 27582 6896
rect 29366 6296 29422 6352
rect 30562 18672 30618 18728
rect 30930 18828 30986 18864
rect 30930 18808 30932 18828
rect 30932 18808 30984 18828
rect 30984 18808 30986 18828
rect 32126 50224 32182 50280
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 33230 36780 33286 36816
rect 33230 36760 33232 36780
rect 33232 36760 33284 36780
rect 33284 36760 33286 36780
rect 33782 36760 33838 36816
rect 33506 30252 33562 30288
rect 33506 30232 33508 30252
rect 33508 30232 33560 30252
rect 33560 30232 33562 30252
rect 29918 3576 29974 3632
rect 32126 22652 32128 22672
rect 32128 22652 32180 22672
rect 32180 22652 32182 22672
rect 32126 22616 32182 22652
rect 32218 20440 32274 20496
rect 32862 20460 32918 20496
rect 32862 20440 32864 20460
rect 32864 20440 32916 20460
rect 32916 20440 32918 20460
rect 32586 17604 32642 17640
rect 32586 17584 32588 17604
rect 32588 17584 32640 17604
rect 32640 17584 32642 17604
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35346 36780 35402 36816
rect 35346 36760 35348 36780
rect 35348 36760 35400 36780
rect 35400 36760 35402 36780
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34334 30252 34390 30288
rect 34334 30232 34336 30252
rect 34336 30232 34388 30252
rect 34388 30232 34390 30252
rect 34058 22652 34060 22672
rect 34060 22652 34112 22672
rect 34112 22652 34114 22672
rect 34058 22616 34114 22652
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34426 6332 34428 6352
rect 34428 6332 34480 6352
rect 34480 6332 34482 6352
rect 34426 6296 34482 6332
rect 57518 57840 57574 57896
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 57886 56480 57942 56536
rect 36082 18844 36084 18864
rect 36084 18844 36136 18864
rect 36136 18844 36138 18864
rect 36082 18808 36138 18844
rect 35622 17620 35624 17640
rect 35624 17620 35676 17640
rect 35676 17620 35678 17640
rect 35622 17584 35678 17620
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35806 15408 35862 15464
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 58162 55140 58218 55176
rect 58162 55120 58164 55140
rect 58164 55120 58216 55140
rect 58216 55120 58218 55140
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 57886 53760 57942 53816
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 57886 52436 57888 52456
rect 57888 52436 57940 52456
rect 57940 52436 57942 52456
rect 57886 52400 57942 52436
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 58162 51040 58218 51096
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 58162 49716 58164 49736
rect 58164 49716 58216 49736
rect 58216 49716 58218 49736
rect 58162 49680 58218 49716
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 58162 48320 58218 48376
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 58162 46996 58164 47016
rect 58164 46996 58216 47016
rect 58216 46996 58218 47016
rect 58162 46960 58218 46996
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 58162 45600 58218 45656
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 58162 44260 58218 44296
rect 58162 44240 58164 44260
rect 58164 44240 58216 44260
rect 58216 44240 58218 44260
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 58162 42880 58218 42936
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 58162 41556 58164 41576
rect 58164 41556 58216 41576
rect 58216 41556 58218 41576
rect 58162 41520 58218 41556
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 58162 40160 58218 40216
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 58162 38820 58218 38856
rect 58162 38800 58164 38820
rect 58164 38800 58216 38820
rect 58216 38800 58218 38820
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 58162 37440 58218 37496
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 58162 36116 58164 36136
rect 58164 36116 58216 36136
rect 58216 36116 58218 36136
rect 58162 36080 58218 36116
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 58162 34720 58218 34776
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 58162 33380 58218 33416
rect 58162 33360 58164 33380
rect 58164 33360 58216 33380
rect 58216 33360 58218 33380
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 58162 32000 58218 32056
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 58162 30676 58164 30696
rect 58164 30676 58216 30696
rect 58216 30676 58218 30696
rect 58162 30640 58218 30676
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 58162 29280 58218 29336
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 58162 27940 58218 27976
rect 58162 27920 58164 27940
rect 58164 27920 58216 27940
rect 58216 27920 58218 27940
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 58162 26560 58218 26616
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 58162 25236 58164 25256
rect 58164 25236 58216 25256
rect 58216 25236 58218 25256
rect 58162 25200 58218 25236
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 58162 23840 58218 23896
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 58162 22500 58218 22536
rect 58162 22480 58164 22500
rect 58164 22480 58216 22500
rect 58216 22480 58218 22500
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 58162 21120 58218 21176
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 58162 19796 58164 19816
rect 58164 19796 58216 19816
rect 58216 19796 58218 19816
rect 58162 19760 58218 19796
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 58162 18400 58218 18456
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 58162 17060 58218 17096
rect 58162 17040 58164 17060
rect 58164 17040 58216 17060
rect 58216 17040 58218 17060
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 58162 15680 58218 15736
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 58162 14356 58164 14376
rect 58164 14356 58216 14376
rect 58216 14356 58218 14376
rect 58162 14320 58218 14356
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 58162 12960 58218 13016
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 58162 11620 58218 11656
rect 58162 11600 58164 11620
rect 58164 11600 58216 11620
rect 58216 11600 58218 11620
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 58162 10240 58218 10296
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 58162 8916 58164 8936
rect 58164 8916 58216 8936
rect 58216 8916 58218 8936
rect 58162 8880 58218 8916
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 58162 7520 58218 7576
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 58162 6180 58218 6216
rect 58162 6160 58164 6180
rect 58164 6160 58216 6180
rect 58216 6160 58218 6180
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 53378 2896 53434 2952
rect 53470 2760 53526 2816
rect 58162 4800 58218 4856
rect 58162 3476 58164 3496
rect 58164 3476 58216 3496
rect 58216 3476 58218 3496
rect 56598 2932 56600 2952
rect 56600 2932 56652 2952
rect 56652 2932 56654 2952
rect 56598 2896 56654 2932
rect 55310 2760 55366 2816
rect 58162 3440 58218 3476
rect 57518 2080 57574 2136
rect 58438 720 58494 776
<< metal3 >>
rect 58433 59258 58499 59261
rect 59200 59258 60000 59288
rect 58433 59256 60000 59258
rect 58433 59200 58438 59256
rect 58494 59200 60000 59256
rect 58433 59198 60000 59200
rect 58433 59195 58499 59198
rect 59200 59168 60000 59198
rect 57513 57898 57579 57901
rect 59200 57898 60000 57928
rect 57513 57896 60000 57898
rect 57513 57840 57518 57896
rect 57574 57840 60000 57896
rect 57513 57838 60000 57840
rect 57513 57835 57579 57838
rect 59200 57808 60000 57838
rect 19570 57696 19886 57697
rect 0 57536 800 57656
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 20069 57218 20135 57221
rect 20478 57218 20484 57220
rect 20069 57216 20484 57218
rect 20069 57160 20074 57216
rect 20130 57160 20484 57216
rect 20069 57158 20484 57160
rect 20069 57155 20135 57158
rect 20478 57156 20484 57158
rect 20548 57156 20554 57220
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 18505 56810 18571 56813
rect 18638 56810 18644 56812
rect 18505 56808 18644 56810
rect 18505 56752 18510 56808
rect 18566 56752 18644 56808
rect 18505 56750 18644 56752
rect 18505 56747 18571 56750
rect 18638 56748 18644 56750
rect 18708 56748 18714 56812
rect 21398 56612 21404 56676
rect 21468 56674 21474 56676
rect 25129 56674 25195 56677
rect 21468 56672 25195 56674
rect 21468 56616 25134 56672
rect 25190 56616 25195 56672
rect 21468 56614 25195 56616
rect 21468 56612 21474 56614
rect 25129 56611 25195 56614
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 57881 56538 57947 56541
rect 59200 56538 60000 56568
rect 57881 56536 60000 56538
rect 57881 56480 57886 56536
rect 57942 56480 60000 56536
rect 57881 56478 60000 56480
rect 57881 56475 57947 56478
rect 59200 56448 60000 56478
rect 0 56040 800 56160
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 16205 55588 16271 55589
rect 16205 55586 16252 55588
rect 16160 55584 16252 55586
rect 16160 55528 16210 55584
rect 16160 55526 16252 55528
rect 16205 55524 16252 55526
rect 16316 55524 16322 55588
rect 18045 55586 18111 55589
rect 20345 55588 20411 55589
rect 18270 55586 18276 55588
rect 18045 55584 18276 55586
rect 18045 55528 18050 55584
rect 18106 55528 18276 55584
rect 18045 55526 18276 55528
rect 16205 55523 16271 55524
rect 18045 55523 18111 55526
rect 18270 55524 18276 55526
rect 18340 55524 18346 55588
rect 20294 55524 20300 55588
rect 20364 55586 20411 55588
rect 22553 55586 22619 55589
rect 22686 55586 22692 55588
rect 20364 55584 20456 55586
rect 20406 55528 20456 55584
rect 20364 55526 20456 55528
rect 22553 55584 22692 55586
rect 22553 55528 22558 55584
rect 22614 55528 22692 55584
rect 22553 55526 22692 55528
rect 20364 55524 20411 55526
rect 20345 55523 20411 55524
rect 22553 55523 22619 55526
rect 22686 55524 22692 55526
rect 22756 55524 22762 55588
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 17125 55316 17191 55317
rect 17125 55314 17172 55316
rect 17080 55312 17172 55314
rect 17080 55256 17130 55312
rect 17080 55254 17172 55256
rect 17125 55252 17172 55254
rect 17236 55252 17242 55316
rect 18454 55252 18460 55316
rect 18524 55314 18530 55316
rect 18965 55314 19031 55317
rect 18524 55312 19031 55314
rect 18524 55256 18970 55312
rect 19026 55256 19031 55312
rect 18524 55254 19031 55256
rect 18524 55252 18530 55254
rect 17125 55251 17191 55252
rect 18965 55251 19031 55254
rect 58157 55178 58223 55181
rect 59200 55178 60000 55208
rect 58157 55176 60000 55178
rect 58157 55120 58162 55176
rect 58218 55120 60000 55176
rect 58157 55118 60000 55120
rect 58157 55115 58223 55118
rect 59200 55088 60000 55118
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 0 54544 800 54664
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 57881 53818 57947 53821
rect 59200 53818 60000 53848
rect 57881 53816 60000 53818
rect 57881 53760 57886 53816
rect 57942 53760 60000 53816
rect 57881 53758 60000 53760
rect 57881 53755 57947 53758
rect 59200 53728 60000 53758
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 0 53048 800 53168
rect 13486 53076 13492 53140
rect 13556 53138 13562 53140
rect 29637 53138 29703 53141
rect 13556 53136 29703 53138
rect 13556 53080 29642 53136
rect 29698 53080 29703 53136
rect 13556 53078 29703 53080
rect 13556 53076 13562 53078
rect 29637 53075 29703 53078
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 57881 52458 57947 52461
rect 59200 52458 60000 52488
rect 57881 52456 60000 52458
rect 57881 52400 57886 52456
rect 57942 52400 60000 52456
rect 57881 52398 60000 52400
rect 57881 52395 57947 52398
rect 59200 52368 60000 52398
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 0 51552 800 51672
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 58157 51098 58223 51101
rect 59200 51098 60000 51128
rect 58157 51096 60000 51098
rect 58157 51040 58162 51096
rect 58218 51040 60000 51096
rect 58157 51038 60000 51040
rect 58157 51035 58223 51038
rect 59200 51008 60000 51038
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 16430 50220 16436 50284
rect 16500 50282 16506 50284
rect 32121 50282 32187 50285
rect 16500 50280 32187 50282
rect 16500 50224 32126 50280
rect 32182 50224 32187 50280
rect 16500 50222 32187 50224
rect 16500 50220 16506 50222
rect 32121 50219 32187 50222
rect 0 50056 800 50176
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 58157 49738 58223 49741
rect 59200 49738 60000 49768
rect 58157 49736 60000 49738
rect 58157 49680 58162 49736
rect 58218 49680 60000 49736
rect 58157 49678 60000 49680
rect 58157 49675 58223 49678
rect 59200 49648 60000 49678
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 0 48560 800 48680
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 58157 48378 58223 48381
rect 59200 48378 60000 48408
rect 58157 48376 60000 48378
rect 58157 48320 58162 48376
rect 58218 48320 60000 48376
rect 58157 48318 60000 48320
rect 58157 48315 58223 48318
rect 59200 48288 60000 48318
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 0 47064 800 47184
rect 58157 47018 58223 47021
rect 59200 47018 60000 47048
rect 58157 47016 60000 47018
rect 58157 46960 58162 47016
rect 58218 46960 60000 47016
rect 58157 46958 60000 46960
rect 58157 46955 58223 46958
rect 59200 46928 60000 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 0 45568 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 58157 45658 58223 45661
rect 59200 45658 60000 45688
rect 58157 45656 60000 45658
rect 58157 45600 58162 45656
rect 58218 45600 60000 45656
rect 58157 45598 60000 45600
rect 58157 45595 58223 45598
rect 59200 45568 60000 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 14774 44916 14780 44980
rect 14844 44978 14850 44980
rect 24945 44978 25011 44981
rect 14844 44976 25011 44978
rect 14844 44920 24950 44976
rect 25006 44920 25011 44976
rect 14844 44918 25011 44920
rect 14844 44916 14850 44918
rect 24945 44915 25011 44918
rect 14590 44780 14596 44844
rect 14660 44842 14666 44844
rect 27153 44842 27219 44845
rect 14660 44840 27219 44842
rect 14660 44784 27158 44840
rect 27214 44784 27219 44840
rect 14660 44782 27219 44784
rect 14660 44780 14666 44782
rect 27153 44779 27219 44782
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 58157 44298 58223 44301
rect 59200 44298 60000 44328
rect 58157 44296 60000 44298
rect 58157 44240 58162 44296
rect 58218 44240 60000 44296
rect 58157 44238 60000 44240
rect 58157 44235 58223 44238
rect 59200 44208 60000 44238
rect 0 44072 800 44192
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 58157 42938 58223 42941
rect 59200 42938 60000 42968
rect 58157 42936 60000 42938
rect 58157 42880 58162 42936
rect 58218 42880 60000 42936
rect 58157 42878 60000 42880
rect 58157 42875 58223 42878
rect 59200 42848 60000 42878
rect 0 42576 800 42696
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 17350 42060 17356 42124
rect 17420 42122 17426 42124
rect 26325 42122 26391 42125
rect 17420 42120 26391 42122
rect 17420 42064 26330 42120
rect 26386 42064 26391 42120
rect 17420 42062 26391 42064
rect 17420 42060 17426 42062
rect 26325 42059 26391 42062
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 58157 41578 58223 41581
rect 59200 41578 60000 41608
rect 58157 41576 60000 41578
rect 58157 41520 58162 41576
rect 58218 41520 60000 41576
rect 58157 41518 60000 41520
rect 58157 41515 58223 41518
rect 59200 41488 60000 41518
rect 19333 41442 19399 41445
rect 19333 41440 19442 41442
rect 19333 41384 19338 41440
rect 19394 41384 19442 41440
rect 19333 41379 19442 41384
rect 0 41080 800 41200
rect 19382 41173 19442 41379
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 19333 41168 19442 41173
rect 19333 41112 19338 41168
rect 19394 41112 19442 41168
rect 19333 41110 19442 41112
rect 19333 41107 19399 41110
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 58157 40218 58223 40221
rect 59200 40218 60000 40248
rect 58157 40216 60000 40218
rect 58157 40160 58162 40216
rect 58218 40160 60000 40216
rect 58157 40158 60000 40160
rect 58157 40155 58223 40158
rect 59200 40128 60000 40158
rect 4210 39744 4526 39745
rect 0 39584 800 39704
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 58157 38858 58223 38861
rect 59200 38858 60000 38888
rect 58157 38856 60000 38858
rect 58157 38800 58162 38856
rect 58218 38800 60000 38856
rect 58157 38798 60000 38800
rect 58157 38795 58223 38798
rect 59200 38768 60000 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 0 38088 800 38208
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 58157 37498 58223 37501
rect 59200 37498 60000 37528
rect 58157 37496 60000 37498
rect 58157 37440 58162 37496
rect 58218 37440 60000 37496
rect 58157 37438 60000 37440
rect 58157 37435 58223 37438
rect 59200 37408 60000 37438
rect 18781 37362 18847 37365
rect 19374 37362 19380 37364
rect 18781 37360 19380 37362
rect 18781 37304 18786 37360
rect 18842 37304 19380 37360
rect 18781 37302 19380 37304
rect 18781 37299 18847 37302
rect 19374 37300 19380 37302
rect 19444 37300 19450 37364
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 33225 36818 33291 36821
rect 33777 36818 33843 36821
rect 35341 36818 35407 36821
rect 33225 36816 35407 36818
rect 33225 36760 33230 36816
rect 33286 36760 33782 36816
rect 33838 36760 35346 36816
rect 35402 36760 35407 36816
rect 33225 36758 35407 36760
rect 33225 36755 33291 36758
rect 33777 36755 33843 36758
rect 35341 36755 35407 36758
rect 0 36592 800 36712
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 58157 36138 58223 36141
rect 59200 36138 60000 36168
rect 58157 36136 60000 36138
rect 58157 36080 58162 36136
rect 58218 36080 60000 36136
rect 58157 36078 60000 36080
rect 58157 36075 58223 36078
rect 59200 36048 60000 36078
rect 22502 35940 22508 36004
rect 22572 36002 22578 36004
rect 22737 36002 22803 36005
rect 22572 36000 22803 36002
rect 22572 35944 22742 36000
rect 22798 35944 22803 36000
rect 22572 35942 22803 35944
rect 22572 35940 22578 35942
rect 22737 35939 22803 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 0 35096 800 35216
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 58157 34778 58223 34781
rect 59200 34778 60000 34808
rect 58157 34776 60000 34778
rect 58157 34720 58162 34776
rect 58218 34720 60000 34776
rect 58157 34718 60000 34720
rect 58157 34715 58223 34718
rect 59200 34688 60000 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 0 33600 800 33720
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 58157 33418 58223 33421
rect 59200 33418 60000 33448
rect 58157 33416 60000 33418
rect 58157 33360 58162 33416
rect 58218 33360 60000 33416
rect 58157 33358 60000 33360
rect 58157 33355 58223 33358
rect 59200 33328 60000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 0 32104 800 32224
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 58157 32058 58223 32061
rect 59200 32058 60000 32088
rect 58157 32056 60000 32058
rect 58157 32000 58162 32056
rect 58218 32000 60000 32056
rect 58157 31998 60000 32000
rect 58157 31995 58223 31998
rect 59200 31968 60000 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 5257 31378 5323 31381
rect 7465 31378 7531 31381
rect 5257 31376 7531 31378
rect 5257 31320 5262 31376
rect 5318 31320 7470 31376
rect 7526 31320 7531 31376
rect 5257 31318 7531 31320
rect 5257 31315 5323 31318
rect 7465 31315 7531 31318
rect 10225 31242 10291 31245
rect 15009 31242 15075 31245
rect 10225 31240 15075 31242
rect 10225 31184 10230 31240
rect 10286 31184 15014 31240
rect 15070 31184 15075 31240
rect 10225 31182 15075 31184
rect 10225 31179 10291 31182
rect 15009 31179 15075 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 0 30608 800 30728
rect 58157 30698 58223 30701
rect 59200 30698 60000 30728
rect 58157 30696 60000 30698
rect 58157 30640 58162 30696
rect 58218 30640 60000 30696
rect 58157 30638 60000 30640
rect 58157 30635 58223 30638
rect 59200 30608 60000 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 33501 30290 33567 30293
rect 34329 30290 34395 30293
rect 33501 30288 34395 30290
rect 33501 30232 33506 30288
rect 33562 30232 34334 30288
rect 34390 30232 34395 30288
rect 33501 30230 34395 30232
rect 33501 30227 33567 30230
rect 34329 30227 34395 30230
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 58157 29338 58223 29341
rect 59200 29338 60000 29368
rect 58157 29336 60000 29338
rect 58157 29280 58162 29336
rect 58218 29280 60000 29336
rect 58157 29278 60000 29280
rect 58157 29275 58223 29278
rect 59200 29248 60000 29278
rect 0 29112 800 29232
rect 12433 29066 12499 29069
rect 21950 29066 21956 29068
rect 12433 29064 21956 29066
rect 12433 29008 12438 29064
rect 12494 29008 21956 29064
rect 12433 29006 21956 29008
rect 12433 29003 12499 29006
rect 21950 29004 21956 29006
rect 22020 29066 22026 29068
rect 27613 29066 27679 29069
rect 22020 29064 27679 29066
rect 22020 29008 27618 29064
rect 27674 29008 27679 29064
rect 22020 29006 27679 29008
rect 22020 29004 22026 29006
rect 27613 29003 27679 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 8477 28522 8543 28525
rect 9397 28522 9463 28525
rect 8477 28520 9463 28522
rect 8477 28464 8482 28520
rect 8538 28464 9402 28520
rect 9458 28464 9463 28520
rect 8477 28462 9463 28464
rect 8477 28459 8543 28462
rect 9397 28459 9463 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 58157 27978 58223 27981
rect 59200 27978 60000 28008
rect 58157 27976 60000 27978
rect 58157 27920 58162 27976
rect 58218 27920 60000 27976
rect 58157 27918 60000 27920
rect 58157 27915 58223 27918
rect 59200 27888 60000 27918
rect 4210 27776 4526 27777
rect 0 27616 800 27736
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 15377 27434 15443 27437
rect 23565 27434 23631 27437
rect 15377 27432 23631 27434
rect 15377 27376 15382 27432
rect 15438 27376 23570 27432
rect 23626 27376 23631 27432
rect 15377 27374 23631 27376
rect 15377 27371 15443 27374
rect 23565 27371 23631 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 58157 26618 58223 26621
rect 59200 26618 60000 26648
rect 58157 26616 60000 26618
rect 58157 26560 58162 26616
rect 58218 26560 60000 26616
rect 58157 26558 60000 26560
rect 58157 26555 58223 26558
rect 59200 26528 60000 26558
rect 4613 26346 4679 26349
rect 5073 26346 5139 26349
rect 7925 26346 7991 26349
rect 4613 26344 7991 26346
rect 4613 26288 4618 26344
rect 4674 26288 5078 26344
rect 5134 26288 7930 26344
rect 7986 26288 7991 26344
rect 4613 26286 7991 26288
rect 4613 26283 4679 26286
rect 5073 26283 5139 26286
rect 7925 26283 7991 26286
rect 0 26120 800 26240
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 58157 25258 58223 25261
rect 59200 25258 60000 25288
rect 58157 25256 60000 25258
rect 58157 25200 58162 25256
rect 58218 25200 60000 25256
rect 58157 25198 60000 25200
rect 58157 25195 58223 25198
rect 59200 25168 60000 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 22553 24852 22619 24853
rect 22502 24850 22508 24852
rect 22462 24790 22508 24850
rect 22572 24848 22619 24852
rect 22614 24792 22619 24848
rect 22502 24788 22508 24790
rect 22572 24788 22619 24792
rect 22553 24787 22619 24788
rect 0 24624 800 24744
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 10685 23898 10751 23901
rect 14641 23898 14707 23901
rect 10685 23896 14707 23898
rect 10685 23840 10690 23896
rect 10746 23840 14646 23896
rect 14702 23840 14707 23896
rect 10685 23838 14707 23840
rect 10685 23835 10751 23838
rect 14641 23835 14707 23838
rect 58157 23898 58223 23901
rect 59200 23898 60000 23928
rect 58157 23896 60000 23898
rect 58157 23840 58162 23896
rect 58218 23840 60000 23896
rect 58157 23838 60000 23840
rect 58157 23835 58223 23838
rect 59200 23808 60000 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23128 800 23248
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 32121 22674 32187 22677
rect 34053 22674 34119 22677
rect 32121 22672 34119 22674
rect 32121 22616 32126 22672
rect 32182 22616 34058 22672
rect 34114 22616 34119 22672
rect 32121 22614 34119 22616
rect 32121 22611 32187 22614
rect 34053 22611 34119 22614
rect 58157 22538 58223 22541
rect 59200 22538 60000 22568
rect 58157 22536 60000 22538
rect 58157 22480 58162 22536
rect 58218 22480 60000 22536
rect 58157 22478 60000 22480
rect 58157 22475 58223 22478
rect 59200 22448 60000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 22001 22268 22067 22269
rect 21950 22266 21956 22268
rect 21910 22206 21956 22266
rect 22020 22264 22067 22268
rect 22062 22208 22067 22264
rect 21950 22204 21956 22206
rect 22020 22204 22067 22208
rect 22001 22203 22067 22204
rect 15837 21994 15903 21997
rect 16941 21994 17007 21997
rect 15837 21992 17007 21994
rect 15837 21936 15842 21992
rect 15898 21936 16946 21992
rect 17002 21936 17007 21992
rect 15837 21934 17007 21936
rect 15837 21931 15903 21934
rect 16941 21931 17007 21934
rect 19570 21792 19886 21793
rect 0 21632 800 21752
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 58157 21178 58223 21181
rect 59200 21178 60000 21208
rect 58157 21176 60000 21178
rect 58157 21120 58162 21176
rect 58218 21120 60000 21176
rect 58157 21118 60000 21120
rect 58157 21115 58223 21118
rect 59200 21088 60000 21118
rect 22829 20770 22895 20773
rect 23473 20770 23539 20773
rect 22829 20768 23539 20770
rect 22829 20712 22834 20768
rect 22890 20712 23478 20768
rect 23534 20712 23539 20768
rect 22829 20710 23539 20712
rect 22829 20707 22895 20710
rect 23473 20707 23539 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 19241 20498 19307 20501
rect 25221 20498 25287 20501
rect 19241 20496 25287 20498
rect 19241 20440 19246 20496
rect 19302 20440 25226 20496
rect 25282 20440 25287 20496
rect 19241 20438 25287 20440
rect 19241 20435 19307 20438
rect 25221 20435 25287 20438
rect 32213 20498 32279 20501
rect 32857 20498 32923 20501
rect 32213 20496 32923 20498
rect 32213 20440 32218 20496
rect 32274 20440 32862 20496
rect 32918 20440 32923 20496
rect 32213 20438 32923 20440
rect 32213 20435 32279 20438
rect 32857 20435 32923 20438
rect 0 20136 800 20256
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 58157 19818 58223 19821
rect 59200 19818 60000 19848
rect 58157 19816 60000 19818
rect 58157 19760 58162 19816
rect 58218 19760 60000 19816
rect 58157 19758 60000 19760
rect 58157 19755 58223 19758
rect 59200 19728 60000 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 30925 18866 30991 18869
rect 36077 18866 36143 18869
rect 30925 18864 36143 18866
rect 30925 18808 30930 18864
rect 30986 18808 36082 18864
rect 36138 18808 36143 18864
rect 30925 18806 36143 18808
rect 30925 18803 30991 18806
rect 36077 18803 36143 18806
rect 0 18640 800 18760
rect 8109 18730 8175 18733
rect 30557 18730 30623 18733
rect 8109 18728 30623 18730
rect 8109 18672 8114 18728
rect 8170 18672 30562 18728
rect 30618 18672 30623 18728
rect 8109 18670 30623 18672
rect 8109 18667 8175 18670
rect 30557 18667 30623 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 58157 18458 58223 18461
rect 59200 18458 60000 18488
rect 58157 18456 60000 18458
rect 58157 18400 58162 18456
rect 58218 18400 60000 18456
rect 58157 18398 60000 18400
rect 58157 18395 58223 18398
rect 59200 18368 60000 18398
rect 10961 18050 11027 18053
rect 18597 18050 18663 18053
rect 10961 18048 18663 18050
rect 10961 17992 10966 18048
rect 11022 17992 18602 18048
rect 18658 17992 18663 18048
rect 10961 17990 18663 17992
rect 10961 17987 11027 17990
rect 18597 17987 18663 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 20805 17642 20871 17645
rect 22921 17642 22987 17645
rect 20805 17640 22987 17642
rect 20805 17584 20810 17640
rect 20866 17584 22926 17640
rect 22982 17584 22987 17640
rect 20805 17582 22987 17584
rect 20805 17579 20871 17582
rect 22921 17579 22987 17582
rect 24945 17642 25011 17645
rect 26969 17642 27035 17645
rect 24945 17640 27035 17642
rect 24945 17584 24950 17640
rect 25006 17584 26974 17640
rect 27030 17584 27035 17640
rect 24945 17582 27035 17584
rect 24945 17579 25011 17582
rect 26969 17579 27035 17582
rect 32581 17642 32647 17645
rect 35617 17642 35683 17645
rect 32581 17640 35683 17642
rect 32581 17584 32586 17640
rect 32642 17584 35622 17640
rect 35678 17584 35683 17640
rect 32581 17582 35683 17584
rect 32581 17579 32647 17582
rect 35617 17579 35683 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 0 17144 800 17264
rect 58157 17098 58223 17101
rect 59200 17098 60000 17128
rect 58157 17096 60000 17098
rect 58157 17040 58162 17096
rect 58218 17040 60000 17096
rect 58157 17038 60000 17040
rect 58157 17035 58223 17038
rect 59200 17008 60000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 11697 16690 11763 16693
rect 16757 16690 16823 16693
rect 11697 16688 16823 16690
rect 11697 16632 11702 16688
rect 11758 16632 16762 16688
rect 16818 16632 16823 16688
rect 11697 16630 16823 16632
rect 11697 16627 11763 16630
rect 16757 16627 16823 16630
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 0 15648 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 58157 15738 58223 15741
rect 59200 15738 60000 15768
rect 58157 15736 60000 15738
rect 58157 15680 58162 15736
rect 58218 15680 60000 15736
rect 58157 15678 60000 15680
rect 58157 15675 58223 15678
rect 59200 15648 60000 15678
rect 9397 15602 9463 15605
rect 24301 15602 24367 15605
rect 9397 15600 24367 15602
rect 9397 15544 9402 15600
rect 9458 15544 24306 15600
rect 24362 15544 24367 15600
rect 9397 15542 24367 15544
rect 9397 15539 9463 15542
rect 24301 15539 24367 15542
rect 27521 15466 27587 15469
rect 35801 15466 35867 15469
rect 27521 15464 35867 15466
rect 27521 15408 27526 15464
rect 27582 15408 35806 15464
rect 35862 15408 35867 15464
rect 27521 15406 35867 15408
rect 27521 15403 27587 15406
rect 35801 15403 35867 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 5942 14724 5948 14788
rect 6012 14786 6018 14788
rect 7741 14786 7807 14789
rect 6012 14784 7807 14786
rect 6012 14728 7746 14784
rect 7802 14728 7807 14784
rect 6012 14726 7807 14728
rect 6012 14724 6018 14726
rect 7741 14723 7807 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 58157 14378 58223 14381
rect 59200 14378 60000 14408
rect 58157 14376 60000 14378
rect 58157 14320 58162 14376
rect 58218 14320 60000 14376
rect 58157 14318 60000 14320
rect 58157 14315 58223 14318
rect 59200 14288 60000 14318
rect 0 14152 800 14272
rect 5809 14242 5875 14245
rect 6494 14242 6500 14244
rect 5809 14240 6500 14242
rect 5809 14184 5814 14240
rect 5870 14184 6500 14240
rect 5809 14182 6500 14184
rect 5809 14179 5875 14182
rect 6494 14180 6500 14182
rect 6564 14180 6570 14244
rect 8886 14180 8892 14244
rect 8956 14242 8962 14244
rect 9673 14242 9739 14245
rect 8956 14240 9739 14242
rect 8956 14184 9678 14240
rect 9734 14184 9739 14240
rect 8956 14182 9739 14184
rect 8956 14180 8962 14182
rect 9673 14179 9739 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 7649 13970 7715 13973
rect 23657 13970 23723 13973
rect 7649 13968 23723 13970
rect 7649 13912 7654 13968
rect 7710 13912 23662 13968
rect 23718 13912 23723 13968
rect 7649 13910 23723 13912
rect 7649 13907 7715 13910
rect 23657 13907 23723 13910
rect 7557 13834 7623 13837
rect 24577 13834 24643 13837
rect 7557 13832 24643 13834
rect 7557 13776 7562 13832
rect 7618 13776 24582 13832
rect 24638 13776 24643 13832
rect 7557 13774 24643 13776
rect 7557 13771 7623 13774
rect 24577 13771 24643 13774
rect 20529 13698 20595 13701
rect 21214 13698 21220 13700
rect 20529 13696 21220 13698
rect 20529 13640 20534 13696
rect 20590 13640 21220 13696
rect 20529 13638 21220 13640
rect 20529 13635 20595 13638
rect 21214 13636 21220 13638
rect 21284 13636 21290 13700
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 58157 13018 58223 13021
rect 59200 13018 60000 13048
rect 58157 13016 60000 13018
rect 58157 12960 58162 13016
rect 58218 12960 60000 13016
rect 58157 12958 60000 12960
rect 58157 12955 58223 12958
rect 59200 12928 60000 12958
rect 0 12656 800 12776
rect 7649 12610 7715 12613
rect 8334 12610 8340 12612
rect 7649 12608 8340 12610
rect 7649 12552 7654 12608
rect 7710 12552 8340 12608
rect 7649 12550 8340 12552
rect 7649 12547 7715 12550
rect 8334 12548 8340 12550
rect 8404 12548 8410 12612
rect 17718 12548 17724 12612
rect 17788 12610 17794 12612
rect 24025 12610 24091 12613
rect 17788 12608 24091 12610
rect 17788 12552 24030 12608
rect 24086 12552 24091 12608
rect 17788 12550 24091 12552
rect 17788 12548 17794 12550
rect 24025 12547 24091 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 18597 12338 18663 12341
rect 19241 12338 19307 12341
rect 18597 12336 19307 12338
rect 18597 12280 18602 12336
rect 18658 12280 19246 12336
rect 19302 12280 19307 12336
rect 18597 12278 19307 12280
rect 18597 12275 18663 12278
rect 19241 12275 19307 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 3366 11596 3372 11660
rect 3436 11658 3442 11660
rect 4889 11658 4955 11661
rect 3436 11656 4955 11658
rect 3436 11600 4894 11656
rect 4950 11600 4955 11656
rect 3436 11598 4955 11600
rect 3436 11596 3442 11598
rect 4889 11595 4955 11598
rect 58157 11658 58223 11661
rect 59200 11658 60000 11688
rect 58157 11656 60000 11658
rect 58157 11600 58162 11656
rect 58218 11600 60000 11656
rect 58157 11598 60000 11600
rect 58157 11595 58223 11598
rect 59200 11568 60000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 0 11160 800 11280
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 58157 10298 58223 10301
rect 59200 10298 60000 10328
rect 58157 10296 60000 10298
rect 58157 10240 58162 10296
rect 58218 10240 60000 10296
rect 58157 10238 60000 10240
rect 58157 10235 58223 10238
rect 59200 10208 60000 10238
rect 16062 9964 16068 10028
rect 16132 10026 16138 10028
rect 21398 10026 21404 10028
rect 16132 9966 21404 10026
rect 16132 9964 16138 9966
rect 21398 9964 21404 9966
rect 21468 9964 21474 10028
rect 10317 9892 10383 9893
rect 10317 9890 10364 9892
rect 10272 9888 10364 9890
rect 10272 9832 10322 9888
rect 10272 9830 10364 9832
rect 10317 9828 10364 9830
rect 10428 9828 10434 9892
rect 10317 9827 10383 9828
rect 19570 9824 19886 9825
rect 0 9664 800 9784
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 58157 8938 58223 8941
rect 59200 8938 60000 8968
rect 58157 8936 60000 8938
rect 58157 8880 58162 8936
rect 58218 8880 60000 8936
rect 58157 8878 60000 8880
rect 58157 8875 58223 8878
rect 59200 8848 60000 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 0 8168 800 8288
rect 10910 8196 10916 8260
rect 10980 8258 10986 8260
rect 12525 8258 12591 8261
rect 13721 8258 13787 8261
rect 10980 8256 13787 8258
rect 10980 8200 12530 8256
rect 12586 8200 13726 8256
rect 13782 8200 13787 8256
rect 10980 8198 13787 8200
rect 10980 8196 10986 8198
rect 12525 8195 12591 8198
rect 13721 8195 13787 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 2957 7986 3023 7989
rect 3969 7986 4035 7989
rect 9765 7986 9831 7989
rect 2957 7984 9831 7986
rect 2957 7928 2962 7984
rect 3018 7928 3974 7984
rect 4030 7928 9770 7984
rect 9826 7928 9831 7984
rect 2957 7926 9831 7928
rect 2957 7923 3023 7926
rect 3969 7923 4035 7926
rect 9765 7923 9831 7926
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 6913 7578 6979 7581
rect 9622 7578 9628 7580
rect 6913 7576 9628 7578
rect 6913 7520 6918 7576
rect 6974 7520 9628 7576
rect 6913 7518 9628 7520
rect 6913 7515 6979 7518
rect 9622 7516 9628 7518
rect 9692 7516 9698 7580
rect 58157 7578 58223 7581
rect 59200 7578 60000 7608
rect 58157 7576 60000 7578
rect 58157 7520 58162 7576
rect 58218 7520 60000 7576
rect 58157 7518 60000 7520
rect 58157 7515 58223 7518
rect 59200 7488 60000 7518
rect 14549 7306 14615 7309
rect 18137 7306 18203 7309
rect 14549 7304 18203 7306
rect 14549 7248 14554 7304
rect 14610 7248 18142 7304
rect 18198 7248 18203 7304
rect 14549 7246 18203 7248
rect 14549 7243 14615 7246
rect 18137 7243 18203 7246
rect 21909 7170 21975 7173
rect 25957 7170 26023 7173
rect 21909 7168 26023 7170
rect 21909 7112 21914 7168
rect 21970 7112 25962 7168
rect 26018 7112 26023 7168
rect 21909 7110 26023 7112
rect 21909 7107 21975 7110
rect 25957 7107 26023 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 10133 6898 10199 6901
rect 14825 6898 14891 6901
rect 10133 6896 14891 6898
rect 10133 6840 10138 6896
rect 10194 6840 14830 6896
rect 14886 6840 14891 6896
rect 10133 6838 14891 6840
rect 10133 6835 10199 6838
rect 14825 6835 14891 6838
rect 16849 6898 16915 6901
rect 27521 6898 27587 6901
rect 16849 6896 27587 6898
rect 16849 6840 16854 6896
rect 16910 6840 27526 6896
rect 27582 6840 27587 6896
rect 16849 6838 27587 6840
rect 16849 6835 16915 6838
rect 27521 6835 27587 6838
rect 0 6672 800 6792
rect 13905 6762 13971 6765
rect 15469 6762 15535 6765
rect 13905 6760 15535 6762
rect 13905 6704 13910 6760
rect 13966 6704 15474 6760
rect 15530 6704 15535 6760
rect 13905 6702 15535 6704
rect 13905 6699 13971 6702
rect 15469 6699 15535 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 29361 6354 29427 6357
rect 34421 6354 34487 6357
rect 29361 6352 34487 6354
rect 29361 6296 29366 6352
rect 29422 6296 34426 6352
rect 34482 6296 34487 6352
rect 29361 6294 34487 6296
rect 29361 6291 29427 6294
rect 34421 6291 34487 6294
rect 58157 6218 58223 6221
rect 59200 6218 60000 6248
rect 58157 6216 60000 6218
rect 58157 6160 58162 6216
rect 58218 6160 60000 6216
rect 58157 6158 60000 6160
rect 58157 6155 58223 6158
rect 59200 6128 60000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 14825 5674 14891 5677
rect 15469 5674 15535 5677
rect 14825 5672 15535 5674
rect 14825 5616 14830 5672
rect 14886 5616 15474 5672
rect 15530 5616 15535 5672
rect 14825 5614 15535 5616
rect 14825 5611 14891 5614
rect 15469 5611 15535 5614
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 0 5176 800 5296
rect 4521 5130 4587 5133
rect 8017 5130 8083 5133
rect 4521 5128 8083 5130
rect 4521 5072 4526 5128
rect 4582 5072 8022 5128
rect 8078 5072 8083 5128
rect 4521 5070 8083 5072
rect 4521 5067 4587 5070
rect 8017 5067 8083 5070
rect 8477 5130 8543 5133
rect 17585 5130 17651 5133
rect 8477 5128 17651 5130
rect 8477 5072 8482 5128
rect 8538 5072 17590 5128
rect 17646 5072 17651 5128
rect 8477 5070 17651 5072
rect 8477 5067 8543 5070
rect 17585 5067 17651 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 58157 4858 58223 4861
rect 59200 4858 60000 4888
rect 58157 4856 60000 4858
rect 58157 4800 58162 4856
rect 58218 4800 60000 4856
rect 58157 4798 60000 4800
rect 58157 4795 58223 4798
rect 59200 4768 60000 4798
rect 4981 4722 5047 4725
rect 7281 4722 7347 4725
rect 4981 4720 7347 4722
rect 4981 4664 4986 4720
rect 5042 4664 7286 4720
rect 7342 4664 7347 4720
rect 4981 4662 7347 4664
rect 4981 4659 5047 4662
rect 7281 4659 7347 4662
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 5901 4314 5967 4317
rect 7189 4314 7255 4317
rect 5901 4312 7255 4314
rect 5901 4256 5906 4312
rect 5962 4256 7194 4312
rect 7250 4256 7255 4312
rect 5901 4254 7255 4256
rect 5901 4251 5967 4254
rect 7189 4251 7255 4254
rect 3601 4178 3667 4181
rect 6361 4178 6427 4181
rect 3601 4176 6427 4178
rect 3601 4120 3606 4176
rect 3662 4120 6366 4176
rect 6422 4120 6427 4176
rect 3601 4118 6427 4120
rect 3601 4115 3667 4118
rect 6361 4115 6427 4118
rect 17677 4178 17743 4181
rect 22686 4178 22692 4180
rect 17677 4176 22692 4178
rect 17677 4120 17682 4176
rect 17738 4120 22692 4176
rect 17677 4118 22692 4120
rect 17677 4115 17743 4118
rect 22686 4116 22692 4118
rect 22756 4116 22762 4180
rect 3785 4042 3851 4045
rect 5809 4042 5875 4045
rect 8937 4044 9003 4045
rect 5942 4042 5948 4044
rect 3785 4040 5642 4042
rect 3785 3984 3790 4040
rect 3846 3984 5642 4040
rect 3785 3982 5642 3984
rect 3785 3979 3851 3982
rect 4210 3840 4526 3841
rect 0 3680 800 3800
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 5582 3770 5642 3982
rect 5809 4040 5948 4042
rect 5809 3984 5814 4040
rect 5870 3984 5948 4040
rect 5809 3982 5948 3984
rect 5809 3979 5875 3982
rect 5942 3980 5948 3982
rect 6012 3980 6018 4044
rect 8886 4042 8892 4044
rect 8846 3982 8892 4042
rect 8956 4040 9003 4044
rect 8998 3984 9003 4040
rect 8886 3980 8892 3982
rect 8956 3980 9003 3984
rect 9622 3980 9628 4044
rect 9692 4042 9698 4044
rect 10041 4042 10107 4045
rect 16389 4042 16455 4045
rect 9692 4040 16455 4042
rect 9692 3984 10046 4040
rect 10102 3984 16394 4040
rect 16450 3984 16455 4040
rect 9692 3982 16455 3984
rect 9692 3980 9698 3982
rect 8937 3979 9003 3980
rect 10041 3979 10107 3982
rect 16389 3979 16455 3982
rect 17125 4042 17191 4045
rect 17350 4042 17356 4044
rect 17125 4040 17356 4042
rect 17125 3984 17130 4040
rect 17186 3984 17356 4040
rect 17125 3982 17356 3984
rect 17125 3979 17191 3982
rect 17350 3980 17356 3982
rect 17420 3980 17426 4044
rect 18137 4042 18203 4045
rect 18270 4042 18276 4044
rect 18137 4040 18276 4042
rect 18137 3984 18142 4040
rect 18198 3984 18276 4040
rect 18137 3982 18276 3984
rect 18137 3979 18203 3982
rect 18270 3980 18276 3982
rect 18340 3980 18346 4044
rect 18454 3980 18460 4044
rect 18524 4042 18530 4044
rect 18597 4042 18663 4045
rect 18524 4040 18663 4042
rect 18524 3984 18602 4040
rect 18658 3984 18663 4040
rect 18524 3982 18663 3984
rect 18524 3980 18530 3982
rect 18597 3979 18663 3982
rect 20989 4042 21055 4045
rect 21214 4042 21220 4044
rect 20989 4040 21220 4042
rect 20989 3984 20994 4040
rect 21050 3984 21220 4040
rect 20989 3982 21220 3984
rect 20989 3979 21055 3982
rect 21214 3980 21220 3982
rect 21284 3980 21290 4044
rect 6729 3906 6795 3909
rect 12893 3906 12959 3909
rect 6729 3904 12959 3906
rect 6729 3848 6734 3904
rect 6790 3848 12898 3904
rect 12954 3848 12959 3904
rect 6729 3846 12959 3848
rect 6729 3843 6795 3846
rect 12893 3843 12959 3846
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 7649 3770 7715 3773
rect 8293 3772 8359 3773
rect 8293 3770 8340 3772
rect 5582 3768 7715 3770
rect 5582 3712 7654 3768
rect 7710 3712 7715 3768
rect 5582 3710 7715 3712
rect 8248 3768 8340 3770
rect 8404 3770 8410 3772
rect 16113 3770 16179 3773
rect 17769 3772 17835 3773
rect 20345 3772 20411 3773
rect 16430 3770 16436 3772
rect 8248 3712 8298 3768
rect 8248 3710 8340 3712
rect 7649 3707 7715 3710
rect 8293 3708 8340 3710
rect 8404 3710 12450 3770
rect 8404 3708 8410 3710
rect 8293 3707 8359 3708
rect 3233 3634 3299 3637
rect 8477 3634 8543 3637
rect 3233 3632 8543 3634
rect 3233 3576 3238 3632
rect 3294 3576 8482 3632
rect 8538 3576 8543 3632
rect 3233 3574 8543 3576
rect 12390 3634 12450 3710
rect 16113 3768 16436 3770
rect 16113 3712 16118 3768
rect 16174 3712 16436 3768
rect 16113 3710 16436 3712
rect 16113 3707 16179 3710
rect 16430 3708 16436 3710
rect 16500 3708 16506 3772
rect 17718 3708 17724 3772
rect 17788 3770 17835 3772
rect 17788 3768 17880 3770
rect 17830 3712 17880 3768
rect 17788 3710 17880 3712
rect 17788 3708 17835 3710
rect 20294 3708 20300 3772
rect 20364 3770 20411 3772
rect 20364 3768 20456 3770
rect 20406 3712 20456 3768
rect 20364 3710 20456 3712
rect 20364 3708 20411 3710
rect 17769 3707 17835 3708
rect 20345 3707 20411 3708
rect 29913 3634 29979 3637
rect 12390 3632 29979 3634
rect 12390 3576 29918 3632
rect 29974 3576 29979 3632
rect 12390 3574 29979 3576
rect 3233 3571 3299 3574
rect 8477 3571 8543 3574
rect 29913 3571 29979 3574
rect 5533 3498 5599 3501
rect 20253 3498 20319 3501
rect 5533 3496 20319 3498
rect 5533 3440 5538 3496
rect 5594 3440 20258 3496
rect 20314 3440 20319 3496
rect 5533 3438 20319 3440
rect 5533 3435 5599 3438
rect 20253 3435 20319 3438
rect 58157 3498 58223 3501
rect 59200 3498 60000 3528
rect 58157 3496 60000 3498
rect 58157 3440 58162 3496
rect 58218 3440 60000 3496
rect 58157 3438 60000 3440
rect 58157 3435 58223 3438
rect 59200 3408 60000 3438
rect 5901 3362 5967 3365
rect 14089 3362 14155 3365
rect 5901 3360 14155 3362
rect 5901 3304 5906 3360
rect 5962 3304 14094 3360
rect 14150 3304 14155 3360
rect 5901 3302 14155 3304
rect 5901 3299 5967 3302
rect 14089 3299 14155 3302
rect 20345 3362 20411 3365
rect 20478 3362 20484 3364
rect 20345 3360 20484 3362
rect 20345 3304 20350 3360
rect 20406 3304 20484 3360
rect 20345 3302 20484 3304
rect 20345 3299 20411 3302
rect 20478 3300 20484 3302
rect 20548 3300 20554 3364
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 2037 3226 2103 3229
rect 6729 3226 6795 3229
rect 10869 3228 10935 3229
rect 10869 3226 10916 3228
rect 2037 3224 6795 3226
rect 2037 3168 2042 3224
rect 2098 3168 6734 3224
rect 6790 3168 6795 3224
rect 2037 3166 6795 3168
rect 10824 3224 10916 3226
rect 10824 3168 10874 3224
rect 10824 3166 10916 3168
rect 2037 3163 2103 3166
rect 6729 3163 6795 3166
rect 10869 3164 10916 3166
rect 10980 3164 10986 3228
rect 14549 3226 14615 3229
rect 16113 3228 16179 3229
rect 14774 3226 14780 3228
rect 14549 3224 14780 3226
rect 14549 3168 14554 3224
rect 14610 3168 14780 3224
rect 14549 3166 14780 3168
rect 10869 3163 10935 3164
rect 14549 3163 14615 3166
rect 14774 3164 14780 3166
rect 14844 3164 14850 3228
rect 16062 3164 16068 3228
rect 16132 3226 16179 3228
rect 16132 3224 16224 3226
rect 16174 3168 16224 3224
rect 16132 3166 16224 3168
rect 16132 3164 16179 3166
rect 17166 3164 17172 3228
rect 17236 3226 17242 3228
rect 18781 3226 18847 3229
rect 19425 3228 19491 3229
rect 19374 3226 19380 3228
rect 17236 3224 18847 3226
rect 17236 3168 18786 3224
rect 18842 3168 18847 3224
rect 17236 3166 18847 3168
rect 19334 3166 19380 3226
rect 19444 3224 19491 3228
rect 19486 3168 19491 3224
rect 17236 3164 17242 3166
rect 16113 3163 16179 3164
rect 18781 3163 18847 3166
rect 19374 3164 19380 3166
rect 19444 3164 19491 3168
rect 19425 3163 19491 3164
rect 20529 3224 20595 3229
rect 20529 3168 20534 3224
rect 20590 3168 20595 3224
rect 20529 3163 20595 3168
rect 3141 3090 3207 3093
rect 7833 3090 7899 3093
rect 3141 3088 7899 3090
rect 3141 3032 3146 3088
rect 3202 3032 7838 3088
rect 7894 3032 7899 3088
rect 3141 3030 7899 3032
rect 3141 3027 3207 3030
rect 7833 3027 7899 3030
rect 19517 3090 19583 3093
rect 20532 3090 20592 3163
rect 19517 3088 20592 3090
rect 19517 3032 19522 3088
rect 19578 3032 20592 3088
rect 19517 3030 20592 3032
rect 19517 3027 19583 3030
rect 1761 2954 1827 2957
rect 6085 2954 6151 2957
rect 1761 2952 6151 2954
rect 1761 2896 1766 2952
rect 1822 2896 6090 2952
rect 6146 2896 6151 2952
rect 1761 2894 6151 2896
rect 1761 2891 1827 2894
rect 6085 2891 6151 2894
rect 53373 2954 53439 2957
rect 56593 2954 56659 2957
rect 53373 2952 56659 2954
rect 53373 2896 53378 2952
rect 53434 2896 56598 2952
rect 56654 2896 56659 2952
rect 53373 2894 56659 2896
rect 53373 2891 53439 2894
rect 56593 2891 56659 2894
rect 4889 2818 4955 2821
rect 5809 2818 5875 2821
rect 4889 2816 5875 2818
rect 4889 2760 4894 2816
rect 4950 2760 5814 2816
rect 5870 2760 5875 2816
rect 4889 2758 5875 2760
rect 4889 2755 4955 2758
rect 5809 2755 5875 2758
rect 53465 2818 53531 2821
rect 55305 2818 55371 2821
rect 53465 2816 55371 2818
rect 53465 2760 53470 2816
rect 53526 2760 55310 2816
rect 55366 2760 55371 2816
rect 53465 2758 55371 2760
rect 53465 2755 53531 2758
rect 55305 2755 55371 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 3233 2682 3299 2685
rect 10409 2684 10475 2685
rect 3366 2682 3372 2684
rect 3233 2680 3372 2682
rect 3233 2624 3238 2680
rect 3294 2624 3372 2680
rect 3233 2622 3372 2624
rect 3233 2619 3299 2622
rect 3366 2620 3372 2622
rect 3436 2620 3442 2684
rect 10358 2620 10364 2684
rect 10428 2682 10475 2684
rect 13445 2684 13511 2685
rect 14549 2684 14615 2685
rect 13445 2682 13492 2684
rect 10428 2680 10520 2682
rect 10470 2624 10520 2680
rect 10428 2622 10520 2624
rect 13400 2680 13492 2682
rect 13400 2624 13450 2680
rect 13400 2622 13492 2624
rect 10428 2620 10475 2622
rect 10409 2619 10475 2620
rect 13445 2620 13492 2622
rect 13556 2620 13562 2684
rect 14549 2682 14596 2684
rect 14504 2680 14596 2682
rect 14504 2624 14554 2680
rect 14504 2622 14596 2624
rect 14549 2620 14596 2622
rect 14660 2620 14666 2684
rect 16246 2620 16252 2684
rect 16316 2682 16322 2684
rect 18045 2682 18111 2685
rect 16316 2680 18111 2682
rect 16316 2624 18050 2680
rect 18106 2624 18111 2680
rect 16316 2622 18111 2624
rect 16316 2620 16322 2622
rect 13445 2619 13511 2620
rect 14549 2619 14615 2620
rect 18045 2619 18111 2622
rect 18638 2620 18644 2684
rect 18708 2682 18714 2684
rect 20161 2682 20227 2685
rect 18708 2680 20227 2682
rect 18708 2624 20166 2680
rect 20222 2624 20227 2680
rect 18708 2622 20227 2624
rect 18708 2620 18714 2622
rect 20161 2619 20227 2622
rect 0 2184 800 2304
rect 6494 2212 6500 2276
rect 6564 2274 6570 2276
rect 6729 2274 6795 2277
rect 6564 2272 6795 2274
rect 6564 2216 6734 2272
rect 6790 2216 6795 2272
rect 6564 2214 6795 2216
rect 6564 2212 6570 2214
rect 6729 2211 6795 2214
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 57513 2138 57579 2141
rect 59200 2138 60000 2168
rect 57513 2136 60000 2138
rect 57513 2080 57518 2136
rect 57574 2080 60000 2136
rect 57513 2078 60000 2080
rect 57513 2075 57579 2078
rect 59200 2048 60000 2078
rect 6085 1322 6151 1325
rect 6269 1322 6335 1325
rect 6085 1320 6335 1322
rect 6085 1264 6090 1320
rect 6146 1264 6274 1320
rect 6330 1264 6335 1320
rect 6085 1262 6335 1264
rect 6085 1259 6151 1262
rect 6269 1259 6335 1262
rect 58433 778 58499 781
rect 59200 778 60000 808
rect 58433 776 60000 778
rect 58433 720 58438 776
rect 58494 720 60000 776
rect 58433 718 60000 720
rect 58433 715 58499 718
rect 59200 688 60000 718
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 20484 57156 20548 57220
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 18644 56748 18708 56812
rect 21404 56612 21468 56676
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 16252 55584 16316 55588
rect 16252 55528 16266 55584
rect 16266 55528 16316 55584
rect 16252 55524 16316 55528
rect 18276 55524 18340 55588
rect 20300 55584 20364 55588
rect 20300 55528 20350 55584
rect 20350 55528 20364 55584
rect 20300 55524 20364 55528
rect 22692 55524 22756 55588
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 17172 55312 17236 55316
rect 17172 55256 17186 55312
rect 17186 55256 17236 55312
rect 17172 55252 17236 55256
rect 18460 55252 18524 55316
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 13492 53076 13556 53140
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 16436 50220 16500 50284
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 14780 44916 14844 44980
rect 14596 44780 14660 44844
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 17356 42060 17420 42124
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19380 37300 19444 37364
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 22508 35940 22572 36004
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 21956 29004 22020 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 22508 24848 22572 24852
rect 22508 24792 22558 24848
rect 22558 24792 22572 24848
rect 22508 24788 22572 24792
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 21956 22264 22020 22268
rect 21956 22208 22006 22264
rect 22006 22208 22020 22264
rect 21956 22204 22020 22208
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 5948 14724 6012 14788
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 6500 14180 6564 14244
rect 8892 14180 8956 14244
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 21220 13636 21284 13700
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 8340 12548 8404 12612
rect 17724 12548 17788 12612
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 3372 11596 3436 11660
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 16068 9964 16132 10028
rect 21404 9964 21468 10028
rect 10364 9888 10428 9892
rect 10364 9832 10378 9888
rect 10378 9832 10428 9888
rect 10364 9828 10428 9832
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 10916 8196 10980 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 9628 7516 9692 7580
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 22692 4116 22756 4180
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 5948 3980 6012 4044
rect 8892 4040 8956 4044
rect 8892 3984 8942 4040
rect 8942 3984 8956 4040
rect 8892 3980 8956 3984
rect 9628 3980 9692 4044
rect 17356 3980 17420 4044
rect 18276 3980 18340 4044
rect 18460 3980 18524 4044
rect 21220 3980 21284 4044
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 8340 3768 8404 3772
rect 8340 3712 8354 3768
rect 8354 3712 8404 3768
rect 8340 3708 8404 3712
rect 16436 3708 16500 3772
rect 17724 3768 17788 3772
rect 17724 3712 17774 3768
rect 17774 3712 17788 3768
rect 17724 3708 17788 3712
rect 20300 3768 20364 3772
rect 20300 3712 20350 3768
rect 20350 3712 20364 3768
rect 20300 3708 20364 3712
rect 20484 3300 20548 3364
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 10916 3224 10980 3228
rect 10916 3168 10930 3224
rect 10930 3168 10980 3224
rect 10916 3164 10980 3168
rect 14780 3164 14844 3228
rect 16068 3224 16132 3228
rect 16068 3168 16118 3224
rect 16118 3168 16132 3224
rect 16068 3164 16132 3168
rect 17172 3164 17236 3228
rect 19380 3224 19444 3228
rect 19380 3168 19430 3224
rect 19430 3168 19444 3224
rect 19380 3164 19444 3168
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 3372 2620 3436 2684
rect 10364 2680 10428 2684
rect 10364 2624 10414 2680
rect 10414 2624 10428 2680
rect 10364 2620 10428 2624
rect 13492 2680 13556 2684
rect 13492 2624 13506 2680
rect 13506 2624 13556 2680
rect 13492 2620 13556 2624
rect 14596 2680 14660 2684
rect 14596 2624 14610 2680
rect 14610 2624 14660 2680
rect 14596 2620 14660 2624
rect 16252 2620 16316 2684
rect 18644 2620 18708 2684
rect 6500 2212 6564 2276
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 18643 56812 18709 56813
rect 18643 56748 18644 56812
rect 18708 56748 18709 56812
rect 18643 56747 18709 56748
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 16251 55588 16317 55589
rect 16251 55524 16252 55588
rect 16316 55524 16317 55588
rect 16251 55523 16317 55524
rect 18275 55588 18341 55589
rect 18275 55524 18276 55588
rect 18340 55524 18341 55588
rect 18275 55523 18341 55524
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 13491 53140 13557 53141
rect 13491 53076 13492 53140
rect 13556 53076 13557 53140
rect 13491 53075 13557 53076
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 5947 14788 6013 14789
rect 5947 14724 5948 14788
rect 6012 14724 6013 14788
rect 5947 14723 6013 14724
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 3371 11660 3437 11661
rect 3371 11596 3372 11660
rect 3436 11596 3437 11660
rect 3371 11595 3437 11596
rect 3374 2685 3434 11595
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 5950 4045 6010 14723
rect 6499 14244 6565 14245
rect 6499 14180 6500 14244
rect 6564 14180 6565 14244
rect 6499 14179 6565 14180
rect 8891 14244 8957 14245
rect 8891 14180 8892 14244
rect 8956 14180 8957 14244
rect 8891 14179 8957 14180
rect 5947 4044 6013 4045
rect 5947 3980 5948 4044
rect 6012 3980 6013 4044
rect 5947 3979 6013 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 3371 2684 3437 2685
rect 3371 2620 3372 2684
rect 3436 2620 3437 2684
rect 3371 2619 3437 2620
rect 4208 2128 4528 2688
rect 6502 2277 6562 14179
rect 8339 12612 8405 12613
rect 8339 12548 8340 12612
rect 8404 12548 8405 12612
rect 8339 12547 8405 12548
rect 8342 3773 8402 12547
rect 8894 4045 8954 14179
rect 10363 9892 10429 9893
rect 10363 9828 10364 9892
rect 10428 9828 10429 9892
rect 10363 9827 10429 9828
rect 9627 7580 9693 7581
rect 9627 7516 9628 7580
rect 9692 7516 9693 7580
rect 9627 7515 9693 7516
rect 9630 4045 9690 7515
rect 8891 4044 8957 4045
rect 8891 3980 8892 4044
rect 8956 3980 8957 4044
rect 8891 3979 8957 3980
rect 9627 4044 9693 4045
rect 9627 3980 9628 4044
rect 9692 3980 9693 4044
rect 9627 3979 9693 3980
rect 8339 3772 8405 3773
rect 8339 3708 8340 3772
rect 8404 3708 8405 3772
rect 8339 3707 8405 3708
rect 10366 2685 10426 9827
rect 10915 8260 10981 8261
rect 10915 8196 10916 8260
rect 10980 8196 10981 8260
rect 10915 8195 10981 8196
rect 10918 3229 10978 8195
rect 10915 3228 10981 3229
rect 10915 3164 10916 3228
rect 10980 3164 10981 3228
rect 10915 3163 10981 3164
rect 13494 2685 13554 53075
rect 14779 44980 14845 44981
rect 14779 44916 14780 44980
rect 14844 44916 14845 44980
rect 14779 44915 14845 44916
rect 14595 44844 14661 44845
rect 14595 44780 14596 44844
rect 14660 44780 14661 44844
rect 14595 44779 14661 44780
rect 14598 2685 14658 44779
rect 14782 3229 14842 44915
rect 16067 10028 16133 10029
rect 16067 9964 16068 10028
rect 16132 9964 16133 10028
rect 16067 9963 16133 9964
rect 16070 3229 16130 9963
rect 14779 3228 14845 3229
rect 14779 3164 14780 3228
rect 14844 3164 14845 3228
rect 14779 3163 14845 3164
rect 16067 3228 16133 3229
rect 16067 3164 16068 3228
rect 16132 3164 16133 3228
rect 16067 3163 16133 3164
rect 16254 2685 16314 55523
rect 17171 55316 17237 55317
rect 17171 55252 17172 55316
rect 17236 55252 17237 55316
rect 17171 55251 17237 55252
rect 16435 50284 16501 50285
rect 16435 50220 16436 50284
rect 16500 50220 16501 50284
rect 16435 50219 16501 50220
rect 16438 3773 16498 50219
rect 16435 3772 16501 3773
rect 16435 3708 16436 3772
rect 16500 3708 16501 3772
rect 16435 3707 16501 3708
rect 17174 3229 17234 55251
rect 17355 42124 17421 42125
rect 17355 42060 17356 42124
rect 17420 42060 17421 42124
rect 17355 42059 17421 42060
rect 17358 4045 17418 42059
rect 17723 12612 17789 12613
rect 17723 12548 17724 12612
rect 17788 12548 17789 12612
rect 17723 12547 17789 12548
rect 17355 4044 17421 4045
rect 17355 3980 17356 4044
rect 17420 3980 17421 4044
rect 17355 3979 17421 3980
rect 17726 3773 17786 12547
rect 18278 4045 18338 55523
rect 18459 55316 18525 55317
rect 18459 55252 18460 55316
rect 18524 55252 18525 55316
rect 18459 55251 18525 55252
rect 18462 4045 18522 55251
rect 18275 4044 18341 4045
rect 18275 3980 18276 4044
rect 18340 3980 18341 4044
rect 18275 3979 18341 3980
rect 18459 4044 18525 4045
rect 18459 3980 18460 4044
rect 18524 3980 18525 4044
rect 18459 3979 18525 3980
rect 17723 3772 17789 3773
rect 17723 3708 17724 3772
rect 17788 3708 17789 3772
rect 17723 3707 17789 3708
rect 17171 3228 17237 3229
rect 17171 3164 17172 3228
rect 17236 3164 17237 3228
rect 17171 3163 17237 3164
rect 18646 2685 18706 56747
rect 19568 56608 19888 57632
rect 20483 57220 20549 57221
rect 20483 57156 20484 57220
rect 20548 57156 20549 57220
rect 20483 57155 20549 57156
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 20299 55588 20365 55589
rect 20299 55524 20300 55588
rect 20364 55524 20365 55588
rect 20299 55523 20365 55524
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19379 37364 19445 37365
rect 19379 37300 19380 37364
rect 19444 37300 19445 37364
rect 19379 37299 19445 37300
rect 19382 3229 19442 37299
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 20302 3773 20362 55523
rect 20299 3772 20365 3773
rect 20299 3708 20300 3772
rect 20364 3708 20365 3772
rect 20299 3707 20365 3708
rect 20486 3365 20546 57155
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 21403 56676 21469 56677
rect 21403 56612 21404 56676
rect 21468 56612 21469 56676
rect 21403 56611 21469 56612
rect 21219 13700 21285 13701
rect 21219 13636 21220 13700
rect 21284 13636 21285 13700
rect 21219 13635 21285 13636
rect 21222 4045 21282 13635
rect 21406 10029 21466 56611
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 22691 55588 22757 55589
rect 22691 55524 22692 55588
rect 22756 55524 22757 55588
rect 22691 55523 22757 55524
rect 22507 36004 22573 36005
rect 22507 35940 22508 36004
rect 22572 35940 22573 36004
rect 22507 35939 22573 35940
rect 21955 29068 22021 29069
rect 21955 29004 21956 29068
rect 22020 29004 22021 29068
rect 21955 29003 22021 29004
rect 21958 22269 22018 29003
rect 22510 24853 22570 35939
rect 22507 24852 22573 24853
rect 22507 24788 22508 24852
rect 22572 24788 22573 24852
rect 22507 24787 22573 24788
rect 21955 22268 22021 22269
rect 21955 22204 21956 22268
rect 22020 22204 22021 22268
rect 21955 22203 22021 22204
rect 21403 10028 21469 10029
rect 21403 9964 21404 10028
rect 21468 9964 21469 10028
rect 21403 9963 21469 9964
rect 22694 4181 22754 55523
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 22691 4180 22757 4181
rect 22691 4116 22692 4180
rect 22756 4116 22757 4180
rect 22691 4115 22757 4116
rect 21219 4044 21285 4045
rect 21219 3980 21220 4044
rect 21284 3980 21285 4044
rect 21219 3979 21285 3980
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 20483 3364 20549 3365
rect 20483 3300 20484 3364
rect 20548 3300 20549 3364
rect 20483 3299 20549 3300
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19379 3228 19445 3229
rect 19379 3164 19380 3228
rect 19444 3164 19445 3228
rect 19379 3163 19445 3164
rect 10363 2684 10429 2685
rect 10363 2620 10364 2684
rect 10428 2620 10429 2684
rect 10363 2619 10429 2620
rect 13491 2684 13557 2685
rect 13491 2620 13492 2684
rect 13556 2620 13557 2684
rect 13491 2619 13557 2620
rect 14595 2684 14661 2685
rect 14595 2620 14596 2684
rect 14660 2620 14661 2684
rect 14595 2619 14661 2620
rect 16251 2684 16317 2685
rect 16251 2620 16252 2684
rect 16316 2620 16317 2684
rect 16251 2619 16317 2620
rect 18643 2684 18709 2685
rect 18643 2620 18644 2684
rect 18708 2620 18709 2684
rect 18643 2619 18709 2620
rect 6499 2276 6565 2277
rect 6499 2212 6500 2276
rect 6564 2212 6565 2276
rect 6499 2211 6565 2212
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A0
timestamp 1649977179
transform -1 0 3312 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A0
timestamp 1649977179
transform 1 0 5796 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A0
timestamp 1649977179
transform 1 0 4232 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A0
timestamp 1649977179
transform 1 0 5520 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A0
timestamp 1649977179
transform 1 0 5060 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A0
timestamp 1649977179
transform 1 0 5704 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A0
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A0
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A0
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A0
timestamp 1649977179
transform 1 0 12420 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A0
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A0
timestamp 1649977179
transform 1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A
timestamp 1649977179
transform -1 0 6256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A
timestamp 1649977179
transform 1 0 17296 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A
timestamp 1649977179
transform -1 0 12604 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B
timestamp 1649977179
transform -1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1649977179
transform -1 0 7636 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1649977179
transform 1 0 12328 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A1
timestamp 1649977179
transform -1 0 5336 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1649977179
transform -1 0 6808 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1649977179
transform 1 0 4968 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1649977179
transform 1 0 6716 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A1
timestamp 1649977179
transform -1 0 4416 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A
timestamp 1649977179
transform 1 0 8188 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A1
timestamp 1649977179
transform -1 0 5888 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A
timestamp 1649977179
transform -1 0 9936 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1649977179
transform -1 0 7268 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A
timestamp 1649977179
transform -1 0 25116 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1649977179
transform -1 0 12328 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A1
timestamp 1649977179
transform 1 0 13892 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A1
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1649977179
transform 1 0 26312 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A1
timestamp 1649977179
transform -1 0 16744 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1649977179
transform -1 0 23920 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A1
timestamp 1649977179
transform -1 0 15732 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1649977179
transform 1 0 23552 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A1
timestamp 1649977179
transform -1 0 14260 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1649977179
transform 1 0 16468 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1649977179
transform 1 0 12512 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A1
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__C1
timestamp 1649977179
transform 1 0 13984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1649977179
transform 1 0 12880 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A1
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__C1
timestamp 1649977179
transform -1 0 13616 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1649977179
transform -1 0 20700 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B
timestamp 1649977179
transform -1 0 20148 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A
timestamp 1649977179
transform -1 0 29072 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1649977179
transform 1 0 29440 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1649977179
transform -1 0 31556 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A1
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__C1
timestamp 1649977179
transform 1 0 28888 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A1
timestamp 1649977179
transform 1 0 27140 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__C1
timestamp 1649977179
transform 1 0 27324 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1649977179
transform 1 0 27140 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__C1
timestamp 1649977179
transform 1 0 27048 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A
timestamp 1649977179
transform 1 0 29716 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1
timestamp 1649977179
transform 1 0 29716 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1
timestamp 1649977179
transform 1 0 29716 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A1
timestamp 1649977179
transform 1 0 35512 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A1
timestamp 1649977179
transform -1 0 37168 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A1
timestamp 1649977179
transform 1 0 35328 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1649977179
transform -1 0 36800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A1
timestamp 1649977179
transform -1 0 36156 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A1
timestamp 1649977179
transform 1 0 33764 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A1
timestamp 1649977179
transform 1 0 32200 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1649977179
transform -1 0 21252 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B
timestamp 1649977179
transform 1 0 20700 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1649977179
transform -1 0 29716 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1649977179
transform -1 0 31372 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A
timestamp 1649977179
transform 1 0 29440 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A1
timestamp 1649977179
transform 1 0 27876 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A
timestamp 1649977179
transform 1 0 30544 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A1
timestamp 1649977179
transform 1 0 28152 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A1
timestamp 1649977179
transform 1 0 26680 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A1
timestamp 1649977179
transform 1 0 29808 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A1
timestamp 1649977179
transform 1 0 30268 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A1
timestamp 1649977179
transform 1 0 31464 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1649977179
transform 1 0 31280 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A1
timestamp 1649977179
transform 1 0 34500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A1
timestamp 1649977179
transform 1 0 33212 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A1
timestamp 1649977179
transform 1 0 33764 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A1
timestamp 1649977179
transform 1 0 33672 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A1
timestamp 1649977179
transform -1 0 31556 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1649977179
transform 1 0 30452 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A1
timestamp 1649977179
transform 1 0 31464 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__C1
timestamp 1649977179
transform 1 0 29624 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A
timestamp 1649977179
transform 1 0 10856 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A
timestamp 1649977179
transform 1 0 17112 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1
timestamp 1649977179
transform 1 0 5060 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__C1
timestamp 1649977179
transform 1 0 6532 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A1
timestamp 1649977179
transform 1 0 5428 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__C1
timestamp 1649977179
transform -1 0 5060 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A1
timestamp 1649977179
transform -1 0 2208 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C1
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A1
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__C1
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A
timestamp 1649977179
transform 1 0 19688 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1649977179
transform 1 0 7544 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__C1
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A1
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__C1
timestamp 1649977179
transform 1 0 19780 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A1
timestamp 1649977179
transform 1 0 21160 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__C1
timestamp 1649977179
transform -1 0 20240 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1649977179
transform 1 0 20516 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__C1
timestamp 1649977179
transform 1 0 18584 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A1
timestamp 1649977179
transform 1 0 20976 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__C1
timestamp 1649977179
transform 1 0 19688 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A1
timestamp 1649977179
transform 1 0 19780 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A1
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A1
timestamp 1649977179
transform 1 0 14352 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1649977179
transform 1 0 19320 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__B
timestamp 1649977179
transform -1 0 18492 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1649977179
transform 1 0 16744 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1649977179
transform -1 0 16468 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1649977179
transform 1 0 8280 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A1
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1649977179
transform 1 0 23552 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A1
timestamp 1649977179
transform 1 0 11040 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__C1
timestamp 1649977179
transform -1 0 12144 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A1
timestamp 1649977179
transform 1 0 12512 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__C1
timestamp 1649977179
transform 1 0 13432 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1649977179
transform 1 0 14628 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__C1
timestamp 1649977179
transform 1 0 15456 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A1
timestamp 1649977179
transform 1 0 26036 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__C1
timestamp 1649977179
transform -1 0 27508 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A1
timestamp 1649977179
transform 1 0 25300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__C1
timestamp 1649977179
transform 1 0 24380 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A
timestamp 1649977179
transform 1 0 23920 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A1
timestamp 1649977179
transform 1 0 25944 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A1
timestamp 1649977179
transform 1 0 25484 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1649977179
transform 1 0 23736 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A1
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A1
timestamp 1649977179
transform 1 0 23736 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1649977179
transform 1 0 15732 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1649977179
transform 1 0 20700 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A
timestamp 1649977179
transform 1 0 20884 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1649977179
transform -1 0 23000 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1649977179
transform 1 0 23276 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A
timestamp 1649977179
transform -1 0 24104 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A1
timestamp 1649977179
transform 1 0 23276 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A
timestamp 1649977179
transform 1 0 14536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A1
timestamp 1649977179
transform -1 0 24288 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A1
timestamp 1649977179
transform -1 0 23276 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A1
timestamp 1649977179
transform -1 0 24564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A
timestamp 1649977179
transform 1 0 18952 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A1
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1649977179
transform 1 0 28336 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1649977179
transform 1 0 33856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A1
timestamp 1649977179
transform -1 0 30728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1649977179
transform 1 0 30544 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A1
timestamp 1649977179
transform -1 0 32292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1649977179
transform 1 0 28888 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A1
timestamp 1649977179
transform 1 0 29992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A
timestamp 1649977179
transform 1 0 26864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A1
timestamp 1649977179
transform -1 0 31648 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1649977179
transform 1 0 26496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A1
timestamp 1649977179
transform 1 0 28888 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1649977179
transform 1 0 19320 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A1
timestamp 1649977179
transform 1 0 22356 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A1
timestamp 1649977179
transform -1 0 24748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1649977179
transform 1 0 19228 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__B
timestamp 1649977179
transform 1 0 18584 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1649977179
transform 1 0 19412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A1
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A1
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__A1
timestamp 1649977179
transform -1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A1
timestamp 1649977179
transform 1 0 18584 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__C1
timestamp 1649977179
transform -1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A1
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__C1
timestamp 1649977179
transform -1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A1
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__C1
timestamp 1649977179
transform 1 0 28244 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A1
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__C1
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A1
timestamp 1649977179
transform -1 0 30820 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__C1
timestamp 1649977179
transform -1 0 29072 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A1
timestamp 1649977179
transform -1 0 27232 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__C1
timestamp 1649977179
transform 1 0 28336 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1
timestamp 1649977179
transform -1 0 27968 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__C1
timestamp 1649977179
transform 1 0 27876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__C1
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1
timestamp 1649977179
transform -1 0 20332 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__C1
timestamp 1649977179
transform -1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A
timestamp 1649977179
transform 1 0 21988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B
timestamp 1649977179
transform -1 0 24564 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A
timestamp 1649977179
transform 1 0 33856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A
timestamp 1649977179
transform -1 0 36800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1
timestamp 1649977179
transform 1 0 34684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__C1
timestamp 1649977179
transform 1 0 34776 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A1
timestamp 1649977179
transform -1 0 40020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__C1
timestamp 1649977179
transform 1 0 37996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A1
timestamp 1649977179
transform -1 0 37904 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__C1
timestamp 1649977179
transform 1 0 36248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A1
timestamp 1649977179
transform 1 0 37812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__C1
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A1
timestamp 1649977179
transform 1 0 37536 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__C1
timestamp 1649977179
transform 1 0 38088 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A1
timestamp 1649977179
transform 1 0 35880 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__C1
timestamp 1649977179
transform -1 0 35512 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A
timestamp 1649977179
transform 1 0 33120 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__A1
timestamp 1649977179
transform 1 0 39192 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A1
timestamp 1649977179
transform -1 0 41216 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A1
timestamp 1649977179
transform 1 0 39192 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__A1
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__A1
timestamp 1649977179
transform 1 0 40940 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A1
timestamp 1649977179
transform -1 0 36156 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A
timestamp 1649977179
transform 1 0 21988 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B
timestamp 1649977179
transform 1 0 22172 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A
timestamp 1649977179
transform -1 0 38088 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A
timestamp 1649977179
transform 1 0 34868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A1
timestamp 1649977179
transform -1 0 34500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__A1
timestamp 1649977179
transform 1 0 35972 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A1
timestamp 1649977179
transform 1 0 34408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1
timestamp 1649977179
transform 1 0 37168 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A1
timestamp 1649977179
transform -1 0 40020 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A1
timestamp 1649977179
transform -1 0 37536 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A1
timestamp 1649977179
transform -1 0 40848 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__A1
timestamp 1649977179
transform -1 0 41124 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A1
timestamp 1649977179
transform -1 0 39376 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A1
timestamp 1649977179
transform -1 0 41032 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__C1
timestamp 1649977179
transform -1 0 41860 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1649977179
transform 1 0 38272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__C1
timestamp 1649977179
transform 1 0 38916 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A1
timestamp 1649977179
transform -1 0 35236 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__C1
timestamp 1649977179
transform 1 0 36340 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A
timestamp 1649977179
transform -1 0 23920 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B
timestamp 1649977179
transform -1 0 22080 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__A
timestamp 1649977179
transform -1 0 27784 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A
timestamp 1649977179
transform 1 0 26312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A1
timestamp 1649977179
transform -1 0 26864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__C1
timestamp 1649977179
transform 1 0 28336 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A1
timestamp 1649977179
transform 1 0 26312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__C1
timestamp 1649977179
transform 1 0 28152 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A1
timestamp 1649977179
transform -1 0 29072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A1
timestamp 1649977179
transform 1 0 29348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A1
timestamp 1649977179
transform 1 0 31188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__A1
timestamp 1649977179
transform 1 0 31924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1282__A1
timestamp 1649977179
transform 1 0 32200 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__A
timestamp 1649977179
transform 1 0 23736 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A1
timestamp 1649977179
transform 1 0 32384 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A1
timestamp 1649977179
transform 1 0 32200 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__A1
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__A1
timestamp 1649977179
transform -1 0 27968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__A1
timestamp 1649977179
transform -1 0 26956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1649977179
transform 1 0 5888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__A
timestamp 1649977179
transform 1 0 20700 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__A
timestamp 1649977179
transform 1 0 17112 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B
timestamp 1649977179
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__A
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A
timestamp 1649977179
transform 1 0 7728 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__A
timestamp 1649977179
transform -1 0 15732 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1304__A
timestamp 1649977179
transform 1 0 8004 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__A1
timestamp 1649977179
transform 1 0 4784 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A
timestamp 1649977179
transform 1 0 5704 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A1
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A1
timestamp 1649977179
transform 1 0 3128 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__A
timestamp 1649977179
transform 1 0 7912 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A1
timestamp 1649977179
transform 1 0 8188 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A1
timestamp 1649977179
transform 1 0 6900 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A
timestamp 1649977179
transform 1 0 21160 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__A
timestamp 1649977179
transform 1 0 19688 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__A
timestamp 1649977179
transform -1 0 19872 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 1649977179
transform 1 0 21160 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A1
timestamp 1649977179
transform 1 0 21160 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__A
timestamp 1649977179
transform 1 0 25392 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__A1
timestamp 1649977179
transform -1 0 24104 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1327__A
timestamp 1649977179
transform 1 0 26312 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A1
timestamp 1649977179
transform -1 0 23736 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__A
timestamp 1649977179
transform 1 0 14720 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__A1
timestamp 1649977179
transform 1 0 21528 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A
timestamp 1649977179
transform -1 0 16100 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__A1
timestamp 1649977179
transform -1 0 21160 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A
timestamp 1649977179
transform 1 0 11500 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__B
timestamp 1649977179
transform -1 0 17940 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A
timestamp 1649977179
transform 1 0 20424 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A1
timestamp 1649977179
transform 1 0 16928 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__A2
timestamp 1649977179
transform 1 0 17480 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__C1
timestamp 1649977179
transform 1 0 18124 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A
timestamp 1649977179
transform 1 0 10212 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__B
timestamp 1649977179
transform 1 0 20424 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A1
timestamp 1649977179
transform 1 0 18676 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__A2
timestamp 1649977179
transform -1 0 19136 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__C1
timestamp 1649977179
transform 1 0 19320 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__A
timestamp 1649977179
transform -1 0 22448 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__B
timestamp 1649977179
transform -1 0 22172 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__A
timestamp 1649977179
transform -1 0 22540 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A
timestamp 1649977179
transform 1 0 19688 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__A1
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__C1
timestamp 1649977179
transform 1 0 17296 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__A1
timestamp 1649977179
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__C1
timestamp 1649977179
transform 1 0 18768 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__A1
timestamp 1649977179
transform 1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__C1
timestamp 1649977179
transform -1 0 16192 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__A
timestamp 1649977179
transform 1 0 16100 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__A1
timestamp 1649977179
transform 1 0 15732 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A1
timestamp 1649977179
transform -1 0 18124 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__A1
timestamp 1649977179
transform -1 0 24472 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__A1
timestamp 1649977179
transform -1 0 25392 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__A1
timestamp 1649977179
transform -1 0 27140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__A
timestamp 1649977179
transform -1 0 13524 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__A1
timestamp 1649977179
transform 1 0 24472 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__C1
timestamp 1649977179
transform -1 0 25024 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__A1
timestamp 1649977179
transform -1 0 25024 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__C1
timestamp 1649977179
transform 1 0 24288 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__A1
timestamp 1649977179
transform 1 0 22816 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__C1
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__A1
timestamp 1649977179
transform -1 0 22724 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__C1
timestamp 1649977179
transform -1 0 22172 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__A
timestamp 1649977179
transform -1 0 9752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__B
timestamp 1649977179
transform -1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__A
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__A
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__A1
timestamp 1649977179
transform 1 0 8004 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__C1
timestamp 1649977179
transform 1 0 8924 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__A1
timestamp 1649977179
transform -1 0 2208 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__C1
timestamp 1649977179
transform 1 0 4600 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A1
timestamp 1649977179
transform 1 0 3128 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__C1
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__A1
timestamp 1649977179
transform 1 0 8004 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__C1
timestamp 1649977179
transform -1 0 7636 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__A1
timestamp 1649977179
transform 1 0 6256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__C1
timestamp 1649977179
transform 1 0 8188 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__A1
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__C1
timestamp 1649977179
transform 1 0 13892 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A1
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__A1
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__A1
timestamp 1649977179
transform 1 0 16928 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A1
timestamp 1649977179
transform 1 0 17480 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A1
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A1
timestamp 1649977179
transform 1 0 9752 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A
timestamp 1649977179
transform -1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__B
timestamp 1649977179
transform -1 0 10672 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__A
timestamp 1649977179
transform -1 0 7912 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__A
timestamp 1649977179
transform 1 0 9936 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__A1
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__A1
timestamp 1649977179
transform 1 0 2852 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__A1
timestamp 1649977179
transform -1 0 3312 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__A1
timestamp 1649977179
transform -1 0 5612 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__A1
timestamp 1649977179
transform -1 0 6624 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A1
timestamp 1649977179
transform 1 0 10672 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__A1
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A1
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__A1
timestamp 1649977179
transform 1 0 11960 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__A
timestamp 1649977179
transform 1 0 12328 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__A1
timestamp 1649977179
transform 1 0 11408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__C1
timestamp 1649977179
transform -1 0 12052 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__A1
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__C1
timestamp 1649977179
transform 1 0 10396 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__A1
timestamp 1649977179
transform 1 0 10120 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__C1
timestamp 1649977179
transform 1 0 10672 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__A
timestamp 1649977179
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__B
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__A
timestamp 1649977179
transform -1 0 14628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__A
timestamp 1649977179
transform 1 0 15640 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__A1
timestamp 1649977179
transform 1 0 11316 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__C1
timestamp 1649977179
transform -1 0 13064 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A1
timestamp 1649977179
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__C1
timestamp 1649977179
transform 1 0 11960 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A
timestamp 1649977179
transform 1 0 14260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__A1
timestamp 1649977179
transform 1 0 10764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__A1
timestamp 1649977179
transform -1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__A1
timestamp 1649977179
transform 1 0 12512 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__A1
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__A1
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__A
timestamp 1649977179
transform 1 0 20424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__A1
timestamp 1649977179
transform -1 0 23092 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__A1
timestamp 1649977179
transform 1 0 21252 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__A1
timestamp 1649977179
transform 1 0 17480 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__A1
timestamp 1649977179
transform 1 0 16744 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__A1
timestamp 1649977179
transform 1 0 17940 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__A
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__A
timestamp 1649977179
transform 1 0 21620 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__A
timestamp 1649977179
transform 1 0 20332 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__A
timestamp 1649977179
transform 1 0 15456 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__A1
timestamp 1649977179
transform -1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__A1
timestamp 1649977179
transform 1 0 11960 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__A1
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__A1
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__A1
timestamp 1649977179
transform 1 0 17572 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__A
timestamp 1649977179
transform -1 0 25760 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__A1
timestamp 1649977179
transform 1 0 28980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__A1
timestamp 1649977179
transform 1 0 29808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__A1
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__A1
timestamp 1649977179
transform 1 0 26312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__A1
timestamp 1649977179
transform -1 0 27784 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__A1
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__C1
timestamp 1649977179
transform 1 0 17204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__A1
timestamp 1649977179
transform 1 0 16744 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__C1
timestamp 1649977179
transform 1 0 17756 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1535__D
timestamp 1649977179
transform 1 0 24932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1541__C1
timestamp 1649977179
transform 1 0 8096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1546__D
timestamp 1649977179
transform 1 0 24196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1554__C1
timestamp 1649977179
transform 1 0 6808 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1559__D
timestamp 1649977179
transform -1 0 25668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1564__A
timestamp 1649977179
transform -1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1567__C1
timestamp 1649977179
transform 1 0 7176 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__A
timestamp 1649977179
transform 1 0 30912 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1585__A
timestamp 1649977179
transform -1 0 32292 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__A2
timestamp 1649977179
transform -1 0 16192 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1599__B1
timestamp 1649977179
transform -1 0 15088 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__A
timestamp 1649977179
transform -1 0 8464 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__A2
timestamp 1649977179
transform -1 0 15640 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__B1
timestamp 1649977179
transform 1 0 15824 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1618__A
timestamp 1649977179
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1620__A1
timestamp 1649977179
transform -1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__A2
timestamp 1649977179
transform 1 0 23000 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1629__B1
timestamp 1649977179
transform -1 0 23276 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__A2
timestamp 1649977179
transform -1 0 22724 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__B1
timestamp 1649977179
transform -1 0 23276 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1646__B1
timestamp 1649977179
transform 1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1654__A2
timestamp 1649977179
transform 1 0 22264 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1654__B1
timestamp 1649977179
transform 1 0 22448 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1656__B
timestamp 1649977179
transform 1 0 21528 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1659__B1
timestamp 1649977179
transform -1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1671__B1
timestamp 1649977179
transform 1 0 10120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1695__B1
timestamp 1649977179
transform -1 0 4508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1708__A
timestamp 1649977179
transform -1 0 2760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2167__A
timestamp 1649977179
transform -1 0 46368 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2168__A
timestamp 1649977179
transform 1 0 25392 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2169__A
timestamp 1649977179
transform 1 0 44344 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2170__A
timestamp 1649977179
transform -1 0 19688 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2171__A
timestamp 1649977179
transform -1 0 20148 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2172__A
timestamp 1649977179
transform -1 0 17940 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2173__A
timestamp 1649977179
transform -1 0 18768 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2174__A
timestamp 1649977179
transform -1 0 20884 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2175__A
timestamp 1649977179
transform -1 0 20240 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2176__A
timestamp 1649977179
transform 1 0 24748 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2177__A
timestamp 1649977179
transform -1 0 34776 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2178__A
timestamp 1649977179
transform -1 0 32936 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2179__A
timestamp 1649977179
transform -1 0 30452 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2180__A
timestamp 1649977179
transform -1 0 27968 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2181__A
timestamp 1649977179
transform -1 0 25484 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2182__A
timestamp 1649977179
transform -1 0 27048 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2183__A
timestamp 1649977179
transform -1 0 26680 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2184__A
timestamp 1649977179
transform 1 0 23368 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2185__A
timestamp 1649977179
transform 1 0 22448 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2186__A
timestamp 1649977179
transform 1 0 20884 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2187__A
timestamp 1649977179
transform 1 0 18952 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2188__A
timestamp 1649977179
transform -1 0 18124 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2189__A
timestamp 1649977179
transform -1 0 16836 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2190__A
timestamp 1649977179
transform 1 0 17112 0 -1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2191__A
timestamp 1649977179
transform 1 0 16192 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2192__A
timestamp 1649977179
transform 1 0 14168 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2193__A
timestamp 1649977179
transform -1 0 20516 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2194__A
timestamp 1649977179
transform -1 0 22448 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2195__A
timestamp 1649977179
transform 1 0 30820 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2196__A
timestamp 1649977179
transform -1 0 36616 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 20424 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 10028 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1__f_wb_clk_i_A
timestamp 1649977179
transform -1 0 12512 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2__f_wb_clk_i_A
timestamp 1649977179
transform -1 0 27600 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3__f_wb_clk_i_A
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_wb_clk_i_A
timestamp 1649977179
transform 1 0 12512 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_wb_clk_i_A
timestamp 1649977179
transform -1 0 6532 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_wb_clk_i_A
timestamp 1649977179
transform 1 0 9108 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_wb_clk_i_A
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_wb_clk_i_A
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_wb_clk_i_A
timestamp 1649977179
transform 1 0 11592 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_wb_clk_i_A
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_wb_clk_i_A
timestamp 1649977179
transform 1 0 16928 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_wb_clk_i_A
timestamp 1649977179
transform 1 0 20240 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_wb_clk_i_A
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_wb_clk_i_A
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_wb_clk_i_A
timestamp 1649977179
transform -1 0 29900 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_wb_clk_i_A
timestamp 1649977179
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_wb_clk_i_A
timestamp 1649977179
transform 1 0 34408 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_wb_clk_i_A
timestamp 1649977179
transform 1 0 38548 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_wb_clk_i_A
timestamp 1649977179
transform -1 0 33580 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_wb_clk_i_A
timestamp 1649977179
transform 1 0 30084 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_wb_clk_i_A
timestamp 1649977179
transform 1 0 27876 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_wb_clk_i_A
timestamp 1649977179
transform 1 0 32476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_wb_clk_i_A
timestamp 1649977179
transform 1 0 37536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_wb_clk_i_A
timestamp 1649977179
transform 1 0 36800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_wb_clk_i_A
timestamp 1649977179
transform 1 0 36524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_wb_clk_i_A
timestamp 1649977179
transform -1 0 33764 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_wb_clk_i_A
timestamp 1649977179
transform 1 0 30360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_wb_clk_i_A
timestamp 1649977179
transform 1 0 26864 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_wb_clk_i_A
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_27_wb_clk_i_A
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_28_wb_clk_i_A
timestamp 1649977179
transform 1 0 15732 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_29_wb_clk_i_A
timestamp 1649977179
transform -1 0 16928 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_30_wb_clk_i_A
timestamp 1649977179
transform 1 0 9660 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_31_wb_clk_i_A
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_32_wb_clk_i_A
timestamp 1649977179
transform 1 0 8096 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_33_wb_clk_i_A
timestamp 1649977179
transform 1 0 4416 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_34_wb_clk_i_A
timestamp 1649977179
transform 1 0 9016 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 13064 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 14260 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 25668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 19412 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 19412 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 20056 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 15548 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 19964 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 20792 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 13064 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 20792 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 26220 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 21712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 23828 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 24564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 25116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 22632 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 27140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 24564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 16836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 5520 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 4416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 19964 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 13156 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 20516 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 1656 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 2576 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 11592 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 10488 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 8096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 2024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 1748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 8924 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 3220 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 9292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 3128 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 6072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 1564 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 3956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 1932 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 2668 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 10856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 2208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 2024 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1649977179
transform 1 0 2576 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output87_A
timestamp 1649977179
transform 1 0 42320 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output97_A
timestamp 1649977179
transform -1 0 4048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16
timestamp 1649977179
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_103 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1649977179
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_172
timestamp 1649977179
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_180
timestamp 1649977179
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_188
timestamp 1649977179
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_201
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_207
timestamp 1649977179
transform 1 0 20148 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_212
timestamp 1649977179
transform 1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_230
timestamp 1649977179
transform 1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_238
timestamp 1649977179
transform 1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1649977179
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_255
timestamp 1649977179
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_283
timestamp 1649977179
transform 1 0 27140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_316
timestamp 1649977179
transform 1 0 30176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_323
timestamp 1649977179
transform 1 0 30820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1649977179
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_340
timestamp 1649977179
transform 1 0 32384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1649977179
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_354
timestamp 1649977179
transform 1 0 33672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_362
timestamp 1649977179
transform 1 0 34408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_382
timestamp 1649977179
transform 1 0 36248 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1649977179
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1649977179
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_424
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_446
timestamp 1649977179
transform 1 0 42136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_466
timestamp 1649977179
transform 1 0 43976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_474
timestamp 1649977179
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_494
timestamp 1649977179
transform 1 0 46552 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1649977179
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_522
timestamp 1649977179
transform 1 0 49128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_530
timestamp 1649977179
transform 1 0 49864 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_550
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_558
timestamp 1649977179
transform 1 0 52440 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1649977179
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_578
timestamp 1649977179
transform 1 0 54280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_586
timestamp 1649977179
transform 1 0 55016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_592
timestamp 1649977179
transform 1 0 55568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_599
timestamp 1649977179
transform 1 0 56212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_606
timestamp 1649977179
transform 1 0 56856 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_614
timestamp 1649977179
transform 1 0 57592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_624
timestamp 1649977179
transform 1 0 58512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_10
timestamp 1649977179
transform 1 0 2024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_36
timestamp 1649977179
transform 1 0 4416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_44
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_61
timestamp 1649977179
transform 1 0 6716 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_72
timestamp 1649977179
transform 1 0 7728 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1649977179
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_97
timestamp 1649977179
transform 1 0 10028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1649977179
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_129
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_133
timestamp 1649977179
transform 1 0 13340 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_140
timestamp 1649977179
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_148
timestamp 1649977179
transform 1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_156
timestamp 1649977179
transform 1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_172
timestamp 1649977179
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_180
timestamp 1649977179
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1649977179
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_196
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_204
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_212
timestamp 1649977179
transform 1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_232
timestamp 1649977179
transform 1 0 22448 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1649977179
transform 1 0 23184 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_244
timestamp 1649977179
transform 1 0 23552 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1649977179
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_285
timestamp 1649977179
transform 1 0 27324 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_289
timestamp 1649977179
transform 1 0 27692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_296
timestamp 1649977179
transform 1 0 28336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_303
timestamp 1649977179
transform 1 0 28980 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_310
timestamp 1649977179
transform 1 0 29624 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_324 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30912 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_340
timestamp 1649977179
transform 1 0 32384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_347
timestamp 1649977179
transform 1 0 33028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_354
timestamp 1649977179
transform 1 0 33672 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_368
timestamp 1649977179
transform 1 0 34960 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_375
timestamp 1649977179
transform 1 0 35604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp 1649977179
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1649977179
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1649977179
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1649977179
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1649977179
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_438
timestamp 1649977179
transform 1 0 41400 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_446
timestamp 1649977179
transform 1 0 42136 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1649977179
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_466
timestamp 1649977179
transform 1 0 43976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_480
timestamp 1649977179
transform 1 0 45264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1649977179
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_494
timestamp 1649977179
transform 1 0 46552 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1649977179
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_515
timestamp 1649977179
transform 1 0 48484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_522
timestamp 1649977179
transform 1 0 49128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_536
timestamp 1649977179
transform 1 0 50416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_543
timestamp 1649977179
transform 1 0 51060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_550
timestamp 1649977179
transform 1 0 51704 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_558
timestamp 1649977179
transform 1 0 52440 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_564
timestamp 1649977179
transform 1 0 52992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_571
timestamp 1649977179
transform 1 0 53636 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_578
timestamp 1649977179
transform 1 0 54280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_585
timestamp 1649977179
transform 1 0 54924 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_592
timestamp 1649977179
transform 1 0 55568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_599
timestamp 1649977179
transform 1 0 56212 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_606
timestamp 1649977179
transform 1 0 56856 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_614
timestamp 1649977179
transform 1 0 57592 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_624
timestamp 1649977179
transform 1 0 58512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1649977179
transform 1 0 5336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_55
timestamp 1649977179
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_69
timestamp 1649977179
transform 1 0 7452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_73
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_104
timestamp 1649977179
transform 1 0 10672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_112
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_118
timestamp 1649977179
transform 1 0 11960 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1649977179
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_129
timestamp 1649977179
transform 1 0 12972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_151
timestamp 1649977179
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_183
timestamp 1649977179
transform 1 0 17940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_187
timestamp 1649977179
transform 1 0 18308 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1649977179
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1649977179
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_214
timestamp 1649977179
transform 1 0 20792 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1649977179
transform 1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_223
timestamp 1649977179
transform 1 0 21620 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_228
timestamp 1649977179
transform 1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1649977179
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1649977179
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1649977179
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_259
timestamp 1649977179
transform 1 0 24932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_266
timestamp 1649977179
transform 1 0 25576 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_273
timestamp 1649977179
transform 1 0 26220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_293
timestamp 1649977179
transform 1 0 28060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_299
timestamp 1649977179
transform 1 0 28612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_303
timestamp 1649977179
transform 1 0 28980 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_341
timestamp 1649977179
transform 1 0 32476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_353
timestamp 1649977179
transform 1 0 33580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_361
timestamp 1649977179
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_369
timestamp 1649977179
transform 1 0 35052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_376
timestamp 1649977179
transform 1 0 35696 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_383
timestamp 1649977179
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_390
timestamp 1649977179
transform 1 0 36984 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_399
timestamp 1649977179
transform 1 0 37812 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_407
timestamp 1649977179
transform 1 0 38548 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_411
timestamp 1649977179
transform 1 0 38916 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1649977179
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_426
timestamp 1649977179
transform 1 0 40296 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_433
timestamp 1649977179
transform 1 0 40940 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_440
timestamp 1649977179
transform 1 0 41584 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_448
timestamp 1649977179
transform 1 0 42320 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_453
timestamp 1649977179
transform 1 0 42780 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_460
timestamp 1649977179
transform 1 0 43424 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1649977179
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_480
timestamp 1649977179
transform 1 0 45264 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_487
timestamp 1649977179
transform 1 0 45908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_494
timestamp 1649977179
transform 1 0 46552 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_510
timestamp 1649977179
transform 1 0 48024 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_517
timestamp 1649977179
transform 1 0 48668 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_529
timestamp 1649977179
transform 1 0 49772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_533
timestamp 1649977179
transform 1 0 50140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_537
timestamp 1649977179
transform 1 0 50508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_544
timestamp 1649977179
transform 1 0 51152 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_551
timestamp 1649977179
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_558
timestamp 1649977179
transform 1 0 52440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_565
timestamp 1649977179
transform 1 0 53084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_572
timestamp 1649977179
transform 1 0 53728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_579
timestamp 1649977179
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_592
timestamp 1649977179
transform 1 0 55568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_599
timestamp 1649977179
transform 1 0 56212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_606
timestamp 1649977179
transform 1 0 56856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_610
timestamp 1649977179
transform 1 0 57224 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_614
timestamp 1649977179
transform 1 0 57592 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1649977179
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_7
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_14
timestamp 1649977179
transform 1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_21
timestamp 1649977179
transform 1 0 3036 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_28
timestamp 1649977179
transform 1 0 3680 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_44
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_52
timestamp 1649977179
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_63
timestamp 1649977179
transform 1 0 6900 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_79
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_88
timestamp 1649977179
transform 1 0 9200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_96
timestamp 1649977179
transform 1 0 9936 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_104
timestamp 1649977179
transform 1 0 10672 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_124
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_132
timestamp 1649977179
transform 1 0 13248 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_136
timestamp 1649977179
transform 1 0 13616 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_143
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_150
timestamp 1649977179
transform 1 0 14904 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_157
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_185
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_191
timestamp 1649977179
transform 1 0 18676 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_195
timestamp 1649977179
transform 1 0 19044 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_215
timestamp 1649977179
transform 1 0 20884 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_232
timestamp 1649977179
transform 1 0 22448 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_239
timestamp 1649977179
transform 1 0 23092 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_246
timestamp 1649977179
transform 1 0 23736 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_255
timestamp 1649977179
transform 1 0 24564 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_263
timestamp 1649977179
transform 1 0 25300 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_267
timestamp 1649977179
transform 1 0 25668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_311
timestamp 1649977179
transform 1 0 29716 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_314
timestamp 1649977179
transform 1 0 29992 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_326
timestamp 1649977179
transform 1 0 31096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_334
timestamp 1649977179
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_383
timestamp 1649977179
transform 1 0 36340 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1649977179
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1649977179
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1649977179
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1649977179
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1649977179
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1649977179
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_517
timestamp 1649977179
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_541
timestamp 1649977179
transform 1 0 50876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_547
timestamp 1649977179
transform 1 0 51428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_554
timestamp 1649977179
transform 1 0 52072 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_564
timestamp 1649977179
transform 1 0 52992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_571
timestamp 1649977179
transform 1 0 53636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_578
timestamp 1649977179
transform 1 0 54280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_585
timestamp 1649977179
transform 1 0 54924 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_592
timestamp 1649977179
transform 1 0 55568 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_599
timestamp 1649977179
transform 1 0 56212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_611
timestamp 1649977179
transform 1 0 57316 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_621
timestamp 1649977179
transform 1 0 58236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_5
timestamp 1649977179
transform 1 0 1564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_11
timestamp 1649977179
transform 1 0 2116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp 1649977179
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_33
timestamp 1649977179
transform 1 0 4140 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_42
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_48
timestamp 1649977179
transform 1 0 5520 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_56
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_64
timestamp 1649977179
transform 1 0 6992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_92
timestamp 1649977179
transform 1 0 9568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_96
timestamp 1649977179
transform 1 0 9936 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_106
timestamp 1649977179
transform 1 0 10856 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_125
timestamp 1649977179
transform 1 0 12604 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1649977179
transform 1 0 12972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_143
timestamp 1649977179
transform 1 0 14260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_150
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_157
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_164
timestamp 1649977179
transform 1 0 16192 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_171
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_178
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_185
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_200
timestamp 1649977179
transform 1 0 19504 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_207
timestamp 1649977179
transform 1 0 20148 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_214
timestamp 1649977179
transform 1 0 20792 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_228
timestamp 1649977179
transform 1 0 22080 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1649977179
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_255
timestamp 1649977179
transform 1 0 24564 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_261
timestamp 1649977179
transform 1 0 25116 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_267
timestamp 1649977179
transform 1 0 25668 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_273
timestamp 1649977179
transform 1 0 26220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_276
timestamp 1649977179
transform 1 0 26496 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_288
timestamp 1649977179
transform 1 0 27600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_300
timestamp 1649977179
transform 1 0 28704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_313
timestamp 1649977179
transform 1 0 29900 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_322
timestamp 1649977179
transform 1 0 30728 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_331
timestamp 1649977179
transform 1 0 31556 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_343
timestamp 1649977179
transform 1 0 32660 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp 1649977179
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1649977179
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1649977179
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1649977179
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1649977179
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1649977179
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1649977179
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1649977179
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_525
timestamp 1649977179
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_531
timestamp 1649977179
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_533
timestamp 1649977179
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_545
timestamp 1649977179
transform 1 0 51244 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_553
timestamp 1649977179
transform 1 0 51980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_558
timestamp 1649977179
transform 1 0 52440 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_565
timestamp 1649977179
transform 1 0 53084 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_572
timestamp 1649977179
transform 1 0 53728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_579
timestamp 1649977179
transform 1 0 54372 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_592
timestamp 1649977179
transform 1 0 55568 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_599
timestamp 1649977179
transform 1 0 56212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_611
timestamp 1649977179
transform 1 0 57316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_623
timestamp 1649977179
transform 1 0 58420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_5
timestamp 1649977179
transform 1 0 1564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_11
timestamp 1649977179
transform 1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_20
timestamp 1649977179
transform 1 0 2944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_28
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_31
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_38
timestamp 1649977179
transform 1 0 4600 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_65
timestamp 1649977179
transform 1 0 7084 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_74
timestamp 1649977179
transform 1 0 7912 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_82
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_90
timestamp 1649977179
transform 1 0 9384 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1649977179
transform 1 0 9752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_101
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_131
timestamp 1649977179
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_138
timestamp 1649977179
transform 1 0 13800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_145
timestamp 1649977179
transform 1 0 14444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_152
timestamp 1649977179
transform 1 0 15088 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1649977179
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1649977179
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1649977179
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_177
timestamp 1649977179
transform 1 0 17388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_189
timestamp 1649977179
transform 1 0 18492 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_5_200
timestamp 1649977179
transform 1 0 19504 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_206
timestamp 1649977179
transform 1 0 20056 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_210
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1649977179
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_228
timestamp 1649977179
transform 1 0 22080 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_245
timestamp 1649977179
transform 1 0 23644 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_262
timestamp 1649977179
transform 1 0 25208 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_268
timestamp 1649977179
transform 1 0 25760 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_289
timestamp 1649977179
transform 1 0 27692 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_295
timestamp 1649977179
transform 1 0 28244 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_307
timestamp 1649977179
transform 1 0 29348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_319
timestamp 1649977179
transform 1 0 30452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_331
timestamp 1649977179
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_355
timestamp 1649977179
transform 1 0 33764 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_379
timestamp 1649977179
transform 1 0 35972 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1649977179
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1649977179
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1649977179
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_517
timestamp 1649977179
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_529
timestamp 1649977179
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_541
timestamp 1649977179
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1649977179
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_561
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_569
timestamp 1649977179
transform 1 0 53452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_575
timestamp 1649977179
transform 1 0 54004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_582
timestamp 1649977179
transform 1 0 54648 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_589
timestamp 1649977179
transform 1 0 55292 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_601
timestamp 1649977179
transform 1 0 56396 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_613
timestamp 1649977179
transform 1 0 57500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_621
timestamp 1649977179
transform 1 0 58236 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_38
timestamp 1649977179
transform 1 0 4600 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_42
timestamp 1649977179
transform 1 0 4968 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_51
timestamp 1649977179
transform 1 0 5796 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_55
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_60
timestamp 1649977179
transform 1 0 6624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_68
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_76
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_92
timestamp 1649977179
transform 1 0 9568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1649977179
transform 1 0 10212 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_106
timestamp 1649977179
transform 1 0 10856 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_114
timestamp 1649977179
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_120
timestamp 1649977179
transform 1 0 12144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_127
timestamp 1649977179
transform 1 0 12788 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_144
timestamp 1649977179
transform 1 0 14352 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_160
timestamp 1649977179
transform 1 0 15824 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_169
timestamp 1649977179
transform 1 0 16652 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_180
timestamp 1649977179
transform 1 0 17664 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_213
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_224
timestamp 1649977179
transform 1 0 21712 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_235
timestamp 1649977179
transform 1 0 22724 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_241
timestamp 1649977179
transform 1 0 23276 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_247
timestamp 1649977179
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_258
timestamp 1649977179
transform 1 0 24840 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_276
timestamp 1649977179
transform 1 0 26496 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_282
timestamp 1649977179
transform 1 0 27048 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_294
timestamp 1649977179
transform 1 0 28152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1649977179
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_311
timestamp 1649977179
transform 1 0 29716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_323
timestamp 1649977179
transform 1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_327
timestamp 1649977179
transform 1 0 31188 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_344
timestamp 1649977179
transform 1 0 32752 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_356
timestamp 1649977179
transform 1 0 33856 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_382
timestamp 1649977179
transform 1 0 36248 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_394
timestamp 1649977179
transform 1 0 37352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_411
timestamp 1649977179
transform 1 0 38916 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1649977179
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1649977179
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1649977179
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1649977179
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1649977179
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1649977179
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1649977179
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_557
timestamp 1649977179
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_569
timestamp 1649977179
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_581
timestamp 1649977179
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_9
timestamp 1649977179
transform 1 0 1932 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_16
timestamp 1649977179
transform 1 0 2576 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_22
timestamp 1649977179
transform 1 0 3128 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_43
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_59
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_66
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_73
timestamp 1649977179
transform 1 0 7820 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_80
timestamp 1649977179
transform 1 0 8464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_87
timestamp 1649977179
transform 1 0 9108 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_91
timestamp 1649977179
transform 1 0 9476 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_124
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_153
timestamp 1649977179
transform 1 0 15180 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_162
timestamp 1649977179
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_172
timestamp 1649977179
transform 1 0 16928 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_196
timestamp 1649977179
transform 1 0 19136 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_211
timestamp 1649977179
transform 1 0 20516 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_214
timestamp 1649977179
transform 1 0 20792 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_235
timestamp 1649977179
transform 1 0 22724 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_246
timestamp 1649977179
transform 1 0 23736 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_252
timestamp 1649977179
transform 1 0 24288 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1649977179
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_284
timestamp 1649977179
transform 1 0 27232 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_290
timestamp 1649977179
transform 1 0 27784 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_302
timestamp 1649977179
transform 1 0 28888 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_326
timestamp 1649977179
transform 1 0 31096 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1649977179
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_364
timestamp 1649977179
transform 1 0 34592 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_376
timestamp 1649977179
transform 1 0 35696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_398
timestamp 1649977179
transform 1 0 37720 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_420
timestamp 1649977179
transform 1 0 39744 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_432
timestamp 1649977179
transform 1 0 40848 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_444
timestamp 1649977179
transform 1 0 41952 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1649977179
transform 1 0 58236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp 1649977179
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_12
timestamp 1649977179
transform 1 0 2208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_18
timestamp 1649977179
transform 1 0 2760 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1649977179
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_31
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_37
timestamp 1649977179
transform 1 0 4508 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_45
timestamp 1649977179
transform 1 0 5244 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_51
timestamp 1649977179
transform 1 0 5796 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_54
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_68
timestamp 1649977179
transform 1 0 7360 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_88
timestamp 1649977179
transform 1 0 9200 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_101
timestamp 1649977179
transform 1 0 10396 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_108
timestamp 1649977179
transform 1 0 11040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_114
timestamp 1649977179
transform 1 0 11592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_122
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_128
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_150
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_158
timestamp 1649977179
transform 1 0 15640 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_172
timestamp 1649977179
transform 1 0 16928 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_178
timestamp 1649977179
transform 1 0 17480 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_181
timestamp 1649977179
transform 1 0 17756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_185
timestamp 1649977179
transform 1 0 18124 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_188
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_199
timestamp 1649977179
transform 1 0 19412 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_203
timestamp 1649977179
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_206
timestamp 1649977179
transform 1 0 20056 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_214
timestamp 1649977179
transform 1 0 20792 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_239
timestamp 1649977179
transform 1 0 23092 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1649977179
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_261
timestamp 1649977179
transform 1 0 25116 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_269
timestamp 1649977179
transform 1 0 25852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_280
timestamp 1649977179
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_292
timestamp 1649977179
transform 1 0 27968 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_329
timestamp 1649977179
transform 1 0 31372 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_341
timestamp 1649977179
transform 1 0 32476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_353
timestamp 1649977179
transform 1 0 33580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_360
timestamp 1649977179
transform 1 0 34224 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_375
timestamp 1649977179
transform 1 0 35604 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_381
timestamp 1649977179
transform 1 0 36156 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_385
timestamp 1649977179
transform 1 0 36524 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_394
timestamp 1649977179
transform 1 0 37352 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_400
timestamp 1649977179
transform 1 0 37904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_404
timestamp 1649977179
transform 1 0 38272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1649977179
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1649977179
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_423
timestamp 1649977179
transform 1 0 40020 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_435
timestamp 1649977179
transform 1 0 41124 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_447
timestamp 1649977179
transform 1 0 42228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_459
timestamp 1649977179
transform 1 0 43332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_471
timestamp 1649977179
transform 1 0 44436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1649977179
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1649977179
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_557
timestamp 1649977179
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_569
timestamp 1649977179
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_581
timestamp 1649977179
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_587
timestamp 1649977179
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_10
timestamp 1649977179
transform 1 0 2024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_16
timestamp 1649977179
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_22
timestamp 1649977179
transform 1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_35
timestamp 1649977179
transform 1 0 4324 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_43
timestamp 1649977179
transform 1 0 5060 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_46
timestamp 1649977179
transform 1 0 5336 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_66
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_78
timestamp 1649977179
transform 1 0 8280 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_82
timestamp 1649977179
transform 1 0 8648 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_85
timestamp 1649977179
transform 1 0 8924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_96
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_102
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_115
timestamp 1649977179
transform 1 0 11684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_139
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_144
timestamp 1649977179
transform 1 0 14352 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_158
timestamp 1649977179
transform 1 0 15640 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_174
timestamp 1649977179
transform 1 0 17112 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_192
timestamp 1649977179
transform 1 0 18768 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_199
timestamp 1649977179
transform 1 0 19412 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_211
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_228
timestamp 1649977179
transform 1 0 22080 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_239
timestamp 1649977179
transform 1 0 23092 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_248
timestamp 1649977179
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_252
timestamp 1649977179
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_255
timestamp 1649977179
transform 1 0 24564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_267
timestamp 1649977179
transform 1 0 25668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1649977179
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_300
timestamp 1649977179
transform 1 0 28704 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_312
timestamp 1649977179
transform 1 0 29808 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_321
timestamp 1649977179
transform 1 0 30636 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_333
timestamp 1649977179
transform 1 0 31740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_357
timestamp 1649977179
transform 1 0 33948 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_376
timestamp 1649977179
transform 1 0 35696 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_384
timestamp 1649977179
transform 1 0 36432 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1649977179
transform 1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_407
timestamp 1649977179
transform 1 0 38548 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_413
timestamp 1649977179
transform 1 0 39100 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_425
timestamp 1649977179
transform 1 0 40204 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_437
timestamp 1649977179
transform 1 0 41308 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1649977179
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1649977179
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1649977179
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1649977179
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1649977179
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_517
timestamp 1649977179
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_529
timestamp 1649977179
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_541
timestamp 1649977179
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_553
timestamp 1649977179
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_559
timestamp 1649977179
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp 1649977179
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_10
timestamp 1649977179
transform 1 0 2024 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1649977179
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_38
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_48
timestamp 1649977179
transform 1 0 5520 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_72
timestamp 1649977179
transform 1 0 7728 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_78
timestamp 1649977179
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_89
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_95
timestamp 1649977179
transform 1 0 9844 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_119
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_127
timestamp 1649977179
transform 1 0 12788 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp 1649977179
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_148
timestamp 1649977179
transform 1 0 14720 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_154
timestamp 1649977179
transform 1 0 15272 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_171
timestamp 1649977179
transform 1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_183
timestamp 1649977179
transform 1 0 17940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1649977179
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_199
timestamp 1649977179
transform 1 0 19412 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_205
timestamp 1649977179
transform 1 0 19964 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_211
timestamp 1649977179
transform 1 0 20516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_225
timestamp 1649977179
transform 1 0 21804 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_231
timestamp 1649977179
transform 1 0 22356 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1649977179
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_258
timestamp 1649977179
transform 1 0 24840 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_262
timestamp 1649977179
transform 1 0 25208 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_279
timestamp 1649977179
transform 1 0 26772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_291
timestamp 1649977179
transform 1 0 27876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_304
timestamp 1649977179
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_332
timestamp 1649977179
transform 1 0 31648 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_344
timestamp 1649977179
transform 1 0 32752 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_356
timestamp 1649977179
transform 1 0 33856 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_376
timestamp 1649977179
transform 1 0 35696 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_388
timestamp 1649977179
transform 1 0 36800 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_394
timestamp 1649977179
transform 1 0 37352 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_406
timestamp 1649977179
transform 1 0 38456 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_418
timestamp 1649977179
transform 1 0 39560 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1649977179
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1649977179
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1649977179
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1649977179
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1649977179
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1649977179
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1649977179
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_525
timestamp 1649977179
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_531
timestamp 1649977179
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_533
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_545
timestamp 1649977179
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_557
timestamp 1649977179
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_569
timestamp 1649977179
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_581
timestamp 1649977179
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1649977179
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_617
timestamp 1649977179
transform 1 0 57868 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_621
timestamp 1649977179
transform 1 0 58236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1649977179
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_33
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_41
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_65
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_78
timestamp 1649977179
transform 1 0 8280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1649977179
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_121
timestamp 1649977179
transform 1 0 12236 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_127
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_130
timestamp 1649977179
transform 1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_136
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_144
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_152
timestamp 1649977179
transform 1 0 15088 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_158
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_172
timestamp 1649977179
transform 1 0 16928 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_184
timestamp 1649977179
transform 1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_196
timestamp 1649977179
transform 1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_213
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_235
timestamp 1649977179
transform 1 0 22724 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_251
timestamp 1649977179
transform 1 0 24196 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_263
timestamp 1649977179
transform 1 0 25300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_275
timestamp 1649977179
transform 1 0 26404 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_290
timestamp 1649977179
transform 1 0 27784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_304
timestamp 1649977179
transform 1 0 29072 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_308
timestamp 1649977179
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_325
timestamp 1649977179
transform 1 0 31004 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_333
timestamp 1649977179
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_346
timestamp 1649977179
transform 1 0 32936 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_358
timestamp 1649977179
transform 1 0 34040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_363
timestamp 1649977179
transform 1 0 34500 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_375
timestamp 1649977179
transform 1 0 35604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_387
timestamp 1649977179
transform 1 0 36708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_402
timestamp 1649977179
transform 1 0 38088 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_414
timestamp 1649977179
transform 1 0 39192 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_426
timestamp 1649977179
transform 1 0 40296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_438
timestamp 1649977179
transform 1 0 41400 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp 1649977179
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1649977179
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1649977179
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1649977179
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1649977179
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1649977179
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_517
timestamp 1649977179
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_541
timestamp 1649977179
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_553
timestamp 1649977179
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_559
timestamp 1649977179
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1649977179
transform 1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_16
timestamp 1649977179
transform 1 0 2576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_20
timestamp 1649977179
transform 1 0 2944 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_23
timestamp 1649977179
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_40
timestamp 1649977179
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_54
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_60
timestamp 1649977179
transform 1 0 6624 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_64
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_70
timestamp 1649977179
transform 1 0 7544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_76
timestamp 1649977179
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_94
timestamp 1649977179
transform 1 0 9752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_100
timestamp 1649977179
transform 1 0 10304 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_108
timestamp 1649977179
transform 1 0 11040 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_118
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_126
timestamp 1649977179
transform 1 0 12696 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_134
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_171
timestamp 1649977179
transform 1 0 16836 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_175
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1649977179
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_213
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_220
timestamp 1649977179
transform 1 0 21344 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_236
timestamp 1649977179
transform 1 0 22816 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_240
timestamp 1649977179
transform 1 0 23184 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_243
timestamp 1649977179
transform 1 0 23460 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_295
timestamp 1649977179
transform 1 0 28244 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1649977179
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_344
timestamp 1649977179
transform 1 0 32752 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_355
timestamp 1649977179
transform 1 0 33764 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_381
timestamp 1649977179
transform 1 0 36156 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_396
timestamp 1649977179
transform 1 0 37536 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_416
timestamp 1649977179
transform 1 0 39376 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1649977179
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1649977179
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1649977179
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1649977179
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1649977179
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_533
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_545
timestamp 1649977179
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_557
timestamp 1649977179
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_569
timestamp 1649977179
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1649977179
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1649977179
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_617
timestamp 1649977179
transform 1 0 57868 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_621
timestamp 1649977179
transform 1 0 58236 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_9
timestamp 1649977179
transform 1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_29
timestamp 1649977179
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_45
timestamp 1649977179
transform 1 0 5244 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_59
timestamp 1649977179
transform 1 0 6532 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1649977179
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_70
timestamp 1649977179
transform 1 0 7544 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_74
timestamp 1649977179
transform 1 0 7912 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_80
timestamp 1649977179
transform 1 0 8464 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_100
timestamp 1649977179
transform 1 0 10304 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_106
timestamp 1649977179
transform 1 0 10856 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_121
timestamp 1649977179
transform 1 0 12236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_138
timestamp 1649977179
transform 1 0 13800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_155
timestamp 1649977179
transform 1 0 15364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_171
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1649977179
transform 1 0 17572 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_183
timestamp 1649977179
transform 1 0 17940 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_191
timestamp 1649977179
transform 1 0 18676 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_203
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_211
timestamp 1649977179
transform 1 0 20516 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1649977179
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_231
timestamp 1649977179
transform 1 0 22356 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_239
timestamp 1649977179
transform 1 0 23092 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_251
timestamp 1649977179
transform 1 0 24196 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_263
timestamp 1649977179
transform 1 0 25300 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_271
timestamp 1649977179
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_314
timestamp 1649977179
transform 1 0 29992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_320
timestamp 1649977179
transform 1 0 30544 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_328
timestamp 1649977179
transform 1 0 31280 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_332
timestamp 1649977179
transform 1 0 31648 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_345
timestamp 1649977179
transform 1 0 32844 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_357
timestamp 1649977179
transform 1 0 33948 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_369
timestamp 1649977179
transform 1 0 35052 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_376
timestamp 1649977179
transform 1 0 35696 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1649977179
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_401
timestamp 1649977179
transform 1 0 37996 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_421
timestamp 1649977179
transform 1 0 39836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_433
timestamp 1649977179
transform 1 0 40940 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_445
timestamp 1649977179
transform 1 0 42044 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1649977179
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1649977179
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1649977179
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1649977179
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1649977179
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_517
timestamp 1649977179
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_529
timestamp 1649977179
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_541
timestamp 1649977179
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_20
timestamp 1649977179
transform 1 0 2944 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_51
timestamp 1649977179
transform 1 0 5796 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_59
timestamp 1649977179
transform 1 0 6532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_71
timestamp 1649977179
transform 1 0 7636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_88
timestamp 1649977179
transform 1 0 9200 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_105
timestamp 1649977179
transform 1 0 10764 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_111
timestamp 1649977179
transform 1 0 11316 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_123
timestamp 1649977179
transform 1 0 12420 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1649977179
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_170
timestamp 1649977179
transform 1 0 16744 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_182
timestamp 1649977179
transform 1 0 17848 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_238
timestamp 1649977179
transform 1 0 23000 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1649977179
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_258
timestamp 1649977179
transform 1 0 24840 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_267
timestamp 1649977179
transform 1 0 25668 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_279
timestamp 1649977179
transform 1 0 26772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_287
timestamp 1649977179
transform 1 0 27508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_296
timestamp 1649977179
transform 1 0 28336 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1649977179
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_317
timestamp 1649977179
transform 1 0 30268 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_329
timestamp 1649977179
transform 1 0 31372 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_341
timestamp 1649977179
transform 1 0 32476 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_353
timestamp 1649977179
transform 1 0 33580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1649977179
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_387
timestamp 1649977179
transform 1 0 36708 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_411
timestamp 1649977179
transform 1 0 38916 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1649977179
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1649977179
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1649977179
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1649977179
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1649977179
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1649977179
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1649977179
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1649977179
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1649977179
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1649977179
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_525
timestamp 1649977179
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1649977179
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_533
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_545
timestamp 1649977179
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_557
timestamp 1649977179
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_569
timestamp 1649977179
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_581
timestamp 1649977179
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_45
timestamp 1649977179
transform 1 0 5244 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_65
timestamp 1649977179
transform 1 0 7084 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_77
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_89
timestamp 1649977179
transform 1 0 9292 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_95
timestamp 1649977179
transform 1 0 9844 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_107
timestamp 1649977179
transform 1 0 10948 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_121
timestamp 1649977179
transform 1 0 12236 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_133
timestamp 1649977179
transform 1 0 13340 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_145
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1649977179
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_177
timestamp 1649977179
transform 1 0 17388 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_189
timestamp 1649977179
transform 1 0 18492 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_196
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_208
timestamp 1649977179
transform 1 0 20240 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_212
timestamp 1649977179
transform 1 0 20608 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1649977179
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_234
timestamp 1649977179
transform 1 0 22632 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_241
timestamp 1649977179
transform 1 0 23276 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_245
timestamp 1649977179
transform 1 0 23644 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_256
timestamp 1649977179
transform 1 0 24656 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1649977179
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_285
timestamp 1649977179
transform 1 0 27324 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_288
timestamp 1649977179
transform 1 0 27600 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_295
timestamp 1649977179
transform 1 0 28244 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_319
timestamp 1649977179
transform 1 0 30452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_332
timestamp 1649977179
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_353
timestamp 1649977179
transform 1 0 33580 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_367
timestamp 1649977179
transform 1 0 34868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_387
timestamp 1649977179
transform 1 0 36708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_401
timestamp 1649977179
transform 1 0 37996 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_407
timestamp 1649977179
transform 1 0 38548 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_419
timestamp 1649977179
transform 1 0 39652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_431
timestamp 1649977179
transform 1 0 40756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_443
timestamp 1649977179
transform 1 0 41860 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1649977179
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1649977179
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1649977179
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1649977179
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1649977179
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_517
timestamp 1649977179
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_529
timestamp 1649977179
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_621
timestamp 1649977179
transform 1 0 58236 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_91
timestamp 1649977179
transform 1 0 9476 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_113
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_125
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_166
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_178
timestamp 1649977179
transform 1 0 17480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_199
timestamp 1649977179
transform 1 0 19412 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_16_210
timestamp 1649977179
transform 1 0 20424 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_214
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_239
timestamp 1649977179
transform 1 0 23092 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1649977179
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_274
timestamp 1649977179
transform 1 0 26312 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_286
timestamp 1649977179
transform 1 0 27416 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_294
timestamp 1649977179
transform 1 0 28152 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_299
timestamp 1649977179
transform 1 0 28612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_317
timestamp 1649977179
transform 1 0 30268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_322
timestamp 1649977179
transform 1 0 30728 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_342
timestamp 1649977179
transform 1 0 32568 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_354
timestamp 1649977179
transform 1 0 33672 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1649977179
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_368
timestamp 1649977179
transform 1 0 34960 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_380
timestamp 1649977179
transform 1 0 36064 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_395
timestamp 1649977179
transform 1 0 37444 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_398
timestamp 1649977179
transform 1 0 37720 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_404
timestamp 1649977179
transform 1 0 38272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_416
timestamp 1649977179
transform 1 0 39376 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1649977179
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1649977179
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1649977179
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1649977179
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1649977179
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1649977179
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_533
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_545
timestamp 1649977179
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_557
timestamp 1649977179
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_569
timestamp 1649977179
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_581
timestamp 1649977179
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_587
timestamp 1649977179
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_14
timestamp 1649977179
transform 1 0 2392 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_34
timestamp 1649977179
transform 1 0 4232 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_42
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 1649977179
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_64
timestamp 1649977179
transform 1 0 6992 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_96
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_157
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_163
timestamp 1649977179
transform 1 0 16100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_173
timestamp 1649977179
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_190
timestamp 1649977179
transform 1 0 18584 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_200
timestamp 1649977179
transform 1 0 19504 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_234
timestamp 1649977179
transform 1 0 22632 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_240
timestamp 1649977179
transform 1 0 23184 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_243
timestamp 1649977179
transform 1 0 23460 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_251
timestamp 1649977179
transform 1 0 24196 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_257
timestamp 1649977179
transform 1 0 24748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_269
timestamp 1649977179
transform 1 0 25852 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_277
timestamp 1649977179
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_297
timestamp 1649977179
transform 1 0 28428 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_309
timestamp 1649977179
transform 1 0 29532 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_320
timestamp 1649977179
transform 1 0 30544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1649977179
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_347
timestamp 1649977179
transform 1 0 33028 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_359
timestamp 1649977179
transform 1 0 34132 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_378
timestamp 1649977179
transform 1 0 35880 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_390
timestamp 1649977179
transform 1 0 36984 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_423
timestamp 1649977179
transform 1 0 40020 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_432
timestamp 1649977179
transform 1 0 40848 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_444
timestamp 1649977179
transform 1 0 41952 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1649977179
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1649977179
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1649977179
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1649977179
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_529
timestamp 1649977179
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_621
timestamp 1649977179
transform 1 0 58236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1649977179
transform 1 0 1748 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_11
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_20
timestamp 1649977179
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_66
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_94
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_100
timestamp 1649977179
transform 1 0 10304 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_108
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_143
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1649977179
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_159
timestamp 1649977179
transform 1 0 15732 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_180
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1649977179
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_206
timestamp 1649977179
transform 1 0 20056 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_217
timestamp 1649977179
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_229
timestamp 1649977179
transform 1 0 22172 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_235
timestamp 1649977179
transform 1 0 22724 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_247
timestamp 1649977179
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 1649977179
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_276
timestamp 1649977179
transform 1 0 26496 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_284
timestamp 1649977179
transform 1 0 27232 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_297
timestamp 1649977179
transform 1 0 28428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_305
timestamp 1649977179
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_313
timestamp 1649977179
transform 1 0 29900 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_316
timestamp 1649977179
transform 1 0 30176 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_328
timestamp 1649977179
transform 1 0 31280 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_340
timestamp 1649977179
transform 1 0 32384 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_346
timestamp 1649977179
transform 1 0 32936 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_354
timestamp 1649977179
transform 1 0 33672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_358
timestamp 1649977179
transform 1 0 34040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_375
timestamp 1649977179
transform 1 0 35604 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_381
timestamp 1649977179
transform 1 0 36156 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_393
timestamp 1649977179
transform 1 0 37260 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_397
timestamp 1649977179
transform 1 0 37628 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_408
timestamp 1649977179
transform 1 0 38640 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_431
timestamp 1649977179
transform 1 0 40756 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_443
timestamp 1649977179
transform 1 0 41860 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_455
timestamp 1649977179
transform 1 0 42964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_467
timestamp 1649977179
transform 1 0 44068 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1649977179
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1649977179
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1649977179
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1649977179
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_525
timestamp 1649977179
transform 1 0 49404 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_531
timestamp 1649977179
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 1649977179
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_18
timestamp 1649977179
transform 1 0 2760 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_24
timestamp 1649977179
transform 1 0 3312 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_35
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_41
timestamp 1649977179
transform 1 0 4876 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_66
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_72
timestamp 1649977179
transform 1 0 7728 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_99
timestamp 1649977179
transform 1 0 10212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_122
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_128
timestamp 1649977179
transform 1 0 12880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_140
timestamp 1649977179
transform 1 0 13984 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_146
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_155
timestamp 1649977179
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_188
timestamp 1649977179
transform 1 0 18400 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1649977179
transform 1 0 19504 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_208
timestamp 1649977179
transform 1 0 20240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_212
timestamp 1649977179
transform 1 0 20608 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_218
timestamp 1649977179
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_227
timestamp 1649977179
transform 1 0 21988 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_233
timestamp 1649977179
transform 1 0 22540 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_245
timestamp 1649977179
transform 1 0 23644 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_250
timestamp 1649977179
transform 1 0 24104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_274
timestamp 1649977179
transform 1 0 26312 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_283
timestamp 1649977179
transform 1 0 27140 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_295
timestamp 1649977179
transform 1 0 28244 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_312
timestamp 1649977179
transform 1 0 29808 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_322
timestamp 1649977179
transform 1 0 30728 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1649977179
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_339
timestamp 1649977179
transform 1 0 32292 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_351
timestamp 1649977179
transform 1 0 33396 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_357
timestamp 1649977179
transform 1 0 33948 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_368
timestamp 1649977179
transform 1 0 34960 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_372
timestamp 1649977179
transform 1 0 35328 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_381
timestamp 1649977179
transform 1 0 36156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1649977179
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_398
timestamp 1649977179
transform 1 0 37720 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_422
timestamp 1649977179
transform 1 0 39928 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_434
timestamp 1649977179
transform 1 0 41032 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_446
timestamp 1649977179
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1649977179
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1649977179
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1649977179
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1649977179
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1649977179
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_517
timestamp 1649977179
transform 1 0 48668 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_529
timestamp 1649977179
transform 1 0 49772 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_541
timestamp 1649977179
transform 1 0 50876 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_553
timestamp 1649977179
transform 1 0 51980 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_49
timestamp 1649977179
transform 1 0 5612 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_72
timestamp 1649977179
transform 1 0 7728 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_78
timestamp 1649977179
transform 1 0 8280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_151
timestamp 1649977179
transform 1 0 14996 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_163
timestamp 1649977179
transform 1 0 16100 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_175
timestamp 1649977179
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_184
timestamp 1649977179
transform 1 0 18032 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_192
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_200
timestamp 1649977179
transform 1 0 19504 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_208
timestamp 1649977179
transform 1 0 20240 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_216
timestamp 1649977179
transform 1 0 20976 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_219
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_227
timestamp 1649977179
transform 1 0 21988 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_231
timestamp 1649977179
transform 1 0 22356 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_237
timestamp 1649977179
transform 1 0 22908 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1649977179
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_261
timestamp 1649977179
transform 1 0 25116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_267
timestamp 1649977179
transform 1 0 25668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_275
timestamp 1649977179
transform 1 0 26404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_280
timestamp 1649977179
transform 1 0 26864 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_292
timestamp 1649977179
transform 1 0 27968 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_298
timestamp 1649977179
transform 1 0 28520 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1649977179
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_318
timestamp 1649977179
transform 1 0 30360 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_326
timestamp 1649977179
transform 1 0 31096 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_338
timestamp 1649977179
transform 1 0 32200 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1649977179
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_369
timestamp 1649977179
transform 1 0 35052 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_393
timestamp 1649977179
transform 1 0 37260 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_399
timestamp 1649977179
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_411
timestamp 1649977179
transform 1 0 38916 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1649977179
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_423
timestamp 1649977179
transform 1 0 40020 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_435
timestamp 1649977179
transform 1 0 41124 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_447
timestamp 1649977179
transform 1 0 42228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_459
timestamp 1649977179
transform 1 0 43332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_471
timestamp 1649977179
transform 1 0 44436 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_617
timestamp 1649977179
transform 1 0 57868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_621
timestamp 1649977179
transform 1 0 58236 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_19
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_23
timestamp 1649977179
transform 1 0 3220 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_35
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1649977179
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_65
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_68
timestamp 1649977179
transform 1 0 7360 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_74
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_86
timestamp 1649977179
transform 1 0 9016 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_98
timestamp 1649977179
transform 1 0 10120 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_147
timestamp 1649977179
transform 1 0 14628 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1649977179
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_192
timestamp 1649977179
transform 1 0 18768 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_196
timestamp 1649977179
transform 1 0 19136 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_199
timestamp 1649977179
transform 1 0 19412 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1649977179
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_229
timestamp 1649977179
transform 1 0 22172 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_240
timestamp 1649977179
transform 1 0 23184 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_244
timestamp 1649977179
transform 1 0 23552 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_251
timestamp 1649977179
transform 1 0 24196 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_267
timestamp 1649977179
transform 1 0 25668 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1649977179
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_297
timestamp 1649977179
transform 1 0 28428 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_325
timestamp 1649977179
transform 1 0 31004 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_333
timestamp 1649977179
transform 1 0 31740 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_355
timestamp 1649977179
transform 1 0 33764 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_358
timestamp 1649977179
transform 1 0 34040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_365
timestamp 1649977179
transform 1 0 34684 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_379
timestamp 1649977179
transform 1 0 35972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_388
timestamp 1649977179
transform 1 0 36800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_397
timestamp 1649977179
transform 1 0 37628 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_408
timestamp 1649977179
transform 1 0 38640 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_412
timestamp 1649977179
transform 1 0 39008 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1649977179
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1649977179
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1649977179
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1649977179
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1649977179
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1649977179
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1649977179
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1649977179
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1649977179
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1649977179
transform 1 0 5336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_52
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_56
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_73
timestamp 1649977179
transform 1 0 7820 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1649977179
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_102
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_108
timestamp 1649977179
transform 1 0 11040 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_116
timestamp 1649977179
transform 1 0 11776 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1649977179
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_170
timestamp 1649977179
transform 1 0 16744 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_176
timestamp 1649977179
transform 1 0 17296 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1649977179
transform 1 0 18400 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_202
timestamp 1649977179
transform 1 0 19688 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1649977179
transform 1 0 20424 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_217
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_232
timestamp 1649977179
transform 1 0 22448 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_243
timestamp 1649977179
transform 1 0 23460 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_259
timestamp 1649977179
transform 1 0 24932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_263
timestamp 1649977179
transform 1 0 25300 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_280
timestamp 1649977179
transform 1 0 26864 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_292
timestamp 1649977179
transform 1 0 27968 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_317
timestamp 1649977179
transform 1 0 30268 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_329
timestamp 1649977179
transform 1 0 31372 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_341
timestamp 1649977179
transform 1 0 32476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_356
timestamp 1649977179
transform 1 0 33856 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_375
timestamp 1649977179
transform 1 0 35604 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_384
timestamp 1649977179
transform 1 0 36432 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_412
timestamp 1649977179
transform 1 0 39008 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_426
timestamp 1649977179
transform 1 0 40296 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_434
timestamp 1649977179
transform 1 0 41032 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_446
timestamp 1649977179
transform 1 0 42136 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_458
timestamp 1649977179
transform 1 0 43240 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_470
timestamp 1649977179
transform 1 0 44344 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1649977179
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1649977179
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1649977179
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1649977179
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_525
timestamp 1649977179
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_531
timestamp 1649977179
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_617
timestamp 1649977179
transform 1 0 57868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_621
timestamp 1649977179
transform 1 0 58236 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_14
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_34
timestamp 1649977179
transform 1 0 4232 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1649977179
transform 1 0 4968 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1649977179
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_66
timestamp 1649977179
transform 1 0 7176 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_88
timestamp 1649977179
transform 1 0 9200 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_101
timestamp 1649977179
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_144
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_150
timestamp 1649977179
transform 1 0 14904 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_162
timestamp 1649977179
transform 1 0 16008 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_187
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_194
timestamp 1649977179
transform 1 0 18952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_200
timestamp 1649977179
transform 1 0 19504 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_206
timestamp 1649977179
transform 1 0 20056 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_229
timestamp 1649977179
transform 1 0 22172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_236
timestamp 1649977179
transform 1 0 22816 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_243
timestamp 1649977179
transform 1 0 23460 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_253
timestamp 1649977179
transform 1 0 24380 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_290
timestamp 1649977179
transform 1 0 27784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_296
timestamp 1649977179
transform 1 0 28336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_304
timestamp 1649977179
transform 1 0 29072 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_309
timestamp 1649977179
transform 1 0 29532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_321
timestamp 1649977179
transform 1 0 30636 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_345
timestamp 1649977179
transform 1 0 32844 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_350
timestamp 1649977179
transform 1 0 33304 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_362
timestamp 1649977179
transform 1 0 34408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_382
timestamp 1649977179
transform 1 0 36248 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1649977179
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_396
timestamp 1649977179
transform 1 0 37536 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_402
timestamp 1649977179
transform 1 0 38088 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_426
timestamp 1649977179
transform 1 0 40296 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_432
timestamp 1649977179
transform 1 0 40848 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_435
timestamp 1649977179
transform 1 0 41124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1649977179
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1649977179
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1649977179
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1649977179
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1649977179
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1649977179
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_16
timestamp 1649977179
transform 1 0 2576 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_64
timestamp 1649977179
transform 1 0 6992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_73
timestamp 1649977179
transform 1 0 7820 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1649977179
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_92
timestamp 1649977179
transform 1 0 9568 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_104
timestamp 1649977179
transform 1 0 10672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1649977179
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_144
timestamp 1649977179
transform 1 0 14352 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_168
timestamp 1649977179
transform 1 0 16560 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_180
timestamp 1649977179
transform 1 0 17664 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_186
timestamp 1649977179
transform 1 0 18216 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_213
timestamp 1649977179
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_220
timestamp 1649977179
transform 1 0 21344 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_228
timestamp 1649977179
transform 1 0 22080 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_235
timestamp 1649977179
transform 1 0 22724 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_242
timestamp 1649977179
transform 1 0 23368 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1649977179
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_255
timestamp 1649977179
transform 1 0 24564 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_267
timestamp 1649977179
transform 1 0 25668 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_279
timestamp 1649977179
transform 1 0 26772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_284
timestamp 1649977179
transform 1 0 27232 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_290
timestamp 1649977179
transform 1 0 27784 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_302
timestamp 1649977179
transform 1 0 28888 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_325
timestamp 1649977179
transform 1 0 31004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_337
timestamp 1649977179
transform 1 0 32108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_343
timestamp 1649977179
transform 1 0 32660 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_349
timestamp 1649977179
transform 1 0 33212 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1649977179
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_383
timestamp 1649977179
transform 1 0 36340 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_387
timestamp 1649977179
transform 1 0 36708 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_390
timestamp 1649977179
transform 1 0 36984 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_399
timestamp 1649977179
transform 1 0 37812 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_411
timestamp 1649977179
transform 1 0 38916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1649977179
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_431
timestamp 1649977179
transform 1 0 40756 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_443
timestamp 1649977179
transform 1 0 41860 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_455
timestamp 1649977179
transform 1 0 42964 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_467
timestamp 1649977179
transform 1 0 44068 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1649977179
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_9
timestamp 1649977179
transform 1 0 1932 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_26
timestamp 1649977179
transform 1 0 3496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1649977179
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_63
timestamp 1649977179
transform 1 0 6900 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_66
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_78
timestamp 1649977179
transform 1 0 8280 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_90
timestamp 1649977179
transform 1 0 9384 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_94
timestamp 1649977179
transform 1 0 9752 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_101
timestamp 1649977179
transform 1 0 10396 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_121
timestamp 1649977179
transform 1 0 12236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_128
timestamp 1649977179
transform 1 0 12880 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_136
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_139
timestamp 1649977179
transform 1 0 13892 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_153
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1649977179
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_174
timestamp 1649977179
transform 1 0 17112 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_183
timestamp 1649977179
transform 1 0 17940 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_200
timestamp 1649977179
transform 1 0 19504 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_209
timestamp 1649977179
transform 1 0 20332 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_216
timestamp 1649977179
transform 1 0 20976 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_229
timestamp 1649977179
transform 1 0 22172 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_232
timestamp 1649977179
transform 1 0 22448 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_248
timestamp 1649977179
transform 1 0 23920 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_260
timestamp 1649977179
transform 1 0 25024 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_272
timestamp 1649977179
transform 1 0 26128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_276
timestamp 1649977179
transform 1 0 26496 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_288
timestamp 1649977179
transform 1 0 27600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_300
timestamp 1649977179
transform 1 0 28704 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_309
timestamp 1649977179
transform 1 0 29532 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_323
timestamp 1649977179
transform 1 0 30820 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_330
timestamp 1649977179
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_369
timestamp 1649977179
transform 1 0 35052 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_380
timestamp 1649977179
transform 1 0 36064 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_400
timestamp 1649977179
transform 1 0 37904 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_406
timestamp 1649977179
transform 1 0 38456 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_426
timestamp 1649977179
transform 1 0 40296 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_438
timestamp 1649977179
transform 1 0 41400 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_446
timestamp 1649977179
transform 1 0 42136 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1649977179
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1649977179
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1649977179
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1649977179
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_621
timestamp 1649977179
transform 1 0 58236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_11
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_37
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_46
timestamp 1649977179
transform 1 0 5336 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_58
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_66
timestamp 1649977179
transform 1 0 7176 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_76
timestamp 1649977179
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_87
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_95
timestamp 1649977179
transform 1 0 9844 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_98
timestamp 1649977179
transform 1 0 10120 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_104
timestamp 1649977179
transform 1 0 10672 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_110
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_122
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1649977179
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_131
timestamp 1649977179
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_149
timestamp 1649977179
transform 1 0 14812 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_152
timestamp 1649977179
transform 1 0 15088 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1649977179
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_176
timestamp 1649977179
transform 1 0 17296 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1649977179
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_201
timestamp 1649977179
transform 1 0 19596 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_207
timestamp 1649977179
transform 1 0 20148 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_213
timestamp 1649977179
transform 1 0 20700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_219
timestamp 1649977179
transform 1 0 21252 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_229
timestamp 1649977179
transform 1 0 22172 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1649977179
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_285
timestamp 1649977179
transform 1 0 27324 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_297
timestamp 1649977179
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1649977179
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_326
timestamp 1649977179
transform 1 0 31096 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_340
timestamp 1649977179
transform 1 0 32384 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_352
timestamp 1649977179
transform 1 0 33488 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_395
timestamp 1649977179
transform 1 0 37444 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_407
timestamp 1649977179
transform 1 0 38548 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1649977179
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_421
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_429
timestamp 1649977179
transform 1 0 40572 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_441
timestamp 1649977179
transform 1 0 41676 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_453
timestamp 1649977179
transform 1 0 42780 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_465
timestamp 1649977179
transform 1 0 43884 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_473
timestamp 1649977179
transform 1 0 44620 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1649977179
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1649977179
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1649977179
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1649977179
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1649977179
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_34
timestamp 1649977179
transform 1 0 4232 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_38
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1649977179
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1649977179
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_83
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_95
timestamp 1649977179
transform 1 0 9844 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1649977179
transform 1 0 10948 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_122
timestamp 1649977179
transform 1 0 12328 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_134
timestamp 1649977179
transform 1 0 13432 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_146
timestamp 1649977179
transform 1 0 14536 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_160
timestamp 1649977179
transform 1 0 15824 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_171
timestamp 1649977179
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_175
timestamp 1649977179
transform 1 0 17204 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_178
timestamp 1649977179
transform 1 0 17480 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_184
timestamp 1649977179
transform 1 0 18032 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_194
timestamp 1649977179
transform 1 0 18952 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_200
timestamp 1649977179
transform 1 0 19504 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_207
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_215
timestamp 1649977179
transform 1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1649977179
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_239
timestamp 1649977179
transform 1 0 23092 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_253
timestamp 1649977179
transform 1 0 24380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_263
timestamp 1649977179
transform 1 0 25300 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_274
timestamp 1649977179
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_286
timestamp 1649977179
transform 1 0 27416 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_292
timestamp 1649977179
transform 1 0 27968 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_304
timestamp 1649977179
transform 1 0 29072 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_316
timestamp 1649977179
transform 1 0 30176 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1649977179
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_381
timestamp 1649977179
transform 1 0 36156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1649977179
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_398
timestamp 1649977179
transform 1 0 37720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_406
timestamp 1649977179
transform 1 0 38456 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_418
timestamp 1649977179
transform 1 0 39560 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_430
timestamp 1649977179
transform 1 0 40664 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_442
timestamp 1649977179
transform 1 0 41768 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1649977179
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1649977179
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1649977179
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1649977179
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1649977179
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1649977179
transform 1 0 58236 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_33
timestamp 1649977179
transform 1 0 4140 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_36
timestamp 1649977179
transform 1 0 4416 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_48
timestamp 1649977179
transform 1 0 5520 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_54
timestamp 1649977179
transform 1 0 6072 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_66
timestamp 1649977179
transform 1 0 7176 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_76
timestamp 1649977179
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_88
timestamp 1649977179
transform 1 0 9200 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_100
timestamp 1649977179
transform 1 0 10304 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_104
timestamp 1649977179
transform 1 0 10672 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_107
timestamp 1649977179
transform 1 0 10948 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_113
timestamp 1649977179
transform 1 0 11500 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_125
timestamp 1649977179
transform 1 0 12604 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_157
timestamp 1649977179
transform 1 0 15548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_169
timestamp 1649977179
transform 1 0 16652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_181
timestamp 1649977179
transform 1 0 17756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_193
timestamp 1649977179
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_205
timestamp 1649977179
transform 1 0 19964 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_241
timestamp 1649977179
transform 1 0 23276 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_249
timestamp 1649977179
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_260
timestamp 1649977179
transform 1 0 25024 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_266
timestamp 1649977179
transform 1 0 25576 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_275
timestamp 1649977179
transform 1 0 26404 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_281
timestamp 1649977179
transform 1 0 26956 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_293
timestamp 1649977179
transform 1 0 28060 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1649977179
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_317
timestamp 1649977179
transform 1 0 30268 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_323
timestamp 1649977179
transform 1 0 30820 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_337
timestamp 1649977179
transform 1 0 32108 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_349
timestamp 1649977179
transform 1 0 33212 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1649977179
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_371
timestamp 1649977179
transform 1 0 35236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_383
timestamp 1649977179
transform 1 0 36340 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_394
timestamp 1649977179
transform 1 0 37352 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_402
timestamp 1649977179
transform 1 0 38088 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_414
timestamp 1649977179
transform 1 0 39192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_421
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_428
timestamp 1649977179
transform 1 0 40480 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_434
timestamp 1649977179
transform 1 0 41032 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_446
timestamp 1649977179
transform 1 0 42136 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_458
timestamp 1649977179
transform 1 0 43240 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_470
timestamp 1649977179
transform 1 0 44344 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_589
timestamp 1649977179
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_601
timestamp 1649977179
transform 1 0 56396 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_613
timestamp 1649977179
transform 1 0 57500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_9
timestamp 1649977179
transform 1 0 1932 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_24
timestamp 1649977179
transform 1 0 3312 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_31
timestamp 1649977179
transform 1 0 3956 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_35
timestamp 1649977179
transform 1 0 4324 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_38
timestamp 1649977179
transform 1 0 4600 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_46
timestamp 1649977179
transform 1 0 5336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_52
timestamp 1649977179
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_59
timestamp 1649977179
transform 1 0 6532 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_72
timestamp 1649977179
transform 1 0 7728 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_80
timestamp 1649977179
transform 1 0 8464 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_121
timestamp 1649977179
transform 1 0 12236 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_127
timestamp 1649977179
transform 1 0 12788 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_130
timestamp 1649977179
transform 1 0 13064 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_142
timestamp 1649977179
transform 1 0 14168 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_154
timestamp 1649977179
transform 1 0 15272 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_173
timestamp 1649977179
transform 1 0 17020 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1649977179
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_185
timestamp 1649977179
transform 1 0 18124 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_189
timestamp 1649977179
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_195
timestamp 1649977179
transform 1 0 19044 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_201
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_204
timestamp 1649977179
transform 1 0 19872 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_211
timestamp 1649977179
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1649977179
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_257
timestamp 1649977179
transform 1 0 24748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_274
timestamp 1649977179
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_309
timestamp 1649977179
transform 1 0 29532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_316
timestamp 1649977179
transform 1 0 30176 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1649977179
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_343
timestamp 1649977179
transform 1 0 32660 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_352
timestamp 1649977179
transform 1 0 33488 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_381
timestamp 1649977179
transform 1 0 36156 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_403
timestamp 1649977179
transform 1 0 38180 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_425
timestamp 1649977179
transform 1 0 40204 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_437
timestamp 1649977179
transform 1 0 41308 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_443
timestamp 1649977179
transform 1 0 41860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1649977179
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1649977179
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1649977179
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1649977179
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1649977179
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_24
timestamp 1649977179
transform 1 0 3312 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_38
timestamp 1649977179
transform 1 0 4600 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_50
timestamp 1649977179
transform 1 0 5704 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_58
timestamp 1649977179
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1649977179
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_115
timestamp 1649977179
transform 1 0 11684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_124
timestamp 1649977179
transform 1 0 12512 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_130
timestamp 1649977179
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_147
timestamp 1649977179
transform 1 0 14628 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_161
timestamp 1649977179
transform 1 0 15916 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_173
timestamp 1649977179
transform 1 0 17020 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_179
timestamp 1649977179
transform 1 0 17572 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_188
timestamp 1649977179
transform 1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_213
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_227
timestamp 1649977179
transform 1 0 21988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_235
timestamp 1649977179
transform 1 0 22724 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1649977179
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_255
timestamp 1649977179
transform 1 0 24564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_261
timestamp 1649977179
transform 1 0 25116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_269
timestamp 1649977179
transform 1 0 25852 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_275
timestamp 1649977179
transform 1 0 26404 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_278
timestamp 1649977179
transform 1 0 26680 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_286
timestamp 1649977179
transform 1 0 27416 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_298
timestamp 1649977179
transform 1 0 28520 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1649977179
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_316
timestamp 1649977179
transform 1 0 30176 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_326
timestamp 1649977179
transform 1 0 31096 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_332
timestamp 1649977179
transform 1 0 31648 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_335
timestamp 1649977179
transform 1 0 31924 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_347
timestamp 1649977179
transform 1 0 33028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_359
timestamp 1649977179
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_387
timestamp 1649977179
transform 1 0 36708 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_399
timestamp 1649977179
transform 1 0 37812 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_411
timestamp 1649977179
transform 1 0 38916 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1649977179
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_423
timestamp 1649977179
transform 1 0 40020 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_435
timestamp 1649977179
transform 1 0 41124 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_444
timestamp 1649977179
transform 1 0 41952 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_456
timestamp 1649977179
transform 1 0 43056 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_468
timestamp 1649977179
transform 1 0 44160 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1649977179
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1649977179
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1649977179
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1649977179
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1649977179
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_617
timestamp 1649977179
transform 1 0 57868 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_621
timestamp 1649977179
transform 1 0 58236 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_36
timestamp 1649977179
transform 1 0 4416 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_49
timestamp 1649977179
transform 1 0 5612 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_67
timestamp 1649977179
transform 1 0 7268 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_78
timestamp 1649977179
transform 1 0 8280 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_87
timestamp 1649977179
transform 1 0 9108 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_118
timestamp 1649977179
transform 1 0 11960 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_126
timestamp 1649977179
transform 1 0 12696 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_138
timestamp 1649977179
transform 1 0 13800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_145
timestamp 1649977179
transform 1 0 14444 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_154
timestamp 1649977179
transform 1 0 15272 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1649977179
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_185
timestamp 1649977179
transform 1 0 18124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_197
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_230
timestamp 1649977179
transform 1 0 22264 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_242
timestamp 1649977179
transform 1 0 23368 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_254
timestamp 1649977179
transform 1 0 24472 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1649977179
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_287
timestamp 1649977179
transform 1 0 27508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_304
timestamp 1649977179
transform 1 0 29072 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_318
timestamp 1649977179
transform 1 0 30360 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_359
timestamp 1649977179
transform 1 0 34132 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_371
timestamp 1649977179
transform 1 0 35236 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_386
timestamp 1649977179
transform 1 0 36616 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_398
timestamp 1649977179
transform 1 0 37720 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_422
timestamp 1649977179
transform 1 0 39928 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_442
timestamp 1649977179
transform 1 0 41768 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1649977179
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1649977179
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1649977179
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1649977179
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1649977179
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_17
timestamp 1649977179
transform 1 0 2668 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1649977179
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_39
timestamp 1649977179
transform 1 0 4692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_47
timestamp 1649977179
transform 1 0 5428 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_50
timestamp 1649977179
transform 1 0 5704 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_56
timestamp 1649977179
transform 1 0 6256 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_62
timestamp 1649977179
transform 1 0 6808 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_72
timestamp 1649977179
transform 1 0 7728 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1649977179
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_89
timestamp 1649977179
transform 1 0 9292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_106
timestamp 1649977179
transform 1 0 10856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_118
timestamp 1649977179
transform 1 0 11960 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_134
timestamp 1649977179
transform 1 0 13432 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_32_151
timestamp 1649977179
transform 1 0 14996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_162
timestamp 1649977179
transform 1 0 16008 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_174
timestamp 1649977179
transform 1 0 17112 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_186
timestamp 1649977179
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_201
timestamp 1649977179
transform 1 0 19596 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_210
timestamp 1649977179
transform 1 0 20424 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_222
timestamp 1649977179
transform 1 0 21528 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_227
timestamp 1649977179
transform 1 0 21988 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_287
timestamp 1649977179
transform 1 0 27508 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_293
timestamp 1649977179
transform 1 0 28060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1649977179
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_320
timestamp 1649977179
transform 1 0 30544 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_332
timestamp 1649977179
transform 1 0 31648 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_340
timestamp 1649977179
transform 1 0 32384 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_348
timestamp 1649977179
transform 1 0 33120 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1649977179
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_381
timestamp 1649977179
transform 1 0 36156 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_392
timestamp 1649977179
transform 1 0 37168 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_403
timestamp 1649977179
transform 1 0 38180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_411
timestamp 1649977179
transform 1 0 38916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_416
timestamp 1649977179
transform 1 0 39376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1649977179
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1649977179
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_457
timestamp 1649977179
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1649977179
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1649977179
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1649977179
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1649977179
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1649977179
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_525
timestamp 1649977179
transform 1 0 49404 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_617
timestamp 1649977179
transform 1 0 57868 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1649977179
transform 1 0 58236 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_63
timestamp 1649977179
transform 1 0 6900 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_73
timestamp 1649977179
transform 1 0 7820 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_79
timestamp 1649977179
transform 1 0 8372 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_91
timestamp 1649977179
transform 1 0 9476 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_103
timestamp 1649977179
transform 1 0 10580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_117
timestamp 1649977179
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_120
timestamp 1649977179
transform 1 0 12144 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_124
timestamp 1649977179
transform 1 0 12512 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_157
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1649977179
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_175
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_184
timestamp 1649977179
transform 1 0 18032 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_192
timestamp 1649977179
transform 1 0 18768 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_202
timestamp 1649977179
transform 1 0 19688 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_214
timestamp 1649977179
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1649977179
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_229
timestamp 1649977179
transform 1 0 22172 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_235
timestamp 1649977179
transform 1 0 22724 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_255
timestamp 1649977179
transform 1 0 24564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_267
timestamp 1649977179
transform 1 0 25668 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_274
timestamp 1649977179
transform 1 0 26312 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_289
timestamp 1649977179
transform 1 0 27692 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_295
timestamp 1649977179
transform 1 0 28244 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_298
timestamp 1649977179
transform 1 0 28520 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_304
timestamp 1649977179
transform 1 0 29072 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_312
timestamp 1649977179
transform 1 0 29808 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_322
timestamp 1649977179
transform 1 0 30728 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_334
timestamp 1649977179
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_348
timestamp 1649977179
transform 1 0 33120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_368
timestamp 1649977179
transform 1 0 34960 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_376
timestamp 1649977179
transform 1 0 35696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1649977179
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_400
timestamp 1649977179
transform 1 0 37904 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_420
timestamp 1649977179
transform 1 0 39744 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1649977179
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1649977179
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1649977179
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1649977179
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1649977179
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1649977179
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1649977179
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1649977179
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_58
timestamp 1649977179
transform 1 0 6440 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_62
timestamp 1649977179
transform 1 0 6808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_73
timestamp 1649977179
transform 1 0 7820 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1649977179
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_93
timestamp 1649977179
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1649977179
transform 1 0 9936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_106
timestamp 1649977179
transform 1 0 10856 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_118
timestamp 1649977179
transform 1 0 11960 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_124
timestamp 1649977179
transform 1 0 12512 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_128
timestamp 1649977179
transform 1 0 12880 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_134
timestamp 1649977179
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_149
timestamp 1649977179
transform 1 0 14812 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_175
timestamp 1649977179
transform 1 0 17204 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_184
timestamp 1649977179
transform 1 0 18032 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_205
timestamp 1649977179
transform 1 0 19964 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_212
timestamp 1649977179
transform 1 0 20608 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_224
timestamp 1649977179
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_231
timestamp 1649977179
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_243
timestamp 1649977179
transform 1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_258
timestamp 1649977179
transform 1 0 24840 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_278
timestamp 1649977179
transform 1 0 26680 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_286
timestamp 1649977179
transform 1 0 27416 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1649977179
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_298
timestamp 1649977179
transform 1 0 28520 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1649977179
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_317
timestamp 1649977179
transform 1 0 30268 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_329
timestamp 1649977179
transform 1 0 31372 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_337
timestamp 1649977179
transform 1 0 32108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_340
timestamp 1649977179
transform 1 0 32384 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_352
timestamp 1649977179
transform 1 0 33488 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1649977179
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1649977179
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1649977179
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1649977179
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1649977179
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1649977179
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_501
timestamp 1649977179
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_513
timestamp 1649977179
transform 1 0 48300 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_525
timestamp 1649977179
transform 1 0 49404 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_9
timestamp 1649977179
transform 1 0 1932 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_18
timestamp 1649977179
transform 1 0 2760 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_24
timestamp 1649977179
transform 1 0 3312 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_36
timestamp 1649977179
transform 1 0 4416 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_42
timestamp 1649977179
transform 1 0 4968 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1649977179
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_73
timestamp 1649977179
transform 1 0 7820 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_79
timestamp 1649977179
transform 1 0 8372 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_91
timestamp 1649977179
transform 1 0 9476 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_102
timestamp 1649977179
transform 1 0 10488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1649977179
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_145
timestamp 1649977179
transform 1 0 14444 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_153
timestamp 1649977179
transform 1 0 15180 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_163
timestamp 1649977179
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_185
timestamp 1649977179
transform 1 0 18124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_197
timestamp 1649977179
transform 1 0 19228 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_209
timestamp 1649977179
transform 1 0 20332 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_212
timestamp 1649977179
transform 1 0 20608 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1649977179
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_245
timestamp 1649977179
transform 1 0 23644 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_257
timestamp 1649977179
transform 1 0 24748 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_269
timestamp 1649977179
transform 1 0 25852 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_277
timestamp 1649977179
transform 1 0 26588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_284
timestamp 1649977179
transform 1 0 27232 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_296
timestamp 1649977179
transform 1 0 28336 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_300
timestamp 1649977179
transform 1 0 28704 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_315
timestamp 1649977179
transform 1 0 30084 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1649977179
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_343
timestamp 1649977179
transform 1 0 32660 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_350
timestamp 1649977179
transform 1 0 33304 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_362
timestamp 1649977179
transform 1 0 34408 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_374
timestamp 1649977179
transform 1 0 35512 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_380
timestamp 1649977179
transform 1 0 36064 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_423
timestamp 1649977179
transform 1 0 40020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_435
timestamp 1649977179
transform 1 0 41124 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1649977179
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_473
timestamp 1649977179
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_485
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1649977179
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1649977179
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_621
timestamp 1649977179
transform 1 0 58236 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_7
timestamp 1649977179
transform 1 0 1748 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1649977179
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_45
timestamp 1649977179
transform 1 0 5244 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_63
timestamp 1649977179
transform 1 0 6900 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_75
timestamp 1649977179
transform 1 0 8004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_87
timestamp 1649977179
transform 1 0 9108 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_36_102
timestamp 1649977179
transform 1 0 10488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_110
timestamp 1649977179
transform 1 0 11224 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_115
timestamp 1649977179
transform 1 0 11684 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_123
timestamp 1649977179
transform 1 0 12420 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_135
timestamp 1649977179
transform 1 0 13524 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_149
timestamp 1649977179
transform 1 0 14812 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_152
timestamp 1649977179
transform 1 0 15088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_156
timestamp 1649977179
transform 1 0 15456 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1649977179
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_168
timestamp 1649977179
transform 1 0 16560 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_180
timestamp 1649977179
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1649977179
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_202
timestamp 1649977179
transform 1 0 19688 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_210
timestamp 1649977179
transform 1 0 20424 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_234
timestamp 1649977179
transform 1 0 22632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_246
timestamp 1649977179
transform 1 0 23736 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_255
timestamp 1649977179
transform 1 0 24564 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_267
timestamp 1649977179
transform 1 0 25668 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_279
timestamp 1649977179
transform 1 0 26772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_282
timestamp 1649977179
transform 1 0 27048 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1649977179
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_342
timestamp 1649977179
transform 1 0 32568 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_352
timestamp 1649977179
transform 1 0 33488 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_384
timestamp 1649977179
transform 1 0 36432 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_396
timestamp 1649977179
transform 1 0 37536 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_408
timestamp 1649977179
transform 1 0 38640 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1649977179
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_429
timestamp 1649977179
transform 1 0 40572 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_441
timestamp 1649977179
transform 1 0 41676 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_453
timestamp 1649977179
transform 1 0 42780 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_465
timestamp 1649977179
transform 1 0 43884 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_473
timestamp 1649977179
transform 1 0 44620 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_10
timestamp 1649977179
transform 1 0 2024 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_30
timestamp 1649977179
transform 1 0 3864 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1649977179
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_76
timestamp 1649977179
transform 1 0 8096 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_83
timestamp 1649977179
transform 1 0 8740 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_95
timestamp 1649977179
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_101
timestamp 1649977179
transform 1 0 10396 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_109
timestamp 1649977179
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_120
timestamp 1649977179
transform 1 0 12144 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_132
timestamp 1649977179
transform 1 0 13248 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_140
timestamp 1649977179
transform 1 0 13984 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_148
timestamp 1649977179
transform 1 0 14720 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_158
timestamp 1649977179
transform 1 0 15640 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1649977179
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_179
timestamp 1649977179
transform 1 0 17572 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_185
timestamp 1649977179
transform 1 0 18124 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_207
timestamp 1649977179
transform 1 0 20148 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1649977179
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_37_230
timestamp 1649977179
transform 1 0 22264 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_238
timestamp 1649977179
transform 1 0 23000 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_246
timestamp 1649977179
transform 1 0 23736 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_257
timestamp 1649977179
transform 1 0 24748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_264
timestamp 1649977179
transform 1 0 25392 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1649977179
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_289
timestamp 1649977179
transform 1 0 27692 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_296
timestamp 1649977179
transform 1 0 28336 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_308
timestamp 1649977179
transform 1 0 29440 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_320
timestamp 1649977179
transform 1 0 30544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_324
timestamp 1649977179
transform 1 0 30912 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1649977179
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_341
timestamp 1649977179
transform 1 0 32476 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_350
timestamp 1649977179
transform 1 0 33304 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_376
timestamp 1649977179
transform 1 0 35696 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1649977179
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_398
timestamp 1649977179
transform 1 0 37720 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_410
timestamp 1649977179
transform 1 0 38824 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_416
timestamp 1649977179
transform 1 0 39376 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_422
timestamp 1649977179
transform 1 0 39928 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_434
timestamp 1649977179
transform 1 0 41032 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_446
timestamp 1649977179
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1649977179
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1649977179
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1649977179
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_621
timestamp 1649977179
transform 1 0 58236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_11
timestamp 1649977179
transform 1 0 2116 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1649977179
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_31
timestamp 1649977179
transform 1 0 3956 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_43
timestamp 1649977179
transform 1 0 5060 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_55
timestamp 1649977179
transform 1 0 6164 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_71
timestamp 1649977179
transform 1 0 7636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_105
timestamp 1649977179
transform 1 0 10764 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_123
timestamp 1649977179
transform 1 0 12420 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_132
timestamp 1649977179
transform 1 0 13248 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_143
timestamp 1649977179
transform 1 0 14260 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_156
timestamp 1649977179
transform 1 0 15456 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_162
timestamp 1649977179
transform 1 0 16008 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_172
timestamp 1649977179
transform 1 0 16928 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_184
timestamp 1649977179
transform 1 0 18032 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_202
timestamp 1649977179
transform 1 0 19688 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_214
timestamp 1649977179
transform 1 0 20792 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_224
timestamp 1649977179
transform 1 0 21712 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_234
timestamp 1649977179
transform 1 0 22632 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1649977179
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_261
timestamp 1649977179
transform 1 0 25116 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_282
timestamp 1649977179
transform 1 0 27048 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_294
timestamp 1649977179
transform 1 0 28152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_306
timestamp 1649977179
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_311
timestamp 1649977179
transform 1 0 29716 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_323
timestamp 1649977179
transform 1 0 30820 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_331
timestamp 1649977179
transform 1 0 31556 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_339
timestamp 1649977179
transform 1 0 32292 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_359
timestamp 1649977179
transform 1 0 34132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_371
timestamp 1649977179
transform 1 0 35236 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_374
timestamp 1649977179
transform 1 0 35512 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_394
timestamp 1649977179
transform 1 0 37352 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_406
timestamp 1649977179
transform 1 0 38456 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_416
timestamp 1649977179
transform 1 0 39376 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_421
timestamp 1649977179
transform 1 0 39836 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_430
timestamp 1649977179
transform 1 0 40664 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_436
timestamp 1649977179
transform 1 0 41216 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_448
timestamp 1649977179
transform 1 0 42320 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_460
timestamp 1649977179
transform 1 0 43424 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_472
timestamp 1649977179
transform 1 0 44528 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1649977179
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_501
timestamp 1649977179
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_513
timestamp 1649977179
transform 1 0 48300 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_525
timestamp 1649977179
transform 1 0 49404 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_531
timestamp 1649977179
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_11
timestamp 1649977179
transform 1 0 2116 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_17
timestamp 1649977179
transform 1 0 2668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_29
timestamp 1649977179
transform 1 0 3772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_41
timestamp 1649977179
transform 1 0 4876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_53
timestamp 1649977179
transform 1 0 5980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1649977179
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_72
timestamp 1649977179
transform 1 0 7728 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_94
timestamp 1649977179
transform 1 0 9752 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_103
timestamp 1649977179
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_121
timestamp 1649977179
transform 1 0 12236 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_143
timestamp 1649977179
transform 1 0 14260 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_187
timestamp 1649977179
transform 1 0 18308 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_199
timestamp 1649977179
transform 1 0 19412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_211
timestamp 1649977179
transform 1 0 20516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_239
timestamp 1649977179
transform 1 0 23092 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_251
timestamp 1649977179
transform 1 0 24196 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1649977179
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_260
timestamp 1649977179
transform 1 0 25024 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 1649977179
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_297
timestamp 1649977179
transform 1 0 28428 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_314
timestamp 1649977179
transform 1 0 29992 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_326
timestamp 1649977179
transform 1 0 31096 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1649977179
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_342
timestamp 1649977179
transform 1 0 32568 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_348
timestamp 1649977179
transform 1 0 33120 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_355
timestamp 1649977179
transform 1 0 33764 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_367
timestamp 1649977179
transform 1 0 34868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_375
timestamp 1649977179
transform 1 0 35604 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_384
timestamp 1649977179
transform 1 0 36432 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_425
timestamp 1649977179
transform 1 0 40204 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_437
timestamp 1649977179
transform 1 0 41308 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_445
timestamp 1649977179
transform 1 0 42044 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1649977179
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1649977179
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1649977179
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_505
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_517
timestamp 1649977179
transform 1 0 48668 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_529
timestamp 1649977179
transform 1 0 49772 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_541
timestamp 1649977179
transform 1 0 50876 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_553
timestamp 1649977179
transform 1 0 51980 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1649977179
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_71
timestamp 1649977179
transform 1 0 7636 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_74
timestamp 1649977179
transform 1 0 7912 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1649977179
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_101
timestamp 1649977179
transform 1 0 10396 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_107
timestamp 1649977179
transform 1 0 10948 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_110
timestamp 1649977179
transform 1 0 11224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_122
timestamp 1649977179
transform 1 0 12328 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_134
timestamp 1649977179
transform 1 0 13432 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_152
timestamp 1649977179
transform 1 0 15088 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_158
timestamp 1649977179
transform 1 0 15640 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_166
timestamp 1649977179
transform 1 0 16376 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_169
timestamp 1649977179
transform 1 0 16652 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_202
timestamp 1649977179
transform 1 0 19688 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_222
timestamp 1649977179
transform 1 0 21528 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_234
timestamp 1649977179
transform 1 0 22632 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1649977179
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_260
timestamp 1649977179
transform 1 0 25024 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_280
timestamp 1649977179
transform 1 0 26864 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_288
timestamp 1649977179
transform 1 0 27600 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_295
timestamp 1649977179
transform 1 0 28244 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1649977179
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_317
timestamp 1649977179
transform 1 0 30268 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_323
timestamp 1649977179
transform 1 0 30820 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_335
timestamp 1649977179
transform 1 0 31924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_347
timestamp 1649977179
transform 1 0 33028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_359
timestamp 1649977179
transform 1 0 34132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1649977179
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1649977179
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_428
timestamp 1649977179
transform 1 0 40480 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_437
timestamp 1649977179
transform 1 0 41308 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_449
timestamp 1649977179
transform 1 0 42412 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_461
timestamp 1649977179
transform 1 0 43516 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_473
timestamp 1649977179
transform 1 0 44620 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1649977179
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_617
timestamp 1649977179
transform 1 0 57868 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1649977179
transform 1 0 58236 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_31
timestamp 1649977179
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_43
timestamp 1649977179
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_59
timestamp 1649977179
transform 1 0 6532 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_71
timestamp 1649977179
transform 1 0 7636 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_83
timestamp 1649977179
transform 1 0 8740 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_89
timestamp 1649977179
transform 1 0 9292 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_101
timestamp 1649977179
transform 1 0 10396 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_107
timestamp 1649977179
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_117
timestamp 1649977179
transform 1 0 11868 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_120
timestamp 1649977179
transform 1 0 12144 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_126
timestamp 1649977179
transform 1 0 12696 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_132
timestamp 1649977179
transform 1 0 13248 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_138
timestamp 1649977179
transform 1 0 13800 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_144
timestamp 1649977179
transform 1 0 14352 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_173
timestamp 1649977179
transform 1 0 17020 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_189
timestamp 1649977179
transform 1 0 18492 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_209
timestamp 1649977179
transform 1 0 20332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_221
timestamp 1649977179
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_239
timestamp 1649977179
transform 1 0 23092 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_251
timestamp 1649977179
transform 1 0 24196 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_254
timestamp 1649977179
transform 1 0 24472 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_266
timestamp 1649977179
transform 1 0 25576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1649977179
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_297
timestamp 1649977179
transform 1 0 28428 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1649977179
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_339
timestamp 1649977179
transform 1 0 32292 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_353
timestamp 1649977179
transform 1 0 33580 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_377
timestamp 1649977179
transform 1 0 35788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1649977179
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_398
timestamp 1649977179
transform 1 0 37720 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_406
timestamp 1649977179
transform 1 0 38456 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_424
timestamp 1649977179
transform 1 0 40112 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_436
timestamp 1649977179
transform 1 0 41216 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1649977179
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1649977179
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1649977179
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1649977179
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_73
timestamp 1649977179
transform 1 0 7820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1649977179
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_96
timestamp 1649977179
transform 1 0 9936 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_120
timestamp 1649977179
transform 1 0 12144 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_126
timestamp 1649977179
transform 1 0 12696 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1649977179
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_143
timestamp 1649977179
transform 1 0 14260 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_149
timestamp 1649977179
transform 1 0 14812 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_155
timestamp 1649977179
transform 1 0 15364 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_173
timestamp 1649977179
transform 1 0 17020 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_180
timestamp 1649977179
transform 1 0 17664 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1649977179
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_199
timestamp 1649977179
transform 1 0 19412 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_211
timestamp 1649977179
transform 1 0 20516 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_239
timestamp 1649977179
transform 1 0 23092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_271
timestamp 1649977179
transform 1 0 26036 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_283
timestamp 1649977179
transform 1 0 27140 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_295
timestamp 1649977179
transform 1 0 28244 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1649977179
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_317
timestamp 1649977179
transform 1 0 30268 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_323
timestamp 1649977179
transform 1 0 30820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_327
timestamp 1649977179
transform 1 0 31188 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_344
timestamp 1649977179
transform 1 0 32752 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_356
timestamp 1649977179
transform 1 0 33856 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_373
timestamp 1649977179
transform 1 0 35420 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_392
timestamp 1649977179
transform 1 0 37168 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_404
timestamp 1649977179
transform 1 0 38272 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_410
timestamp 1649977179
transform 1 0 38824 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1649977179
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_429
timestamp 1649977179
transform 1 0 40572 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_435
timestamp 1649977179
transform 1 0 41124 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_447
timestamp 1649977179
transform 1 0 42228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_459
timestamp 1649977179
transform 1 0 43332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_471
timestamp 1649977179
transform 1 0 44436 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_617
timestamp 1649977179
transform 1 0 57868 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_621
timestamp 1649977179
transform 1 0 58236 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_32
timestamp 1649977179
transform 1 0 4048 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_44
timestamp 1649977179
transform 1 0 5152 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_65
timestamp 1649977179
transform 1 0 7084 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_71
timestamp 1649977179
transform 1 0 7636 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_77
timestamp 1649977179
transform 1 0 8188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_87
timestamp 1649977179
transform 1 0 9108 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_43_95
timestamp 1649977179
transform 1 0 9844 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_101
timestamp 1649977179
transform 1 0 10396 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_106
timestamp 1649977179
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_130
timestamp 1649977179
transform 1 0 13064 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_138
timestamp 1649977179
transform 1 0 13800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_146
timestamp 1649977179
transform 1 0 14536 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_160
timestamp 1649977179
transform 1 0 15824 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_172
timestamp 1649977179
transform 1 0 16928 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_188
timestamp 1649977179
transform 1 0 18400 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_197
timestamp 1649977179
transform 1 0 19228 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_206
timestamp 1649977179
transform 1 0 20056 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_214
timestamp 1649977179
transform 1 0 20792 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1649977179
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_233
timestamp 1649977179
transform 1 0 22540 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_239
timestamp 1649977179
transform 1 0 23092 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_251
timestamp 1649977179
transform 1 0 24196 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_259
timestamp 1649977179
transform 1 0 24932 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_264
timestamp 1649977179
transform 1 0 25392 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_283
timestamp 1649977179
transform 1 0 27140 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_309
timestamp 1649977179
transform 1 0 29532 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_318
timestamp 1649977179
transform 1 0 30360 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_330
timestamp 1649977179
transform 1 0 31464 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_345
timestamp 1649977179
transform 1 0 32844 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_362
timestamp 1649977179
transform 1 0 34408 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_374
timestamp 1649977179
transform 1 0 35512 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_386
timestamp 1649977179
transform 1 0 36616 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_396
timestamp 1649977179
transform 1 0 37536 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_404
timestamp 1649977179
transform 1 0 38272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_423
timestamp 1649977179
transform 1 0 40020 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_435
timestamp 1649977179
transform 1 0 41124 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1649977179
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_9
timestamp 1649977179
transform 1 0 1932 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_12
timestamp 1649977179
transform 1 0 2208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1649977179
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_34
timestamp 1649977179
transform 1 0 4232 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_40
timestamp 1649977179
transform 1 0 4784 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_52
timestamp 1649977179
transform 1 0 5888 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_58
timestamp 1649977179
transform 1 0 6440 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_70
timestamp 1649977179
transform 1 0 7544 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_74
timestamp 1649977179
transform 1 0 7912 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_89
timestamp 1649977179
transform 1 0 9292 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_93
timestamp 1649977179
transform 1 0 9660 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_101
timestamp 1649977179
transform 1 0 10396 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_106
timestamp 1649977179
transform 1 0 10856 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_114
timestamp 1649977179
transform 1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_118
timestamp 1649977179
transform 1 0 11960 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_129
timestamp 1649977179
transform 1 0 12972 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_135
timestamp 1649977179
transform 1 0 13524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_167
timestamp 1649977179
transform 1 0 16468 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_176
timestamp 1649977179
transform 1 0 17296 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1649977179
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_199
timestamp 1649977179
transform 1 0 19412 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_211
timestamp 1649977179
transform 1 0 20516 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_215
timestamp 1649977179
transform 1 0 20884 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_264
timestamp 1649977179
transform 1 0 25392 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_276
timestamp 1649977179
transform 1 0 26496 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_285
timestamp 1649977179
transform 1 0 27324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_297
timestamp 1649977179
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1649977179
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_311
timestamp 1649977179
transform 1 0 29716 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_317
timestamp 1649977179
transform 1 0 30268 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_329
timestamp 1649977179
transform 1 0 31372 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_337
timestamp 1649977179
transform 1 0 32108 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_340
timestamp 1649977179
transform 1 0 32384 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_351
timestamp 1649977179
transform 1 0 33396 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_381
timestamp 1649977179
transform 1 0 36156 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_393
timestamp 1649977179
transform 1 0 37260 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_399
timestamp 1649977179
transform 1 0 37812 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1649977179
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_426
timestamp 1649977179
transform 1 0 40296 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_432
timestamp 1649977179
transform 1 0 40848 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_444
timestamp 1649977179
transform 1 0 41952 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_456
timestamp 1649977179
transform 1 0 43056 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_468
timestamp 1649977179
transform 1 0 44160 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1649977179
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1649977179
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_501
timestamp 1649977179
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_513
timestamp 1649977179
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1649977179
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1649977179
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_24
timestamp 1649977179
transform 1 0 3312 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_33
timestamp 1649977179
transform 1 0 4140 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_49
timestamp 1649977179
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_73
timestamp 1649977179
transform 1 0 7820 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_85
timestamp 1649977179
transform 1 0 8924 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_89
timestamp 1649977179
transform 1 0 9292 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_94
timestamp 1649977179
transform 1 0 9752 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1649977179
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_124
timestamp 1649977179
transform 1 0 12512 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_138
timestamp 1649977179
transform 1 0 13800 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_150
timestamp 1649977179
transform 1 0 14904 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1649977179
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_173
timestamp 1649977179
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_190
timestamp 1649977179
transform 1 0 18584 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_210
timestamp 1649977179
transform 1 0 20424 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1649977179
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_230
timestamp 1649977179
transform 1 0 22264 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_250
timestamp 1649977179
transform 1 0 24104 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_258
timestamp 1649977179
transform 1 0 24840 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1649977179
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_289
timestamp 1649977179
transform 1 0 27692 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_307
timestamp 1649977179
transform 1 0 29348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_315
timestamp 1649977179
transform 1 0 30084 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_323
timestamp 1649977179
transform 1 0 30820 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_326
timestamp 1649977179
transform 1 0 31096 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1649977179
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_348
timestamp 1649977179
transform 1 0 33120 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_364
timestamp 1649977179
transform 1 0 34592 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_409
timestamp 1649977179
transform 1 0 38732 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_433
timestamp 1649977179
transform 1 0 40940 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_445
timestamp 1649977179
transform 1 0 42044 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1649977179
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1649977179
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1649977179
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1649977179
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_621
timestamp 1649977179
transform 1 0 58236 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_21
timestamp 1649977179
transform 1 0 3036 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1649977179
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_31
timestamp 1649977179
transform 1 0 3956 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_39
timestamp 1649977179
transform 1 0 4692 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_50
timestamp 1649977179
transform 1 0 5704 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_62
timestamp 1649977179
transform 1 0 6808 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_73
timestamp 1649977179
transform 1 0 7820 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_81
timestamp 1649977179
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_87
timestamp 1649977179
transform 1 0 9108 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_96
timestamp 1649977179
transform 1 0 9936 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_108
timestamp 1649977179
transform 1 0 11040 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_116
timestamp 1649977179
transform 1 0 11776 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_136
timestamp 1649977179
transform 1 0 13616 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_147
timestamp 1649977179
transform 1 0 14628 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_150
timestamp 1649977179
transform 1 0 14904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_158
timestamp 1649977179
transform 1 0 15640 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_166
timestamp 1649977179
transform 1 0 16376 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_170
timestamp 1649977179
transform 1 0 16744 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_178
timestamp 1649977179
transform 1 0 17480 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1649977179
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1649977179
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_205
timestamp 1649977179
transform 1 0 19964 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_210
timestamp 1649977179
transform 1 0 20424 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_234
timestamp 1649977179
transform 1 0 22632 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_246
timestamp 1649977179
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_256
timestamp 1649977179
transform 1 0 24656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_268
timestamp 1649977179
transform 1 0 25760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_292
timestamp 1649977179
transform 1 0 27968 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_300
timestamp 1649977179
transform 1 0 28704 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1649977179
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_322
timestamp 1649977179
transform 1 0 30728 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_336
timestamp 1649977179
transform 1 0 32016 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_347
timestamp 1649977179
transform 1 0 33028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_356
timestamp 1649977179
transform 1 0 33856 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_381
timestamp 1649977179
transform 1 0 36156 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_393
timestamp 1649977179
transform 1 0 37260 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_405
timestamp 1649977179
transform 1 0 38364 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_417
timestamp 1649977179
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_421
timestamp 1649977179
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_445
timestamp 1649977179
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_457
timestamp 1649977179
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1649977179
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1649977179
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1649977179
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_489
timestamp 1649977179
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_501
timestamp 1649977179
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_513
timestamp 1649977179
transform 1 0 48300 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1649977179
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_31
timestamp 1649977179
transform 1 0 3956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_43
timestamp 1649977179
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_68
timestamp 1649977179
transform 1 0 7360 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_74
timestamp 1649977179
transform 1 0 7912 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_90
timestamp 1649977179
transform 1 0 9384 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1649977179
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_118
timestamp 1649977179
transform 1 0 11960 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_124
timestamp 1649977179
transform 1 0 12512 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_132
timestamp 1649977179
transform 1 0 13248 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_143
timestamp 1649977179
transform 1 0 14260 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_147
timestamp 1649977179
transform 1 0 14628 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1649977179
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_172
timestamp 1649977179
transform 1 0 16928 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_194
timestamp 1649977179
transform 1 0 18952 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_198
timestamp 1649977179
transform 1 0 19320 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_209
timestamp 1649977179
transform 1 0 20332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_221
timestamp 1649977179
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_233
timestamp 1649977179
transform 1 0 22540 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_241
timestamp 1649977179
transform 1 0 23276 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_246
timestamp 1649977179
transform 1 0 23736 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_254
timestamp 1649977179
transform 1 0 24472 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_260
timestamp 1649977179
transform 1 0 25024 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_272
timestamp 1649977179
transform 1 0 26128 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_310
timestamp 1649977179
transform 1 0 29624 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_317
timestamp 1649977179
transform 1 0 30268 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_321
timestamp 1649977179
transform 1 0 30636 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1649977179
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_339
timestamp 1649977179
transform 1 0 32292 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_351
timestamp 1649977179
transform 1 0 33396 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_364
timestamp 1649977179
transform 1 0 34592 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_376
timestamp 1649977179
transform 1 0 35696 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1649977179
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_417
timestamp 1649977179
transform 1 0 39468 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1649977179
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1649977179
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1649977179
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1649977179
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1649977179
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1649977179
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_621
timestamp 1649977179
transform 1 0 58236 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_21
timestamp 1649977179
transform 1 0 3036 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_31
timestamp 1649977179
transform 1 0 3956 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_43
timestamp 1649977179
transform 1 0 5060 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_55
timestamp 1649977179
transform 1 0 6164 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_67
timestamp 1649977179
transform 1 0 7268 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_71
timestamp 1649977179
transform 1 0 7636 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1649977179
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_94
timestamp 1649977179
transform 1 0 9752 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_100
timestamp 1649977179
transform 1 0 10304 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_106
timestamp 1649977179
transform 1 0 10856 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_118
timestamp 1649977179
transform 1 0 11960 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_122
timestamp 1649977179
transform 1 0 12328 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_130
timestamp 1649977179
transform 1 0 13064 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_136
timestamp 1649977179
transform 1 0 13616 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_146
timestamp 1649977179
transform 1 0 14536 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_158
timestamp 1649977179
transform 1 0 15640 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_162
timestamp 1649977179
transform 1 0 16008 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_167
timestamp 1649977179
transform 1 0 16468 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_179
timestamp 1649977179
transform 1 0 17572 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_191
timestamp 1649977179
transform 1 0 18676 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_201
timestamp 1649977179
transform 1 0 19596 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_204
timestamp 1649977179
transform 1 0 19872 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_212
timestamp 1649977179
transform 1 0 20608 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_218
timestamp 1649977179
transform 1 0 21160 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_226
timestamp 1649977179
transform 1 0 21896 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_238
timestamp 1649977179
transform 1 0 23000 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1649977179
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_260
timestamp 1649977179
transform 1 0 25024 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_266
timestamp 1649977179
transform 1 0 25576 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_276
timestamp 1649977179
transform 1 0 26496 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_284
timestamp 1649977179
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1649977179
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_311
timestamp 1649977179
transform 1 0 29716 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_325
timestamp 1649977179
transform 1 0 31004 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_331
timestamp 1649977179
transform 1 0 31556 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_343
timestamp 1649977179
transform 1 0 32660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_356
timestamp 1649977179
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_372
timestamp 1649977179
transform 1 0 35328 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_380
timestamp 1649977179
transform 1 0 36064 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_393
timestamp 1649977179
transform 1 0 37260 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_410
timestamp 1649977179
transform 1 0 38824 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_418
timestamp 1649977179
transform 1 0 39560 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_457
timestamp 1649977179
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1649977179
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1649977179
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1649977179
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1649977179
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_513
timestamp 1649977179
transform 1 0 48300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_525
timestamp 1649977179
transform 1 0 49404 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_531
timestamp 1649977179
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_26
timestamp 1649977179
transform 1 0 3496 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_41
timestamp 1649977179
transform 1 0 4876 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_52
timestamp 1649977179
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_89
timestamp 1649977179
transform 1 0 9292 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_96
timestamp 1649977179
transform 1 0 9936 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1649977179
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_139
timestamp 1649977179
transform 1 0 13892 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_143
timestamp 1649977179
transform 1 0 14260 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_146
timestamp 1649977179
transform 1 0 14536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_155
timestamp 1649977179
transform 1 0 15364 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_163
timestamp 1649977179
transform 1 0 16100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_187
timestamp 1649977179
transform 1 0 18308 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_204
timestamp 1649977179
transform 1 0 19872 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_212
timestamp 1649977179
transform 1 0 20608 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1649977179
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_231
timestamp 1649977179
transform 1 0 22356 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_236
timestamp 1649977179
transform 1 0 22816 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_248
timestamp 1649977179
transform 1 0 23920 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_254
timestamp 1649977179
transform 1 0 24472 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_262
timestamp 1649977179
transform 1 0 25208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_270
timestamp 1649977179
transform 1 0 25944 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1649977179
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_295
timestamp 1649977179
transform 1 0 28244 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_319
timestamp 1649977179
transform 1 0 30452 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_328
timestamp 1649977179
transform 1 0 31280 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_345
timestamp 1649977179
transform 1 0 32844 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_356
timestamp 1649977179
transform 1 0 33856 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_368
timestamp 1649977179
transform 1 0 34960 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_376
timestamp 1649977179
transform 1 0 35696 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1649977179
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_423
timestamp 1649977179
transform 1 0 40020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_435
timestamp 1649977179
transform 1 0 41124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1649977179
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1649977179
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1649977179
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1649977179
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1649977179
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_40
timestamp 1649977179
transform 1 0 4784 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_52
timestamp 1649977179
transform 1 0 5888 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_64
timestamp 1649977179
transform 1 0 6992 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_67
timestamp 1649977179
transform 1 0 7268 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_79
timestamp 1649977179
transform 1 0 8372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_92
timestamp 1649977179
transform 1 0 9568 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_98
timestamp 1649977179
transform 1 0 10120 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_102
timestamp 1649977179
transform 1 0 10488 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_119
timestamp 1649977179
transform 1 0 12052 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_131
timestamp 1649977179
transform 1 0 13156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_143
timestamp 1649977179
transform 1 0 14260 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_151
timestamp 1649977179
transform 1 0 14996 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_157
timestamp 1649977179
transform 1 0 15548 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_169
timestamp 1649977179
transform 1 0 16652 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_174
timestamp 1649977179
transform 1 0 17112 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_180
timestamp 1649977179
transform 1 0 17664 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1649977179
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_200
timestamp 1649977179
transform 1 0 19504 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_208
timestamp 1649977179
transform 1 0 20240 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_216
timestamp 1649977179
transform 1 0 20976 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_224
timestamp 1649977179
transform 1 0 21712 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_228
timestamp 1649977179
transform 1 0 22080 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_236
timestamp 1649977179
transform 1 0 22816 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_244
timestamp 1649977179
transform 1 0 23552 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1649977179
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_264
timestamp 1649977179
transform 1 0 25392 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_284
timestamp 1649977179
transform 1 0 27232 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_296
timestamp 1649977179
transform 1 0 28336 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1649977179
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_316
timestamp 1649977179
transform 1 0 30176 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_323
timestamp 1649977179
transform 1 0 30820 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_329
timestamp 1649977179
transform 1 0 31372 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_341
timestamp 1649977179
transform 1 0 32476 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1649977179
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_368
timestamp 1649977179
transform 1 0 34960 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_382
timestamp 1649977179
transform 1 0 36248 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_388
timestamp 1649977179
transform 1 0 36800 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_416
timestamp 1649977179
transform 1 0 39376 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_433
timestamp 1649977179
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_445
timestamp 1649977179
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_457
timestamp 1649977179
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1649977179
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1649977179
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_617
timestamp 1649977179
transform 1 0 57868 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_621
timestamp 1649977179
transform 1 0 58236 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_11
timestamp 1649977179
transform 1 0 2116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_30
timestamp 1649977179
transform 1 0 3864 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_73
timestamp 1649977179
transform 1 0 7820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_85
timestamp 1649977179
transform 1 0 8924 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_97
timestamp 1649977179
transform 1 0 10028 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_103
timestamp 1649977179
transform 1 0 10580 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_121
timestamp 1649977179
transform 1 0 12236 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_127
timestamp 1649977179
transform 1 0 12788 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_139
timestamp 1649977179
transform 1 0 13892 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_151
timestamp 1649977179
transform 1 0 14996 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_160
timestamp 1649977179
transform 1 0 15824 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_173
timestamp 1649977179
transform 1 0 17020 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_176
timestamp 1649977179
transform 1 0 17296 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_196
timestamp 1649977179
transform 1 0 19136 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_208
timestamp 1649977179
transform 1 0 20240 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_236
timestamp 1649977179
transform 1 0 22816 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_248
timestamp 1649977179
transform 1 0 23920 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_256
timestamp 1649977179
transform 1 0 24656 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_260
timestamp 1649977179
transform 1 0 25024 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_265
timestamp 1649977179
transform 1 0 25484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_283
timestamp 1649977179
transform 1 0 27140 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_313
timestamp 1649977179
transform 1 0 29900 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_326
timestamp 1649977179
transform 1 0 31096 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1649977179
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_343
timestamp 1649977179
transform 1 0 32660 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_357
timestamp 1649977179
transform 1 0 33948 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_368
timestamp 1649977179
transform 1 0 34960 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_374
timestamp 1649977179
transform 1 0 35512 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_386
timestamp 1649977179
transform 1 0 36616 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_398
timestamp 1649977179
transform 1 0 37720 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_410
timestamp 1649977179
transform 1 0 38824 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_422
timestamp 1649977179
transform 1 0 39928 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_434
timestamp 1649977179
transform 1 0 41032 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_446
timestamp 1649977179
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1649977179
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1649977179
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1649977179
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1649977179
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1649977179
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1649977179
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_11
timestamp 1649977179
transform 1 0 2116 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_19
timestamp 1649977179
transform 1 0 2852 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_47
timestamp 1649977179
transform 1 0 5428 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_73
timestamp 1649977179
transform 1 0 7820 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_78
timestamp 1649977179
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_87
timestamp 1649977179
transform 1 0 9108 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_99
timestamp 1649977179
transform 1 0 10212 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1649977179
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_143
timestamp 1649977179
transform 1 0 14260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_174
timestamp 1649977179
transform 1 0 17112 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_180
timestamp 1649977179
transform 1 0 17664 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_183
timestamp 1649977179
transform 1 0 17940 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1649977179
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_201
timestamp 1649977179
transform 1 0 19596 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_204
timestamp 1649977179
transform 1 0 19872 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_218
timestamp 1649977179
transform 1 0 21160 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_240
timestamp 1649977179
transform 1 0 23184 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_246
timestamp 1649977179
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_255
timestamp 1649977179
transform 1 0 24564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_267
timestamp 1649977179
transform 1 0 25668 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_271
timestamp 1649977179
transform 1 0 26036 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_288
timestamp 1649977179
transform 1 0 27600 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_300
timestamp 1649977179
transform 1 0 28704 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_312
timestamp 1649977179
transform 1 0 29808 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_323
timestamp 1649977179
transform 1 0 30820 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_335
timestamp 1649977179
transform 1 0 31924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_355
timestamp 1649977179
transform 1 0 33764 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_374
timestamp 1649977179
transform 1 0 35512 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_386
timestamp 1649977179
transform 1 0 36616 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_392
timestamp 1649977179
transform 1 0 37168 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_416
timestamp 1649977179
transform 1 0 39376 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_445
timestamp 1649977179
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_457
timestamp 1649977179
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1649977179
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1649977179
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_617
timestamp 1649977179
transform 1 0 57868 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_621
timestamp 1649977179
transform 1 0 58236 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_11
timestamp 1649977179
transform 1 0 2116 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_19
timestamp 1649977179
transform 1 0 2852 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_31
timestamp 1649977179
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_45
timestamp 1649977179
transform 1 0 5244 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1649977179
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_61
timestamp 1649977179
transform 1 0 6716 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_73
timestamp 1649977179
transform 1 0 7820 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_83
timestamp 1649977179
transform 1 0 8740 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_89
timestamp 1649977179
transform 1 0 9292 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_101
timestamp 1649977179
transform 1 0 10396 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1649977179
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_118
timestamp 1649977179
transform 1 0 11960 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_124
timestamp 1649977179
transform 1 0 12512 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_136
timestamp 1649977179
transform 1 0 13616 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_142
timestamp 1649977179
transform 1 0 14168 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_148
timestamp 1649977179
transform 1 0 14720 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_157
timestamp 1649977179
transform 1 0 15548 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1649977179
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1649977179
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1649977179
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_235
timestamp 1649977179
transform 1 0 22724 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_243
timestamp 1649977179
transform 1 0 23460 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_247
timestamp 1649977179
transform 1 0 23828 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_250
timestamp 1649977179
transform 1 0 24104 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_258
timestamp 1649977179
transform 1 0 24840 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_310
timestamp 1649977179
transform 1 0 29624 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_319
timestamp 1649977179
transform 1 0 30452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_330
timestamp 1649977179
transform 1 0 31464 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_340
timestamp 1649977179
transform 1 0 32384 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_352
timestamp 1649977179
transform 1 0 33488 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_364
timestamp 1649977179
transform 1 0 34592 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_376
timestamp 1649977179
transform 1 0 35696 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_382
timestamp 1649977179
transform 1 0 36248 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1649977179
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_417
timestamp 1649977179
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_429
timestamp 1649977179
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1649977179
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1649977179
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_449
timestamp 1649977179
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_461
timestamp 1649977179
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_473
timestamp 1649977179
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_485
timestamp 1649977179
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1649977179
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1649977179
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_9
timestamp 1649977179
transform 1 0 1932 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_18
timestamp 1649977179
transform 1 0 2760 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1649977179
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_49
timestamp 1649977179
transform 1 0 5612 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_70
timestamp 1649977179
transform 1 0 7544 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_79
timestamp 1649977179
transform 1 0 8372 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_105
timestamp 1649977179
transform 1 0 10764 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_111
timestamp 1649977179
transform 1 0 11316 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_128
timestamp 1649977179
transform 1 0 12880 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_143
timestamp 1649977179
transform 1 0 14260 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_155
timestamp 1649977179
transform 1 0 15364 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_167
timestamp 1649977179
transform 1 0 16468 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_171
timestamp 1649977179
transform 1 0 16836 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_174
timestamp 1649977179
transform 1 0 17112 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_188
timestamp 1649977179
transform 1 0 18400 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_224
timestamp 1649977179
transform 1 0 21712 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_237
timestamp 1649977179
transform 1 0 22908 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1649977179
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_263
timestamp 1649977179
transform 1 0 25300 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_275
timestamp 1649977179
transform 1 0 26404 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_287
timestamp 1649977179
transform 1 0 27508 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_299
timestamp 1649977179
transform 1 0 28612 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_303
timestamp 1649977179
transform 1 0 28980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_327
timestamp 1649977179
transform 1 0 31188 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_339
timestamp 1649977179
transform 1 0 32292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_351
timestamp 1649977179
transform 1 0 33396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_373
timestamp 1649977179
transform 1 0 35420 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_376
timestamp 1649977179
transform 1 0 35696 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_388
timestamp 1649977179
transform 1 0 36800 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_412
timestamp 1649977179
transform 1 0 39008 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_433
timestamp 1649977179
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_445
timestamp 1649977179
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_457
timestamp 1649977179
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1649977179
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1649977179
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_11
timestamp 1649977179
transform 1 0 2116 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_28
timestamp 1649977179
transform 1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_40
timestamp 1649977179
transform 1 0 4784 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1649977179
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_73
timestamp 1649977179
transform 1 0 7820 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_79
timestamp 1649977179
transform 1 0 8372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_95
timestamp 1649977179
transform 1 0 9844 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_104
timestamp 1649977179
transform 1 0 10672 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_121
timestamp 1649977179
transform 1 0 12236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_129
timestamp 1649977179
transform 1 0 12972 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_146
timestamp 1649977179
transform 1 0 14536 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_155
timestamp 1649977179
transform 1 0 15364 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_159
timestamp 1649977179
transform 1 0 15732 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1649977179
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_173
timestamp 1649977179
transform 1 0 17020 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_194
timestamp 1649977179
transform 1 0 18952 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_214
timestamp 1649977179
transform 1 0 20792 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1649977179
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_235
timestamp 1649977179
transform 1 0 22724 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_246
timestamp 1649977179
transform 1 0 23736 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_266
timestamp 1649977179
transform 1 0 25576 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_278
timestamp 1649977179
transform 1 0 26680 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_303
timestamp 1649977179
transform 1 0 28980 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_315
timestamp 1649977179
transform 1 0 30084 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_321
timestamp 1649977179
transform 1 0 30636 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 1649977179
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_342
timestamp 1649977179
transform 1 0 32568 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_354
timestamp 1649977179
transform 1 0 33672 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_364
timestamp 1649977179
transform 1 0 34592 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_388
timestamp 1649977179
transform 1 0 36800 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_417
timestamp 1649977179
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_429
timestamp 1649977179
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1649977179
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1649977179
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_621
timestamp 1649977179
transform 1 0 58236 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_31
timestamp 1649977179
transform 1 0 3956 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_43
timestamp 1649977179
transform 1 0 5060 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_55
timestamp 1649977179
transform 1 0 6164 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_58
timestamp 1649977179
transform 1 0 6440 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_70
timestamp 1649977179
transform 1 0 7544 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_79
timestamp 1649977179
transform 1 0 8372 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_157
timestamp 1649977179
transform 1 0 15548 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_163
timestamp 1649977179
transform 1 0 16100 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_172
timestamp 1649977179
transform 1 0 16928 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_184
timestamp 1649977179
transform 1 0 18032 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1649977179
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_199
timestamp 1649977179
transform 1 0 19412 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_205
timestamp 1649977179
transform 1 0 19964 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_217
timestamp 1649977179
transform 1 0 21068 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_229
timestamp 1649977179
transform 1 0 22172 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_241
timestamp 1649977179
transform 1 0 23276 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1649977179
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_316
timestamp 1649977179
transform 1 0 30176 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_324
timestamp 1649977179
transform 1 0 30912 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_328
timestamp 1649977179
transform 1 0 31280 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_331
timestamp 1649977179
transform 1 0 31556 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_343
timestamp 1649977179
transform 1 0 32660 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_351
timestamp 1649977179
transform 1 0 33396 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1649977179
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_383
timestamp 1649977179
transform 1 0 36340 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_395
timestamp 1649977179
transform 1 0 37444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_407
timestamp 1649977179
transform 1 0 38548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_31
timestamp 1649977179
transform 1 0 3956 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_40
timestamp 1649977179
transform 1 0 4784 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1649977179
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_61
timestamp 1649977179
transform 1 0 6716 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_78
timestamp 1649977179
transform 1 0 8280 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_90
timestamp 1649977179
transform 1 0 9384 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_102
timestamp 1649977179
transform 1 0 10488 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_110
timestamp 1649977179
transform 1 0 11224 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_130
timestamp 1649977179
transform 1 0 13064 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_142
timestamp 1649977179
transform 1 0 14168 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_156
timestamp 1649977179
transform 1 0 15456 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_174
timestamp 1649977179
transform 1 0 17112 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_180
timestamp 1649977179
transform 1 0 17664 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_184
timestamp 1649977179
transform 1 0 18032 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_190
timestamp 1649977179
transform 1 0 18584 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_198
timestamp 1649977179
transform 1 0 19320 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_204
timestamp 1649977179
transform 1 0 19872 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_216
timestamp 1649977179
transform 1 0 20976 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_243
timestamp 1649977179
transform 1 0 23460 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_267
timestamp 1649977179
transform 1 0 25668 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_285
timestamp 1649977179
transform 1 0 27324 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_297
timestamp 1649977179
transform 1 0 28428 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_306
timestamp 1649977179
transform 1 0 29256 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_310
timestamp 1649977179
transform 1 0 29624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_313
timestamp 1649977179
transform 1 0 29900 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_325
timestamp 1649977179
transform 1 0 31004 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_333
timestamp 1649977179
transform 1 0 31740 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_350
timestamp 1649977179
transform 1 0 33304 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_364
timestamp 1649977179
transform 1 0 34592 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_384
timestamp 1649977179
transform 1 0 36432 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_417
timestamp 1649977179
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_429
timestamp 1649977179
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1649977179
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_621
timestamp 1649977179
transform 1 0 58236 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_9
timestamp 1649977179
transform 1 0 1932 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_12
timestamp 1649977179
transform 1 0 2208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1649977179
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_37
timestamp 1649977179
transform 1 0 4508 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_43
timestamp 1649977179
transform 1 0 5060 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_49
timestamp 1649977179
transform 1 0 5612 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_61
timestamp 1649977179
transform 1 0 6716 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_73
timestamp 1649977179
transform 1 0 7820 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_81
timestamp 1649977179
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_93
timestamp 1649977179
transform 1 0 9660 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_101
timestamp 1649977179
transform 1 0 10396 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_108
timestamp 1649977179
transform 1 0 11040 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_114
timestamp 1649977179
transform 1 0 11592 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_120
timestamp 1649977179
transform 1 0 12144 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_132
timestamp 1649977179
transform 1 0 13248 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_145
timestamp 1649977179
transform 1 0 14444 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_173
timestamp 1649977179
transform 1 0 17020 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_185
timestamp 1649977179
transform 1 0 18124 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_193
timestamp 1649977179
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_201
timestamp 1649977179
transform 1 0 19596 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_207
timestamp 1649977179
transform 1 0 20148 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_229
timestamp 1649977179
transform 1 0 22172 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_238
timestamp 1649977179
transform 1 0 23000 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1649977179
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_261
timestamp 1649977179
transform 1 0 25116 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_273
timestamp 1649977179
transform 1 0 26220 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_281
timestamp 1649977179
transform 1 0 26956 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_284
timestamp 1649977179
transform 1 0 27232 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1649977179
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_317
timestamp 1649977179
transform 1 0 30268 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_331
timestamp 1649977179
transform 1 0 31556 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_351
timestamp 1649977179
transform 1 0 33396 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1649977179
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_373
timestamp 1649977179
transform 1 0 35420 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_385
timestamp 1649977179
transform 1 0 36524 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_397
timestamp 1649977179
transform 1 0 37628 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_409
timestamp 1649977179
transform 1 0 38732 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_417
timestamp 1649977179
transform 1 0 39468 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_31
timestamp 1649977179
transform 1 0 3956 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_40
timestamp 1649977179
transform 1 0 4784 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_52
timestamp 1649977179
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_72
timestamp 1649977179
transform 1 0 7728 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_84
timestamp 1649977179
transform 1 0 8832 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_96
timestamp 1649977179
transform 1 0 9936 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1649977179
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_129
timestamp 1649977179
transform 1 0 12972 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_140
timestamp 1649977179
transform 1 0 13984 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_152
timestamp 1649977179
transform 1 0 15088 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1649977179
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_174
timestamp 1649977179
transform 1 0 17112 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_186
timestamp 1649977179
transform 1 0 18216 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_200
timestamp 1649977179
transform 1 0 19504 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_212
timestamp 1649977179
transform 1 0 20608 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_218
timestamp 1649977179
transform 1 0 21160 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_241
timestamp 1649977179
transform 1 0 23276 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_253
timestamp 1649977179
transform 1 0 24380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_257
timestamp 1649977179
transform 1 0 24748 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_266
timestamp 1649977179
transform 1 0 25576 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_272
timestamp 1649977179
transform 1 0 26128 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_313
timestamp 1649977179
transform 1 0 29900 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_327
timestamp 1649977179
transform 1 0 31188 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_340
timestamp 1649977179
transform 1 0 32384 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_352
timestamp 1649977179
transform 1 0 33488 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_360
timestamp 1649977179
transform 1 0 34224 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_365
timestamp 1649977179
transform 1 0 34684 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_377
timestamp 1649977179
transform 1 0 35788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1649977179
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_43
timestamp 1649977179
transform 1 0 5060 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_49
timestamp 1649977179
transform 1 0 5612 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_57
timestamp 1649977179
transform 1 0 6348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_63
timestamp 1649977179
transform 1 0 6900 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_75
timestamp 1649977179
transform 1 0 8004 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_87
timestamp 1649977179
transform 1 0 9108 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_101
timestamp 1649977179
transform 1 0 10396 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_113
timestamp 1649977179
transform 1 0 11500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_119
timestamp 1649977179
transform 1 0 12052 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_123
timestamp 1649977179
transform 1 0 12420 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_131
timestamp 1649977179
transform 1 0 13156 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_173
timestamp 1649977179
transform 1 0 17020 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1649977179
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_201
timestamp 1649977179
transform 1 0 19596 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_204
timestamp 1649977179
transform 1 0 19872 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_218
timestamp 1649977179
transform 1 0 21160 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_230
timestamp 1649977179
transform 1 0 22264 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_242
timestamp 1649977179
transform 1 0 23368 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1649977179
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_262
timestamp 1649977179
transform 1 0 25208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_266
timestamp 1649977179
transform 1 0 25576 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_283
timestamp 1649977179
transform 1 0 27140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_295
timestamp 1649977179
transform 1 0 28244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_318
timestamp 1649977179
transform 1 0 30360 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_338
timestamp 1649977179
transform 1 0 32200 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_350
timestamp 1649977179
transform 1 0 33304 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_362
timestamp 1649977179
transform 1 0 34408 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_617
timestamp 1649977179
transform 1 0 57868 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_621
timestamp 1649977179
transform 1 0 58236 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_35
timestamp 1649977179
transform 1 0 4324 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_41
timestamp 1649977179
transform 1 0 4876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_53
timestamp 1649977179
transform 1 0 5980 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_73
timestamp 1649977179
transform 1 0 7820 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_87
timestamp 1649977179
transform 1 0 9108 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_95
timestamp 1649977179
transform 1 0 9844 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_106
timestamp 1649977179
transform 1 0 10856 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_118
timestamp 1649977179
transform 1 0 11960 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_134
timestamp 1649977179
transform 1 0 13432 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_138
timestamp 1649977179
transform 1 0 13800 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_141
timestamp 1649977179
transform 1 0 14076 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_151
timestamp 1649977179
transform 1 0 14996 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_163
timestamp 1649977179
transform 1 0 16100 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_187
timestamp 1649977179
transform 1 0 18308 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_199
timestamp 1649977179
transform 1 0 19412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_211
timestamp 1649977179
transform 1 0 20516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_229
timestamp 1649977179
transform 1 0 22172 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_232
timestamp 1649977179
transform 1 0 22448 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_243
timestamp 1649977179
transform 1 0 23460 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_251
timestamp 1649977179
transform 1 0 24196 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_255
timestamp 1649977179
transform 1 0 24564 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_265
timestamp 1649977179
transform 1 0 25484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_277
timestamp 1649977179
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_287
timestamp 1649977179
transform 1 0 27508 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_295
timestamp 1649977179
transform 1 0 28244 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_301
timestamp 1649977179
transform 1 0 28796 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_309
timestamp 1649977179
transform 1 0 29532 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_313
timestamp 1649977179
transform 1 0 29900 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_325
timestamp 1649977179
transform 1 0 31004 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 1649977179
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_45
timestamp 1649977179
transform 1 0 5244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_57
timestamp 1649977179
transform 1 0 6348 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_60
timestamp 1649977179
transform 1 0 6624 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_72
timestamp 1649977179
transform 1 0 7728 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_92
timestamp 1649977179
transform 1 0 9568 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_112
timestamp 1649977179
transform 1 0 11408 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_136
timestamp 1649977179
transform 1 0 13616 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_149
timestamp 1649977179
transform 1 0 14812 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_158
timestamp 1649977179
transform 1 0 15640 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_164
timestamp 1649977179
transform 1 0 16192 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_170
timestamp 1649977179
transform 1 0 16744 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_176
timestamp 1649977179
transform 1 0 17296 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_179
timestamp 1649977179
transform 1 0 17572 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_187
timestamp 1649977179
transform 1 0 18308 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_191
timestamp 1649977179
transform 1 0 18676 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_229
timestamp 1649977179
transform 1 0 22172 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_234
timestamp 1649977179
transform 1 0 22632 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_240
timestamp 1649977179
transform 1 0 23184 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_263
timestamp 1649977179
transform 1 0 25300 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_272
timestamp 1649977179
transform 1 0 26128 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_280
timestamp 1649977179
transform 1 0 26864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_285
timestamp 1649977179
transform 1 0 27324 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_297
timestamp 1649977179
transform 1 0 28428 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1649977179
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_314
timestamp 1649977179
transform 1 0 29992 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_322
timestamp 1649977179
transform 1 0 30728 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_330
timestamp 1649977179
transform 1 0 31464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_344
timestamp 1649977179
transform 1 0 32752 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_352
timestamp 1649977179
transform 1 0 33488 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_360
timestamp 1649977179
transform 1 0 34224 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_382
timestamp 1649977179
transform 1 0 36248 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_394
timestamp 1649977179
transform 1 0 37352 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_406
timestamp 1649977179
transform 1 0 38456 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_418
timestamp 1649977179
transform 1 0 39560 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_617
timestamp 1649977179
transform 1 0 57868 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_621
timestamp 1649977179
transform 1 0 58236 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_67
timestamp 1649977179
transform 1 0 7268 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_76
timestamp 1649977179
transform 1 0 8096 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_88
timestamp 1649977179
transform 1 0 9200 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_100
timestamp 1649977179
transform 1 0 10304 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_117
timestamp 1649977179
transform 1 0 11868 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_122
timestamp 1649977179
transform 1 0 12328 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_136
timestamp 1649977179
transform 1 0 13616 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_140
timestamp 1649977179
transform 1 0 13984 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_157
timestamp 1649977179
transform 1 0 15548 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_165
timestamp 1649977179
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_177
timestamp 1649977179
transform 1 0 17388 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_189
timestamp 1649977179
transform 1 0 18492 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_198
timestamp 1649977179
transform 1 0 19320 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_202
timestamp 1649977179
transform 1 0 19688 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_235
timestamp 1649977179
transform 1 0 22724 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_241
timestamp 1649977179
transform 1 0 23276 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_267
timestamp 1649977179
transform 1 0 25668 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_276
timestamp 1649977179
transform 1 0 26496 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_283
timestamp 1649977179
transform 1 0 27140 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_287
timestamp 1649977179
transform 1 0 27508 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_304
timestamp 1649977179
transform 1 0 29072 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_316
timestamp 1649977179
transform 1 0 30176 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_332
timestamp 1649977179
transform 1 0 31648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_350
timestamp 1649977179
transform 1 0 33304 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_356
timestamp 1649977179
transform 1 0 33856 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_368
timestamp 1649977179
transform 1 0 34960 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_377
timestamp 1649977179
transform 1 0 35788 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_389
timestamp 1649977179
transform 1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_44
timestamp 1649977179
transform 1 0 5152 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_52
timestamp 1649977179
transform 1 0 5888 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_69
timestamp 1649977179
transform 1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1649977179
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_113
timestamp 1649977179
transform 1 0 11500 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_116
timestamp 1649977179
transform 1 0 11776 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_126
timestamp 1649977179
transform 1 0 12696 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_134
timestamp 1649977179
transform 1 0 13432 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_157
timestamp 1649977179
transform 1 0 15548 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_174
timestamp 1649977179
transform 1 0 17112 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_182
timestamp 1649977179
transform 1 0 17848 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1649977179
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_208
timestamp 1649977179
transform 1 0 20240 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_228
timestamp 1649977179
transform 1 0 22080 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_234
timestamp 1649977179
transform 1 0 22632 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_242
timestamp 1649977179
transform 1 0 23368 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1649977179
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_269
timestamp 1649977179
transform 1 0 25852 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_281
timestamp 1649977179
transform 1 0 26956 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_287
timestamp 1649977179
transform 1 0 27508 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_293
timestamp 1649977179
transform 1 0 28060 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_296
timestamp 1649977179
transform 1 0 28336 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_311
timestamp 1649977179
transform 1 0 29716 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_323
timestamp 1649977179
transform 1 0 30820 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_331
timestamp 1649977179
transform 1 0 31556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_336
timestamp 1649977179
transform 1 0 32016 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1649977179
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_385
timestamp 1649977179
transform 1 0 36524 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_397
timestamp 1649977179
transform 1 0 37628 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_409
timestamp 1649977179
transform 1 0 38732 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_417
timestamp 1649977179
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1649977179
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1649977179
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_11
timestamp 1649977179
transform 1 0 2116 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_30
timestamp 1649977179
transform 1 0 3864 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_42
timestamp 1649977179
transform 1 0 4968 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_59
timestamp 1649977179
transform 1 0 6532 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_71
timestamp 1649977179
transform 1 0 7636 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_83
timestamp 1649977179
transform 1 0 8740 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_90
timestamp 1649977179
transform 1 0 9384 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_102
timestamp 1649977179
transform 1 0 10488 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_107
timestamp 1649977179
transform 1 0 10948 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_120
timestamp 1649977179
transform 1 0 12144 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_128
timestamp 1649977179
transform 1 0 12880 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_138
timestamp 1649977179
transform 1 0 13800 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_150
timestamp 1649977179
transform 1 0 14904 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_162
timestamp 1649977179
transform 1 0 16008 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_173
timestamp 1649977179
transform 1 0 17020 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_182
timestamp 1649977179
transform 1 0 17848 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_190
timestamp 1649977179
transform 1 0 18584 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_201
timestamp 1649977179
transform 1 0 19596 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_213
timestamp 1649977179
transform 1 0 20700 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_219
timestamp 1649977179
transform 1 0 21252 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_235
timestamp 1649977179
transform 1 0 22724 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_241
timestamp 1649977179
transform 1 0 23276 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_267
timestamp 1649977179
transform 1 0 25668 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1649977179
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_298
timestamp 1649977179
transform 1 0 28520 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_307
timestamp 1649977179
transform 1 0 29348 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_311
timestamp 1649977179
transform 1 0 29716 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_314
timestamp 1649977179
transform 1 0 29992 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_326
timestamp 1649977179
transform 1 0 31096 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_332
timestamp 1649977179
transform 1 0 31648 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_348
timestamp 1649977179
transform 1 0 33120 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_354
timestamp 1649977179
transform 1 0 33672 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_357
timestamp 1649977179
transform 1 0 33948 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_369
timestamp 1649977179
transform 1 0 35052 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_381
timestamp 1649977179
transform 1 0 36156 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_389
timestamp 1649977179
transform 1 0 36892 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_621
timestamp 1649977179
transform 1 0 58236 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_12
timestamp 1649977179
transform 1 0 2208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_24
timestamp 1649977179
transform 1 0 3312 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_62
timestamp 1649977179
transform 1 0 6808 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_80
timestamp 1649977179
transform 1 0 8464 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_93
timestamp 1649977179
transform 1 0 9660 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_105
timestamp 1649977179
transform 1 0 10764 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_114
timestamp 1649977179
transform 1 0 11592 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_125
timestamp 1649977179
transform 1 0 12604 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_136
timestamp 1649977179
transform 1 0 13616 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_213
timestamp 1649977179
transform 1 0 20700 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_225
timestamp 1649977179
transform 1 0 21804 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_237
timestamp 1649977179
transform 1 0 22908 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_249
timestamp 1649977179
transform 1 0 24012 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_280
timestamp 1649977179
transform 1 0 26864 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_292
timestamp 1649977179
transform 1 0 27968 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1649977179
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_313
timestamp 1649977179
transform 1 0 29900 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_319
timestamp 1649977179
transform 1 0 30452 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_339
timestamp 1649977179
transform 1 0 32292 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_359
timestamp 1649977179
transform 1 0 34132 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1649977179
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1649977179
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_11
timestamp 1649977179
transform 1 0 2116 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_30
timestamp 1649977179
transform 1 0 3864 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_36
timestamp 1649977179
transform 1 0 4416 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_52
timestamp 1649977179
transform 1 0 5888 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_59
timestamp 1649977179
transform 1 0 6532 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_68
timestamp 1649977179
transform 1 0 7360 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_80
timestamp 1649977179
transform 1 0 8464 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_106
timestamp 1649977179
transform 1 0 10856 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_67_115
timestamp 1649977179
transform 1 0 11684 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_127
timestamp 1649977179
transform 1 0 12788 0 -1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_145
timestamp 1649977179
transform 1 0 14444 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_157
timestamp 1649977179
transform 1 0 15548 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_165
timestamp 1649977179
transform 1 0 16284 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1649977179
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_289
timestamp 1649977179
transform 1 0 27692 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_311
timestamp 1649977179
transform 1 0 29716 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_331
timestamp 1649977179
transform 1 0 31556 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_621
timestamp 1649977179
transform 1 0 58236 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_37
timestamp 1649977179
transform 1 0 4508 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_50
timestamp 1649977179
transform 1 0 5704 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_70
timestamp 1649977179
transform 1 0 7544 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_82
timestamp 1649977179
transform 1 0 8648 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_105
timestamp 1649977179
transform 1 0 10764 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_114
timestamp 1649977179
transform 1 0 11592 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_122
timestamp 1649977179
transform 1 0 12328 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_136
timestamp 1649977179
transform 1 0 13616 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_159
timestamp 1649977179
transform 1 0 15732 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_167
timestamp 1649977179
transform 1 0 16468 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_185
timestamp 1649977179
transform 1 0 18124 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_192
timestamp 1649977179
transform 1 0 18768 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_213
timestamp 1649977179
transform 1 0 20700 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_225
timestamp 1649977179
transform 1 0 21804 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_237
timestamp 1649977179
transform 1 0 22908 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_249
timestamp 1649977179
transform 1 0 24012 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_269
timestamp 1649977179
transform 1 0 25852 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_281
timestamp 1649977179
transform 1 0 26956 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_299
timestamp 1649977179
transform 1 0 28612 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_313
timestamp 1649977179
transform 1 0 29900 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_319
timestamp 1649977179
transform 1 0 30452 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_331
timestamp 1649977179
transform 1 0 31556 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_340
timestamp 1649977179
transform 1 0 32384 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_352
timestamp 1649977179
transform 1 0 33488 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_31
timestamp 1649977179
transform 1 0 3956 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_40
timestamp 1649977179
transform 1 0 4784 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_46
timestamp 1649977179
transform 1 0 5336 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_52
timestamp 1649977179
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_65
timestamp 1649977179
transform 1 0 7084 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_85
timestamp 1649977179
transform 1 0 8924 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_121
timestamp 1649977179
transform 1 0 12236 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_127
timestamp 1649977179
transform 1 0 12788 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_139
timestamp 1649977179
transform 1 0 13892 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_156
timestamp 1649977179
transform 1 0 15456 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_183
timestamp 1649977179
transform 1 0 17940 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_207
timestamp 1649977179
transform 1 0 20148 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_213
timestamp 1649977179
transform 1 0 20700 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_220
timestamp 1649977179
transform 1 0 21344 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_233
timestamp 1649977179
transform 1 0 22540 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_242
timestamp 1649977179
transform 1 0 23368 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_246
timestamp 1649977179
transform 1 0 23736 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_263
timestamp 1649977179
transform 1 0 25300 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_275
timestamp 1649977179
transform 1 0 26404 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_301
timestamp 1649977179
transform 1 0 28796 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_313
timestamp 1649977179
transform 1 0 29900 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_325
timestamp 1649977179
transform 1 0 31004 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_333
timestamp 1649977179
transform 1 0 31740 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_60
timestamp 1649977179
transform 1 0 6624 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_64
timestamp 1649977179
transform 1 0 6992 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_67
timestamp 1649977179
transform 1 0 7268 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_79
timestamp 1649977179
transform 1 0 8372 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_114
timestamp 1649977179
transform 1 0 11592 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_70_134
timestamp 1649977179
transform 1 0 13432 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_148
timestamp 1649977179
transform 1 0 14720 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_160
timestamp 1649977179
transform 1 0 15824 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_178
timestamp 1649977179
transform 1 0 17480 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_186
timestamp 1649977179
transform 1 0 18216 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_192
timestamp 1649977179
transform 1 0 18768 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_205
timestamp 1649977179
transform 1 0 19964 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_213
timestamp 1649977179
transform 1 0 20700 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_230
timestamp 1649977179
transform 1 0 22264 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_236
timestamp 1649977179
transform 1 0 22816 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_258
timestamp 1649977179
transform 1 0 24840 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_270
timestamp 1649977179
transform 1 0 25944 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_282
timestamp 1649977179
transform 1 0 27048 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_294
timestamp 1649977179
transform 1 0 28152 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_306
timestamp 1649977179
transform 1 0 29256 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_340
timestamp 1649977179
transform 1 0 32384 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_352
timestamp 1649977179
transform 1 0 33488 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_617
timestamp 1649977179
transform 1 0 57868 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_621
timestamp 1649977179
transform 1 0 58236 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_89
timestamp 1649977179
transform 1 0 9292 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_100
timestamp 1649977179
transform 1 0 10304 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_106
timestamp 1649977179
transform 1 0 10856 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_135
timestamp 1649977179
transform 1 0 13524 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_141
timestamp 1649977179
transform 1 0 14076 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_153
timestamp 1649977179
transform 1 0 15180 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_163
timestamp 1649977179
transform 1 0 16100 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_171
timestamp 1649977179
transform 1 0 16836 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_183
timestamp 1649977179
transform 1 0 17940 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_202
timestamp 1649977179
transform 1 0 19688 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_214
timestamp 1649977179
transform 1 0 20792 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_220
timestamp 1649977179
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_230
timestamp 1649977179
transform 1 0 22264 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_244
timestamp 1649977179
transform 1 0 23552 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_250
timestamp 1649977179
transform 1 0 24104 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_262
timestamp 1649977179
transform 1 0 25208 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_274
timestamp 1649977179
transform 1 0 26312 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1649977179
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_617
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_117
timestamp 1649977179
transform 1 0 11868 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_124
timestamp 1649977179
transform 1 0 12512 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_136
timestamp 1649977179
transform 1 0 13616 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_143
timestamp 1649977179
transform 1 0 14260 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_152
timestamp 1649977179
transform 1 0 15088 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_164
timestamp 1649977179
transform 1 0 16192 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_170
timestamp 1649977179
transform 1 0 16744 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_182
timestamp 1649977179
transform 1 0 17848 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_194
timestamp 1649977179
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_202
timestamp 1649977179
transform 1 0 19688 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_208
timestamp 1649977179
transform 1 0 20240 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_220
timestamp 1649977179
transform 1 0 21344 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_232
timestamp 1649977179
transform 1 0 22448 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_246
timestamp 1649977179
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_617
timestamp 1649977179
transform 1 0 57868 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_621
timestamp 1649977179
transform 1 0 58236 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_73_133
timestamp 1649977179
transform 1 0 13340 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_145
timestamp 1649977179
transform 1 0 14444 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_155
timestamp 1649977179
transform 1 0 15364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1649977179
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1649977179
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1649977179
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1649977179
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1649977179
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1649977179
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1649977179
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1649977179
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1649977179
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_621
timestamp 1649977179
transform 1 0 58236 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1649977179
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1649977179
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1649977179
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_621
timestamp 1649977179
transform 1 0 58236 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1649977179
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1649977179
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1649977179
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_617
timestamp 1649977179
transform 1 0 57868 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_621
timestamp 1649977179
transform 1 0 58236 0 1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1649977179
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1649977179
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_617
timestamp 1649977179
transform 1 0 57868 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_621
timestamp 1649977179
transform 1 0 58236 0 1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1649977179
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1649977179
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1649977179
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1649977179
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1649977179
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1649977179
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1649977179
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1649977179
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1649977179
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_621
timestamp 1649977179
transform 1 0 58236 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1649977179
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1649977179
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1649977179
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1649977179
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1649977179
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1649977179
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1649977179
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1649977179
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1649977179
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1649977179
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1649977179
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1649977179
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1649977179
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1649977179
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1649977179
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1649977179
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_621
timestamp 1649977179
transform 1 0 58236 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1649977179
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1649977179
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1649977179
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1649977179
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1649977179
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1649977179
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1649977179
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1649977179
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1649977179
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1649977179
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1649977179
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1649977179
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1649977179
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1649977179
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1649977179
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1649977179
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1649977179
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1649977179
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1649977179
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1649977179
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1649977179
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1649977179
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1649977179
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1649977179
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1649977179
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1649977179
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1649977179
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1649977179
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1649977179
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1649977179
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1649977179
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1649977179
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1649977179
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_617
timestamp 1649977179
transform 1 0 57868 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_621
timestamp 1649977179
transform 1 0 58236 0 1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1649977179
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1649977179
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1649977179
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1649977179
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1649977179
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1649977179
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1649977179
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1649977179
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1649977179
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1649977179
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1649977179
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1649977179
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1649977179
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1649977179
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1649977179
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1649977179
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_92_617
timestamp 1649977179
transform 1 0 57868 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_621
timestamp 1649977179
transform 1 0 58236 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1649977179
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1649977179
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1649977179
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1649977179
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1649977179
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1649977179
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1649977179
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1649977179
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1649977179
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1649977179
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1649977179
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1649977179
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1649977179
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1649977179
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1649977179
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1649977179
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1649977179
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1649977179
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1649977179
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1649977179
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1649977179
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1649977179
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1649977179
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1649977179
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1649977179
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_621
timestamp 1649977179
transform 1 0 58236 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1649977179
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1649977179
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1649977179
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1649977179
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1649977179
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1649977179
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1649977179
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1649977179
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1649977179
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_173
timestamp 1649977179
transform 1 0 17020 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_176
timestamp 1649977179
transform 1 0 17296 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_188
timestamp 1649977179
transform 1 0 18400 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_97_196
timestamp 1649977179
transform 1 0 19136 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_97_202
timestamp 1649977179
transform 1 0 19688 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_214
timestamp 1649977179
transform 1 0 20792 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_222
timestamp 1649977179
transform 1 0 21528 0 -1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1649977179
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1649977179
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1649977179
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1649977179
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1649977179
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1649977179
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1649977179
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1649977179
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1649977179
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1649977179
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1649977179
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1649977179
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_97_617
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_621
timestamp 1649977179
transform 1 0 58236 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1649977179
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1649977179
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1649977179
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_153
timestamp 1649977179
transform 1 0 15180 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_98_161
timestamp 1649977179
transform 1 0 15916 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_98_166
timestamp 1649977179
transform 1 0 16376 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_170
timestamp 1649977179
transform 1 0 16744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_174
timestamp 1649977179
transform 1 0 17112 0 1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_182
timestamp 1649977179
transform 1 0 17848 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_185
timestamp 1649977179
transform 1 0 18124 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_192
timestamp 1649977179
transform 1 0 18768 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_197
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_201
timestamp 1649977179
transform 1 0 19596 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_205
timestamp 1649977179
transform 1 0 19964 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_211
timestamp 1649977179
transform 1 0 20516 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_217
timestamp 1649977179
transform 1 0 21068 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_98_229
timestamp 1649977179
transform 1 0 22172 0 1 55488
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_98_234
timestamp 1649977179
transform 1 0 22632 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_246
timestamp 1649977179
transform 1 0 23736 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_98_253
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_98_259
timestamp 1649977179
transform 1 0 24932 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_98_263
timestamp 1649977179
transform 1 0 25300 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_98_266
timestamp 1649977179
transform 1 0 25576 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_272
timestamp 1649977179
transform 1 0 26128 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_276
timestamp 1649977179
transform 1 0 26496 0 1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_282
timestamp 1649977179
transform 1 0 27048 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_294
timestamp 1649977179
transform 1 0 28152 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_98_306
timestamp 1649977179
transform 1 0 29256 0 1 55488
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1649977179
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1649977179
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1649977179
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1649977179
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1649977179
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1649977179
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1649977179
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1649977179
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1649977179
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1649977179
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1649977179
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1649977179
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1649977179
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1649977179
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1649977179
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1649977179
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1649977179
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1649977179
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1649977179
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1649977179
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_125
timestamp 1649977179
transform 1 0 12604 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_133
timestamp 1649977179
transform 1 0 13340 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_138
timestamp 1649977179
transform 1 0 13800 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_144
timestamp 1649977179
transform 1 0 14352 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_156
timestamp 1649977179
transform 1 0 15456 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_160
timestamp 1649977179
transform 1 0 15824 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_164
timestamp 1649977179
transform 1 0 16192 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_171
timestamp 1649977179
transform 1 0 16836 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_178
timestamp 1649977179
transform 1 0 17480 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_185
timestamp 1649977179
transform 1 0 18124 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_192
timestamp 1649977179
transform 1 0 18768 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_199
timestamp 1649977179
transform 1 0 19412 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_206
timestamp 1649977179
transform 1 0 20056 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_213
timestamp 1649977179
transform 1 0 20700 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_220
timestamp 1649977179
transform 1 0 21344 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_230
timestamp 1649977179
transform 1 0 22264 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_237
timestamp 1649977179
transform 1 0 22908 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_241
timestamp 1649977179
transform 1 0 23276 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_244
timestamp 1649977179
transform 1 0 23552 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_251
timestamp 1649977179
transform 1 0 24196 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_99_262
timestamp 1649977179
transform 1 0 25208 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_269
timestamp 1649977179
transform 1 0 25852 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_276
timestamp 1649977179
transform 1 0 26496 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_281
timestamp 1649977179
transform 1 0 26956 0 -1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_286
timestamp 1649977179
transform 1 0 27416 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_292
timestamp 1649977179
transform 1 0 27968 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_304
timestamp 1649977179
transform 1 0 29072 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_99_313
timestamp 1649977179
transform 1 0 29900 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_319
timestamp 1649977179
transform 1 0 30452 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_325
timestamp 1649977179
transform 1 0 31004 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_332
timestamp 1649977179
transform 1 0 31648 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_340
timestamp 1649977179
transform 1 0 32384 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_346
timestamp 1649977179
transform 1 0 32936 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_354
timestamp 1649977179
transform 1 0 33672 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_360
timestamp 1649977179
transform 1 0 34224 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_99_366
timestamp 1649977179
transform 1 0 34776 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_374
timestamp 1649977179
transform 1 0 35512 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_380
timestamp 1649977179
transform 1 0 36064 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_99_386
timestamp 1649977179
transform 1 0 36616 0 -1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_461
timestamp 1649977179
transform 1 0 43516 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_99_469
timestamp 1649977179
transform 1 0 44252 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_472
timestamp 1649977179
transform 1 0 44528 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_479
timestamp 1649977179
transform 1 0 45172 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_486
timestamp 1649977179
transform 1 0 45816 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_99_492
timestamp 1649977179
transform 1 0 46368 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_99_617
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_621
timestamp 1649977179
transform 1 0 58236 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1649977179
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1649977179
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1649977179
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1649977179
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1649977179
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1649977179
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1649977179
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_177
timestamp 1649977179
transform 1 0 17388 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_183
timestamp 1649977179
transform 1 0 17940 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_100_190
timestamp 1649977179
transform 1 0 18584 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_100_200
timestamp 1649977179
transform 1 0 19504 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_100_208
timestamp 1649977179
transform 1 0 20240 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_212
timestamp 1649977179
transform 1 0 20608 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_215
timestamp 1649977179
transform 1 0 20884 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_227
timestamp 1649977179
transform 1 0 21988 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_232
timestamp 1649977179
transform 1 0 22448 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_244
timestamp 1649977179
transform 1 0 23552 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_100_253
timestamp 1649977179
transform 1 0 24380 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_261
timestamp 1649977179
transform 1 0 25116 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_265
timestamp 1649977179
transform 1 0 25484 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_272
timestamp 1649977179
transform 1 0 26128 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_278
timestamp 1649977179
transform 1 0 26680 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_290
timestamp 1649977179
transform 1 0 27784 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_302
timestamp 1649977179
transform 1 0 28888 0 1 56576
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1649977179
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1649977179
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1649977179
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1649977179
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1649977179
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1649977179
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1649977179
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_100_445
timestamp 1649977179
transform 1 0 42044 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_450
timestamp 1649977179
transform 1 0 42504 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_462
timestamp 1649977179
transform 1 0 43608 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_474
timestamp 1649977179
transform 1 0 44712 0 1 56576
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1649977179
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1649977179
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1649977179
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1649977179
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1649977179
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_100_609
timestamp 1649977179
transform 1 0 57132 0 1 56576
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_614
timestamp 1649977179
transform 1 0 57592 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_100_621
timestamp 1649977179
transform 1 0 58236 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_3
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_7
timestamp 1649977179
transform 1 0 1748 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_12
timestamp 1649977179
transform 1 0 2208 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_18
timestamp 1649977179
transform 1 0 2760 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_26
timestamp 1649977179
transform 1 0 3496 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_33
timestamp 1649977179
transform 1 0 4140 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_41
timestamp 1649977179
transform 1 0 4876 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_46
timestamp 1649977179
transform 1 0 5336 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_54
timestamp 1649977179
transform 1 0 6072 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_63
timestamp 1649977179
transform 1 0 6900 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_75
timestamp 1649977179
transform 1 0 8004 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_80
timestamp 1649977179
transform 1 0 8464 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_85
timestamp 1649977179
transform 1 0 8924 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_97
timestamp 1649977179
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_109
timestamp 1649977179
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_117
timestamp 1649977179
transform 1 0 11868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_125
timestamp 1649977179
transform 1 0 12604 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_101_131
timestamp 1649977179
transform 1 0 13156 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_139
timestamp 1649977179
transform 1 0 13892 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_101_141
timestamp 1649977179
transform 1 0 14076 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_101_148
timestamp 1649977179
transform 1 0 14720 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_160
timestamp 1649977179
transform 1 0 15824 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_173
timestamp 1649977179
transform 1 0 17020 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_177
timestamp 1649977179
transform 1 0 17388 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_182
timestamp 1649977179
transform 1 0 17848 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_192
timestamp 1649977179
transform 1 0 18768 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_201
timestamp 1649977179
transform 1 0 19596 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_207
timestamp 1649977179
transform 1 0 20148 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_211
timestamp 1649977179
transform 1 0 20516 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_216
timestamp 1649977179
transform 1 0 20976 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_225
timestamp 1649977179
transform 1 0 21804 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_233
timestamp 1649977179
transform 1 0 22540 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_245
timestamp 1649977179
transform 1 0 23644 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_251
timestamp 1649977179
transform 1 0 24196 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_257
timestamp 1649977179
transform 1 0 24748 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_267
timestamp 1649977179
transform 1 0 25668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_279
timestamp 1649977179
transform 1 0 26772 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_285
timestamp 1649977179
transform 1 0 27324 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_301
timestamp 1649977179
transform 1 0 28796 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_307
timestamp 1649977179
transform 1 0 29348 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_309
timestamp 1649977179
transform 1 0 29532 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_313
timestamp 1649977179
transform 1 0 29900 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_318
timestamp 1649977179
transform 1 0 30360 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_330
timestamp 1649977179
transform 1 0 31464 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_341
timestamp 1649977179
transform 1 0 32476 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_347
timestamp 1649977179
transform 1 0 33028 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_352
timestamp 1649977179
transform 1 0 33488 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_369
timestamp 1649977179
transform 1 0 35052 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_381
timestamp 1649977179
transform 1 0 36156 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_386
timestamp 1649977179
transform 1 0 36616 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_101_393
timestamp 1649977179
transform 1 0 37260 0 -1 57664
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_101_403
timestamp 1649977179
transform 1 0 38180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_415
timestamp 1649977179
transform 1 0 39284 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_419
timestamp 1649977179
transform 1 0 39652 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_425
timestamp 1649977179
transform 1 0 40204 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_101_437
timestamp 1649977179
transform 1 0 41308 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_445
timestamp 1649977179
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_101_449
timestamp 1649977179
transform 1 0 42412 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_454
timestamp 1649977179
transform 1 0 42872 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_466
timestamp 1649977179
transform 1 0 43976 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_471
timestamp 1649977179
transform 1 0 44436 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_475
timestamp 1649977179
transform 1 0 44804 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_477
timestamp 1649977179
transform 1 0 44988 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_483
timestamp 1649977179
transform 1 0 45540 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_101_488
timestamp 1649977179
transform 1 0 46000 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_500
timestamp 1649977179
transform 1 0 47104 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_509
timestamp 1649977179
transform 1 0 47932 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_517
timestamp 1649977179
transform 1 0 48668 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_521
timestamp 1649977179
transform 1 0 49036 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_529
timestamp 1649977179
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_101_533
timestamp 1649977179
transform 1 0 50140 0 -1 57664
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_101_538
timestamp 1649977179
transform 1 0 50600 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_550
timestamp 1649977179
transform 1 0 51704 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_555
timestamp 1649977179
transform 1 0 52164 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_559
timestamp 1649977179
transform 1 0 52532 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_561
timestamp 1649977179
transform 1 0 52716 0 -1 57664
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_572
timestamp 1649977179
transform 1 0 53728 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_584
timestamp 1649977179
transform 1 0 54832 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_592
timestamp 1649977179
transform 1 0 55568 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_101_600
timestamp 1649977179
transform 1 0 56304 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_101_606
timestamp 1649977179
transform 1 0 56856 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_614
timestamp 1649977179
transform 1 0 57592 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_617
timestamp 1649977179
transform 1 0 57868 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_621
timestamp 1649977179
transform 1 0 58236 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0855_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4968 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0856_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6440 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or4_4  _0857_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10856 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _0858_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0859_
timestamp 1649977179
transform -1 0 7820 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0860_
timestamp 1649977179
transform 1 0 8188 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0861_
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0862_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _0863_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14996 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0864_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _0865_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _0866_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0867_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4416 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0868_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0869_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2944 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0870_
timestamp 1649977179
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0871_
timestamp 1649977179
transform -1 0 12420 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0872_
timestamp 1649977179
transform 1 0 2944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0873_
timestamp 1649977179
transform 1 0 4968 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0874_
timestamp 1649977179
transform -1 0 2760 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0875_
timestamp 1649977179
transform -1 0 2392 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0876_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1649977179
transform 1 0 2852 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0878_
timestamp 1649977179
transform 1 0 3680 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0879_
timestamp 1649977179
transform 1 0 4784 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0880_
timestamp 1649977179
transform 1 0 2024 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0881_
timestamp 1649977179
transform 1 0 2392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0882_
timestamp 1649977179
transform 1 0 3864 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0884_
timestamp 1649977179
transform 1 0 2208 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0885_
timestamp 1649977179
transform 1 0 5336 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0886_
timestamp 1649977179
transform 1 0 4508 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0887_
timestamp 1649977179
transform 1 0 1932 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0888_
timestamp 1649977179
transform -1 0 2852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0889_
timestamp 1649977179
transform -1 0 4324 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0890_
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1649977179
transform -1 0 2944 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0892_
timestamp 1649977179
transform -1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0893_
timestamp 1649977179
transform 1 0 9936 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0894_
timestamp 1649977179
transform 1 0 8004 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0895_
timestamp 1649977179
transform -1 0 9200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0896_
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0897_
timestamp 1649977179
transform -1 0 2944 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0898_
timestamp 1649977179
transform -1 0 1932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0899_
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0900_
timestamp 1649977179
transform 1 0 12972 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0901_
timestamp 1649977179
transform -1 0 14444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0902_
timestamp 1649977179
transform 1 0 2392 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0903_
timestamp 1649977179
transform -1 0 2576 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0904_
timestamp 1649977179
transform -1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0905_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0906_
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0907_
timestamp 1649977179
transform 1 0 6624 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0908_
timestamp 1649977179
transform 1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0909_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7268 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0910_
timestamp 1649977179
transform -1 0 14352 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0911_
timestamp 1649977179
transform 1 0 17848 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_4  _0912_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0913_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0914_
timestamp 1649977179
transform -1 0 11776 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0915_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8004 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0916_
timestamp 1649977179
transform -1 0 8464 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1649977179
transform -1 0 11960 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0918_
timestamp 1649977179
transform 1 0 9108 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0919_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4784 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0920_
timestamp 1649977179
transform 1 0 4968 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0921_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0922_
timestamp 1649977179
transform -1 0 7728 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0923_
timestamp 1649977179
transform -1 0 2208 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0924_
timestamp 1649977179
transform 1 0 4232 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0925_
timestamp 1649977179
transform -1 0 7820 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0926_
timestamp 1649977179
transform -1 0 5796 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0927_
timestamp 1649977179
transform 1 0 2576 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0928_
timestamp 1649977179
transform -1 0 8464 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0929_
timestamp 1649977179
transform -1 0 6808 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0930_
timestamp 1649977179
transform -1 0 5704 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _0931_
timestamp 1649977179
transform -1 0 10856 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0932_
timestamp 1649977179
transform -1 0 7360 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0933_
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0934_
timestamp 1649977179
transform -1 0 25484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0935_
timestamp 1649977179
transform 1 0 13524 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0936_
timestamp 1649977179
transform -1 0 12604 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1649977179
transform -1 0 12512 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0938_
timestamp 1649977179
transform 1 0 12696 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0939_
timestamp 1649977179
transform 1 0 12788 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1649977179
transform -1 0 26220 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0941_
timestamp 1649977179
transform 1 0 14904 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0942_
timestamp 1649977179
transform -1 0 16100 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0943_
timestamp 1649977179
transform -1 0 25208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0944_
timestamp 1649977179
transform 1 0 14628 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0945_
timestamp 1649977179
transform -1 0 16192 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0946_
timestamp 1649977179
transform -1 0 25024 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0947_
timestamp 1649977179
transform 1 0 14260 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0948_
timestamp 1649977179
transform 1 0 14444 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0949_
timestamp 1649977179
transform 1 0 24104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0950_
timestamp 1649977179
transform 1 0 12880 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0951_
timestamp 1649977179
transform 1 0 12880 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0952_
timestamp 1649977179
transform -1 0 17020 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0953_
timestamp 1649977179
transform 1 0 12512 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0954_
timestamp 1649977179
transform 1 0 13064 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0955_
timestamp 1649977179
transform 1 0 12880 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0956_
timestamp 1649977179
transform -1 0 13800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0958_
timestamp 1649977179
transform 1 0 13156 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _0959_
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0960_
timestamp 1649977179
transform -1 0 20976 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0961_
timestamp 1649977179
transform -1 0 30728 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0962_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29992 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0963_
timestamp 1649977179
transform 1 0 30176 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0964_
timestamp 1649977179
transform 1 0 17020 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0965_
timestamp 1649977179
transform 1 0 30820 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0966_
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0967_
timestamp 1649977179
transform -1 0 29992 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0968_
timestamp 1649977179
transform -1 0 30176 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0969_
timestamp 1649977179
transform -1 0 28796 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0970_
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0971_
timestamp 1649977179
transform -1 0 29256 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0972_
timestamp 1649977179
transform 1 0 27692 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0973_
timestamp 1649977179
transform 1 0 29900 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0974_
timestamp 1649977179
transform 1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0975_
timestamp 1649977179
transform -1 0 31188 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0976_
timestamp 1649977179
transform -1 0 31004 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0977_
timestamp 1649977179
transform 1 0 29808 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0978_
timestamp 1649977179
transform -1 0 31004 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0979_
timestamp 1649977179
transform 1 0 35328 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0980_
timestamp 1649977179
transform -1 0 34960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0981_
timestamp 1649977179
transform 1 0 35788 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0982_
timestamp 1649977179
transform -1 0 36800 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0983_
timestamp 1649977179
transform 1 0 35052 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0984_
timestamp 1649977179
transform -1 0 36616 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0985_
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0986_
timestamp 1649977179
transform -1 0 36616 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0987_
timestamp 1649977179
transform 1 0 35236 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0988_
timestamp 1649977179
transform -1 0 30084 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0989_
timestamp 1649977179
transform -1 0 36800 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0990_
timestamp 1649977179
transform 1 0 35972 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0991_
timestamp 1649977179
transform -1 0 36892 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0992_
timestamp 1649977179
transform 1 0 34960 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0993_
timestamp 1649977179
transform -1 0 34592 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0994_
timestamp 1649977179
transform -1 0 33856 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0995_
timestamp 1649977179
transform -1 0 33120 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _0996_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0997_
timestamp 1649977179
transform -1 0 21344 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0998_
timestamp 1649977179
transform 1 0 30084 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0999_
timestamp 1649977179
transform 1 0 30544 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1000_
timestamp 1649977179
transform -1 0 30912 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1001_
timestamp 1649977179
transform 1 0 29992 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1002_
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1649977179
transform 1 0 28612 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1004_
timestamp 1649977179
transform 1 0 28428 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1005_
timestamp 1649977179
transform -1 0 29348 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1006_
timestamp 1649977179
transform -1 0 31648 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1007_
timestamp 1649977179
transform 1 0 28336 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1008_
timestamp 1649977179
transform -1 0 28520 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1009_
timestamp 1649977179
transform 1 0 27232 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1649977179
transform 1 0 29992 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1011_
timestamp 1649977179
transform -1 0 31096 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1012_
timestamp 1649977179
transform 1 0 31924 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1013_
timestamp 1649977179
transform 1 0 30820 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1014_
timestamp 1649977179
transform 1 0 32384 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1015_
timestamp 1649977179
transform -1 0 32384 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1016_
timestamp 1649977179
transform -1 0 33304 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1017_
timestamp 1649977179
transform -1 0 33120 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1649977179
transform 1 0 33764 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1019_
timestamp 1649977179
transform 1 0 31832 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1020_
timestamp 1649977179
transform -1 0 35420 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1021_
timestamp 1649977179
transform 1 0 33764 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1022_
timestamp 1649977179
transform -1 0 34592 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1649977179
transform 1 0 35328 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1024_
timestamp 1649977179
transform -1 0 35052 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1025_
timestamp 1649977179
transform 1 0 33764 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1026_
timestamp 1649977179
transform -1 0 34960 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1027_
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1028_
timestamp 1649977179
transform 1 0 31924 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1029_
timestamp 1649977179
transform 1 0 32200 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1030_
timestamp 1649977179
transform 1 0 29716 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1031_
timestamp 1649977179
transform -1 0 31924 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _1032_
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1033_
timestamp 1649977179
transform -1 0 10488 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1034_
timestamp 1649977179
transform -1 0 9752 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1035_
timestamp 1649977179
transform 1 0 9476 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1036_
timestamp 1649977179
transform -1 0 8740 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1037_
timestamp 1649977179
transform 1 0 10672 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1038_
timestamp 1649977179
transform -1 0 17112 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1649977179
transform 1 0 5612 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1040_
timestamp 1649977179
transform 1 0 5520 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1041_
timestamp 1649977179
transform -1 0 7820 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1042_
timestamp 1649977179
transform -1 0 4784 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1043_
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1044_
timestamp 1649977179
transform -1 0 4784 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1045_
timestamp 1649977179
transform 1 0 2576 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1046_
timestamp 1649977179
transform 1 0 7912 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1047_
timestamp 1649977179
transform 1 0 6348 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1048_
timestamp 1649977179
transform 1 0 6440 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1049_
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1050_
timestamp 1649977179
transform -1 0 25116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1051_
timestamp 1649977179
transform -1 0 19320 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1052_
timestamp 1649977179
transform 1 0 7268 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1053_
timestamp 1649977179
transform 1 0 15824 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1054_
timestamp 1649977179
transform 1 0 17480 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1055_
timestamp 1649977179
transform 1 0 19780 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1056_
timestamp 1649977179
transform -1 0 20700 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1057_
timestamp 1649977179
transform 1 0 18308 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1058_
timestamp 1649977179
transform 1 0 20056 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1059_
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1060_
timestamp 1649977179
transform -1 0 19964 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 1649977179
transform 1 0 19688 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1062_
timestamp 1649977179
transform -1 0 20608 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1063_
timestamp 1649977179
transform -1 0 18584 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1064_
timestamp 1649977179
transform -1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1065_
timestamp 1649977179
transform -1 0 18032 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1066_
timestamp 1649977179
transform 1 0 15088 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1067_
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1068_
timestamp 1649977179
transform 1 0 14904 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1069_
timestamp 1649977179
transform -1 0 15640 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1070_
timestamp 1649977179
transform -1 0 18952 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1071_
timestamp 1649977179
transform -1 0 18492 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1072_
timestamp 1649977179
transform -1 0 16744 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1073_
timestamp 1649977179
transform -1 0 15824 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1074_
timestamp 1649977179
transform 1 0 16836 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1075_
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1076_
timestamp 1649977179
transform -1 0 10580 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1077_
timestamp 1649977179
transform 1 0 9200 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1078_
timestamp 1649977179
transform -1 0 9292 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1079_
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1080_
timestamp 1649977179
transform 1 0 11776 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1081_
timestamp 1649977179
transform 1 0 23092 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1082_
timestamp 1649977179
transform 1 0 11592 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1083_
timestamp 1649977179
transform -1 0 13800 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1084_
timestamp 1649977179
transform 1 0 12696 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1085_
timestamp 1649977179
transform -1 0 15364 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1086_
timestamp 1649977179
transform 1 0 14352 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1087_
timestamp 1649977179
transform -1 0 25300 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1088_
timestamp 1649977179
transform -1 0 23736 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1089_
timestamp 1649977179
transform 1 0 25668 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1090_
timestamp 1649977179
transform 1 0 26220 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1091_
timestamp 1649977179
transform 1 0 26036 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1092_
timestamp 1649977179
transform 1 0 24564 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1093_
timestamp 1649977179
transform 1 0 24748 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1094_
timestamp 1649977179
transform -1 0 23920 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1095_
timestamp 1649977179
transform -1 0 25576 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1096_
timestamp 1649977179
transform 1 0 23552 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1097_
timestamp 1649977179
transform -1 0 25116 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1098_
timestamp 1649977179
transform 1 0 23460 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1099_
timestamp 1649977179
transform -1 0 25116 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1649977179
transform 1 0 24196 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1101_
timestamp 1649977179
transform -1 0 25668 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1102_
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1103_
timestamp 1649977179
transform -1 0 25392 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1104_
timestamp 1649977179
transform 1 0 15916 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1105_
timestamp 1649977179
transform 1 0 20884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1106_
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1107_
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1108_
timestamp 1649977179
transform 1 0 23000 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1109_
timestamp 1649977179
transform -1 0 24656 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1110_
timestamp 1649977179
transform -1 0 23920 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1111_
timestamp 1649977179
transform -1 0 24840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1649977179
transform -1 0 24840 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1113_
timestamp 1649977179
transform -1 0 23920 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1114_
timestamp 1649977179
transform 1 0 23460 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1115_
timestamp 1649977179
transform 1 0 14720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1117_
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1118_
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1119_
timestamp 1649977179
transform -1 0 23920 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1120_
timestamp 1649977179
transform 1 0 23184 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1121_
timestamp 1649977179
transform 1 0 18308 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1122_
timestamp 1649977179
transform 1 0 26036 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1123_
timestamp 1649977179
transform -1 0 25668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1124_
timestamp 1649977179
transform 1 0 19136 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1125_
timestamp 1649977179
transform -1 0 25668 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1126_
timestamp 1649977179
transform -1 0 25484 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1649977179
transform 1 0 28796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1128_
timestamp 1649977179
transform 1 0 28244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1129_
timestamp 1649977179
transform -1 0 28244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1649977179
transform 1 0 31188 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1131_
timestamp 1649977179
transform 1 0 34040 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1132_
timestamp 1649977179
transform -1 0 33028 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1133_
timestamp 1649977179
transform -1 0 31648 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1134_
timestamp 1649977179
transform 1 0 30728 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1135_
timestamp 1649977179
transform 1 0 32476 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1136_
timestamp 1649977179
transform -1 0 33396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1137_
timestamp 1649977179
transform 1 0 29900 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1138_
timestamp 1649977179
transform 1 0 30084 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1139_
timestamp 1649977179
transform -1 0 31280 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1140_
timestamp 1649977179
transform 1 0 27048 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1649977179
transform 1 0 31188 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1142_
timestamp 1649977179
transform -1 0 32844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1143_
timestamp 1649977179
transform 1 0 27048 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1144_
timestamp 1649977179
transform 1 0 29532 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1145_
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1146_
timestamp 1649977179
transform 1 0 19872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1649977179
transform -1 0 22632 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1148_
timestamp 1649977179
transform -1 0 27692 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1149_
timestamp 1649977179
transform 1 0 21896 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1150_
timestamp 1649977179
transform 1 0 19872 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1151_
timestamp 1649977179
transform -1 0 26312 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1152_
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1153_
timestamp 1649977179
transform -1 0 19688 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1154_
timestamp 1649977179
transform 1 0 20056 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1155_
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1156_
timestamp 1649977179
transform -1 0 21068 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1157_
timestamp 1649977179
transform -1 0 16744 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1158_
timestamp 1649977179
transform 1 0 20148 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1159_
timestamp 1649977179
transform 1 0 19872 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1160_
timestamp 1649977179
transform 1 0 20148 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1161_
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1162_
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1163_
timestamp 1649977179
transform -1 0 16376 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1164_
timestamp 1649977179
transform 1 0 12972 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1649977179
transform -1 0 14536 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1166_
timestamp 1649977179
transform 1 0 14260 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1649977179
transform -1 0 19688 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1168_
timestamp 1649977179
transform 1 0 28060 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1169_
timestamp 1649977179
transform 1 0 18768 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1170_
timestamp 1649977179
transform 1 0 17572 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1171_
timestamp 1649977179
transform 1 0 18032 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1172_
timestamp 1649977179
transform 1 0 25576 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1173_
timestamp 1649977179
transform 1 0 23000 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1174_
timestamp 1649977179
transform 1 0 28612 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1175_
timestamp 1649977179
transform -1 0 30268 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1176_
timestamp 1649977179
transform 1 0 29900 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1177_
timestamp 1649977179
transform -1 0 31372 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1178_
timestamp 1649977179
transform 1 0 27784 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1179_
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1180_
timestamp 1649977179
transform 1 0 27876 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1181_
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1182_
timestamp 1649977179
transform 1 0 27600 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1183_
timestamp 1649977179
transform 1 0 25852 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1184_
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1185_
timestamp 1649977179
transform 1 0 20700 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1186_
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1187_
timestamp 1649977179
transform -1 0 22264 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1188_
timestamp 1649977179
transform 1 0 20700 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _1189_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1190_
timestamp 1649977179
transform -1 0 23460 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1191_
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1192_
timestamp 1649977179
transform -1 0 34684 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1193_
timestamp 1649977179
transform 1 0 39836 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1194_
timestamp 1649977179
transform 1 0 35788 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1195_
timestamp 1649977179
transform -1 0 38640 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1196_
timestamp 1649977179
transform -1 0 36892 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1197_
timestamp 1649977179
transform 1 0 35328 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1198_
timestamp 1649977179
transform 1 0 38640 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1199_
timestamp 1649977179
transform 1 0 35236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1200_
timestamp 1649977179
transform 1 0 38364 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1201_
timestamp 1649977179
transform -1 0 37720 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1202_
timestamp 1649977179
transform -1 0 37352 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1203_
timestamp 1649977179
transform 1 0 37536 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1204_
timestamp 1649977179
transform 1 0 38916 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1205_
timestamp 1649977179
transform 1 0 40388 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1206_
timestamp 1649977179
transform 1 0 38640 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1207_
timestamp 1649977179
transform -1 0 40572 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1208_
timestamp 1649977179
transform -1 0 39560 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1649977179
transform -1 0 37720 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1210_
timestamp 1649977179
transform 1 0 36064 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1211_
timestamp 1649977179
transform 1 0 40020 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1212_
timestamp 1649977179
transform 1 0 33304 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1213_
timestamp 1649977179
transform -1 0 40756 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1214_
timestamp 1649977179
transform 1 0 39928 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1215_
timestamp 1649977179
transform 1 0 40848 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1216_
timestamp 1649977179
transform 1 0 40572 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1217_
timestamp 1649977179
transform 1 0 40112 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1218_
timestamp 1649977179
transform 1 0 40204 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1219_
timestamp 1649977179
transform 1 0 41492 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1220_
timestamp 1649977179
transform 1 0 40388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1221_
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1222_
timestamp 1649977179
transform -1 0 41860 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 1649977179
transform -1 0 36800 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1224_
timestamp 1649977179
transform -1 0 35972 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1225_
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1226_
timestamp 1649977179
transform -1 0 22816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1227_
timestamp 1649977179
transform -1 0 35420 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1228_
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1229_
timestamp 1649977179
transform -1 0 38640 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1230_
timestamp 1649977179
transform 1 0 35972 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1231_
timestamp 1649977179
transform 1 0 37444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1232_
timestamp 1649977179
transform -1 0 35696 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1233_
timestamp 1649977179
transform 1 0 34868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1234_
timestamp 1649977179
transform -1 0 34224 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1235_
timestamp 1649977179
transform 1 0 34868 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1236_
timestamp 1649977179
transform -1 0 36524 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1237_
timestamp 1649977179
transform 1 0 34960 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1238_
timestamp 1649977179
transform 1 0 37076 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1239_
timestamp 1649977179
transform -1 0 38088 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1649977179
transform 1 0 37352 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1241_
timestamp 1649977179
transform 1 0 39100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1242_
timestamp 1649977179
transform -1 0 38916 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1243_
timestamp 1649977179
transform 1 0 37720 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1244_
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1245_
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1246_
timestamp 1649977179
transform 1 0 37536 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1247_
timestamp 1649977179
transform 1 0 38916 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1248_
timestamp 1649977179
transform -1 0 41124 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1249_
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1250_
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1251_
timestamp 1649977179
transform 1 0 39468 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1252_
timestamp 1649977179
transform 1 0 39836 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1253_
timestamp 1649977179
transform 1 0 40020 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1254_
timestamp 1649977179
transform 1 0 40664 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1255_
timestamp 1649977179
transform 1 0 40572 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1256_
timestamp 1649977179
transform 1 0 37352 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1257_
timestamp 1649977179
transform -1 0 38916 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1258_
timestamp 1649977179
transform -1 0 37720 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1259_
timestamp 1649977179
transform -1 0 36340 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1260_
timestamp 1649977179
transform -1 0 23368 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1261_
timestamp 1649977179
transform 1 0 23000 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1262_
timestamp 1649977179
transform -1 0 27232 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1263_
timestamp 1649977179
transform -1 0 30820 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1264_
timestamp 1649977179
transform -1 0 27600 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1265_
timestamp 1649977179
transform 1 0 31188 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1266_
timestamp 1649977179
transform -1 0 27784 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1267_
timestamp 1649977179
transform 1 0 27232 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1268_
timestamp 1649977179
transform -1 0 28796 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1269_
timestamp 1649977179
transform 1 0 27232 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1270_
timestamp 1649977179
transform 1 0 29348 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1271_
timestamp 1649977179
transform -1 0 33856 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1272_
timestamp 1649977179
transform -1 0 30360 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1273_
timestamp 1649977179
transform 1 0 29072 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1274_
timestamp 1649977179
transform 1 0 29900 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1275_
timestamp 1649977179
transform 1 0 29808 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1276_
timestamp 1649977179
transform 1 0 31372 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1277_
timestamp 1649977179
transform 1 0 30728 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1278_
timestamp 1649977179
transform -1 0 30820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 1649977179
transform -1 0 33488 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1280_
timestamp 1649977179
transform -1 0 33212 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1281_
timestamp 1649977179
transform 1 0 33856 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1282_
timestamp 1649977179
transform -1 0 33488 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1649977179
transform 1 0 31832 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1284_
timestamp 1649977179
transform 1 0 14168 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1285_
timestamp 1649977179
transform 1 0 24748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1286_
timestamp 1649977179
transform -1 0 33304 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1287_
timestamp 1649977179
transform 1 0 32660 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1288_
timestamp 1649977179
transform -1 0 33120 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1289_
timestamp 1649977179
transform 1 0 32200 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1290_
timestamp 1649977179
transform -1 0 33028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1291_
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1292_
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1293_
timestamp 1649977179
transform -1 0 26312 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1294_
timestamp 1649977179
transform 1 0 25668 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1295_
timestamp 1649977179
transform 1 0 4968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1296_
timestamp 1649977179
transform 1 0 20976 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1297_
timestamp 1649977179
transform -1 0 16744 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1298_
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _1299_
timestamp 1649977179
transform -1 0 13248 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1300_
timestamp 1649977179
transform -1 0 7728 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1649977179
transform -1 0 16560 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1649977179
transform 1 0 8464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1303_
timestamp 1649977179
transform -1 0 4692 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1304_
timestamp 1649977179
transform -1 0 7636 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1305_
timestamp 1649977179
transform 1 0 3680 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1306_
timestamp 1649977179
transform 1 0 5336 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1307_
timestamp 1649977179
transform -1 0 2024 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1308_
timestamp 1649977179
transform 1 0 2300 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1309_
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1649977179
transform 1 0 2208 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1311_
timestamp 1649977179
transform 1 0 2024 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1312_
timestamp 1649977179
transform 1 0 8096 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1313_
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1314_
timestamp 1649977179
transform -1 0 8004 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1315_
timestamp 1649977179
transform 1 0 6072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1316_
timestamp 1649977179
transform 1 0 5428 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1317_
timestamp 1649977179
transform -1 0 6900 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1318_
timestamp 1649977179
transform 1 0 21344 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1319_
timestamp 1649977179
transform 1 0 19872 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1320_
timestamp 1649977179
transform 1 0 20240 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1321_
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1322_
timestamp 1649977179
transform -1 0 22724 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1323_
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1324_
timestamp 1649977179
transform -1 0 25944 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1325_
timestamp 1649977179
transform -1 0 23368 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1326_
timestamp 1649977179
transform -1 0 23644 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1327_
timestamp 1649977179
transform -1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1328_
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1329_
timestamp 1649977179
transform -1 0 23552 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1330_
timestamp 1649977179
transform 1 0 15272 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1331_
timestamp 1649977179
transform 1 0 22080 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1332_
timestamp 1649977179
transform 1 0 21988 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1333_
timestamp 1649977179
transform 1 0 16100 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1649977179
transform -1 0 23000 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1335_
timestamp 1649977179
transform 1 0 21528 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1336_
timestamp 1649977179
transform 1 0 12052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1649977179
transform 1 0 18308 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1338_
timestamp 1649977179
transform -1 0 20976 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1339_
timestamp 1649977179
transform 1 0 18032 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1340_
timestamp 1649977179
transform 1 0 9476 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1341_
timestamp 1649977179
transform 1 0 20608 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1342_
timestamp 1649977179
transform 1 0 19504 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_4  _1343_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1649977179
transform 1 0 22448 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1345_
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1346_
timestamp 1649977179
transform -1 0 21988 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1347_
timestamp 1649977179
transform -1 0 21988 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1348_
timestamp 1649977179
transform -1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1349_
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1350_
timestamp 1649977179
transform 1 0 20240 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1351_
timestamp 1649977179
transform -1 0 17940 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1352_
timestamp 1649977179
transform -1 0 17296 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1353_
timestamp 1649977179
transform -1 0 19504 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 1649977179
transform -1 0 18768 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1355_
timestamp 1649977179
transform -1 0 17112 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1356_
timestamp 1649977179
transform 1 0 15456 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1357_
timestamp 1649977179
transform -1 0 17572 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1358_
timestamp 1649977179
transform 1 0 16652 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1359_
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1360_
timestamp 1649977179
transform -1 0 19044 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1361_
timestamp 1649977179
transform -1 0 18400 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1362_
timestamp 1649977179
transform 1 0 23828 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1363_
timestamp 1649977179
transform -1 0 25392 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1364_
timestamp 1649977179
transform -1 0 25024 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1365_
timestamp 1649977179
transform -1 0 25576 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 1649977179
transform -1 0 26036 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1367_
timestamp 1649977179
transform -1 0 25392 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1368_
timestamp 1649977179
transform 1 0 26864 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1369_
timestamp 1649977179
transform -1 0 26496 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1370_
timestamp 1649977179
transform -1 0 26220 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1371_
timestamp 1649977179
transform -1 0 12972 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1372_
timestamp 1649977179
transform -1 0 10856 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1373_
timestamp 1649977179
transform -1 0 25760 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1374_
timestamp 1649977179
transform -1 0 26404 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1375_
timestamp 1649977179
transform -1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1376_
timestamp 1649977179
transform 1 0 21896 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1377_
timestamp 1649977179
transform 1 0 23000 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1378_
timestamp 1649977179
transform -1 0 24840 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1379_
timestamp 1649977179
transform -1 0 23460 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1380_
timestamp 1649977179
transform -1 0 10396 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1381_
timestamp 1649977179
transform 1 0 10120 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1382_
timestamp 1649977179
transform -1 0 9660 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1383_
timestamp 1649977179
transform -1 0 8280 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1384_
timestamp 1649977179
transform 1 0 11224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1385_
timestamp 1649977179
transform -1 0 12236 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1386_
timestamp 1649977179
transform -1 0 9844 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1387_
timestamp 1649977179
transform 1 0 7360 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1388_
timestamp 1649977179
transform 1 0 8188 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1389_
timestamp 1649977179
transform -1 0 4232 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1390_
timestamp 1649977179
transform 1 0 10488 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1391_
timestamp 1649977179
transform 1 0 2576 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1649977179
transform -1 0 4140 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1393_
timestamp 1649977179
transform 1 0 2576 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1394_
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1395_
timestamp 1649977179
transform -1 0 7084 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1396_
timestamp 1649977179
transform -1 0 8372 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1397_
timestamp 1649977179
transform 1 0 6808 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1398_
timestamp 1649977179
transform 1 0 14812 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1399_
timestamp 1649977179
transform 1 0 14536 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1400_
timestamp 1649977179
transform -1 0 15640 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1401_
timestamp 1649977179
transform -1 0 14812 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1402_
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1403_
timestamp 1649977179
transform 1 0 11960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1404_
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1405_
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1406_
timestamp 1649977179
transform -1 0 18492 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1407_
timestamp 1649977179
transform -1 0 18308 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1408_
timestamp 1649977179
transform 1 0 17480 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1409_
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1410_
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1411_
timestamp 1649977179
transform 1 0 14904 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1412_
timestamp 1649977179
transform -1 0 14536 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1413_
timestamp 1649977179
transform -1 0 11960 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1414_
timestamp 1649977179
transform -1 0 9936 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1415_
timestamp 1649977179
transform -1 0 11040 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1416_
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1417_
timestamp 1649977179
transform -1 0 11040 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1418_
timestamp 1649977179
transform 1 0 8280 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1419_
timestamp 1649977179
transform -1 0 9660 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1420_
timestamp 1649977179
transform -1 0 9568 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1421_
timestamp 1649977179
transform -1 0 9108 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 1649977179
transform -1 0 4692 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1423_
timestamp 1649977179
transform 1 0 2760 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1424_
timestamp 1649977179
transform -1 0 2852 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1425_
timestamp 1649977179
transform 1 0 2116 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1426_
timestamp 1649977179
transform -1 0 2852 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1427_
timestamp 1649977179
transform 1 0 2024 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1428_
timestamp 1649977179
transform 1 0 4416 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1429_
timestamp 1649977179
transform 1 0 4324 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1430_
timestamp 1649977179
transform -1 0 8096 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1431_
timestamp 1649977179
transform 1 0 9936 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1432_
timestamp 1649977179
transform 1 0 6992 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1433_
timestamp 1649977179
transform 1 0 9476 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1434_
timestamp 1649977179
transform -1 0 9568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1435_
timestamp 1649977179
transform 1 0 9200 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1436_
timestamp 1649977179
transform 1 0 9568 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1437_
timestamp 1649977179
transform -1 0 11592 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1438_
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1440_
timestamp 1649977179
transform -1 0 12236 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1441_
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1442_
timestamp 1649977179
transform -1 0 11500 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1443_
timestamp 1649977179
transform 1 0 10580 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1444_
timestamp 1649977179
transform 1 0 11960 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1445_
timestamp 1649977179
transform -1 0 11960 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1446_
timestamp 1649977179
transform 1 0 10304 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1447_
timestamp 1649977179
transform 1 0 10212 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1448_
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1449_
timestamp 1649977179
transform 1 0 8924 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1450_
timestamp 1649977179
transform 1 0 9016 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1451_
timestamp 1649977179
transform -1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1452_
timestamp 1649977179
transform 1 0 14260 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1453_
timestamp 1649977179
transform -1 0 14444 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1454_
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1455_
timestamp 1649977179
transform 1 0 14904 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1456_
timestamp 1649977179
transform -1 0 16008 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1457_
timestamp 1649977179
transform -1 0 15548 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1458_
timestamp 1649977179
transform -1 0 12512 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1459_
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1460_
timestamp 1649977179
transform -1 0 11960 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1461_
timestamp 1649977179
transform 1 0 11224 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1462_
timestamp 1649977179
transform 1 0 11868 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1463_
timestamp 1649977179
transform 1 0 14444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1464_
timestamp 1649977179
transform 1 0 11868 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1465_
timestamp 1649977179
transform 1 0 13156 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1466_
timestamp 1649977179
transform -1 0 14168 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1467_
timestamp 1649977179
transform 1 0 12972 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1468_
timestamp 1649977179
transform 1 0 12696 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1469_
timestamp 1649977179
transform -1 0 18492 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1470_
timestamp 1649977179
transform -1 0 18308 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1471_
timestamp 1649977179
transform -1 0 19688 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1472_
timestamp 1649977179
transform -1 0 18768 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1473_
timestamp 1649977179
transform -1 0 19228 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1474_
timestamp 1649977179
transform -1 0 18768 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1475_
timestamp 1649977179
transform 1 0 20884 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1476_
timestamp 1649977179
transform -1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1477_
timestamp 1649977179
transform -1 0 22540 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1478_
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1479_
timestamp 1649977179
transform -1 0 22540 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1480_
timestamp 1649977179
transform -1 0 20056 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1481_
timestamp 1649977179
transform 1 0 17664 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp 1649977179
transform -1 0 18032 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1483_
timestamp 1649977179
transform 1 0 16928 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1484_
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1485_
timestamp 1649977179
transform -1 0 18768 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _1486_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7636 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1487_
timestamp 1649977179
transform 1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1488_
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1489_
timestamp 1649977179
transform -1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1490_
timestamp 1649977179
transform 1 0 17848 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1491_
timestamp 1649977179
transform 1 0 20884 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1492_
timestamp 1649977179
transform 1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1493_
timestamp 1649977179
transform -1 0 17112 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1494_
timestamp 1649977179
transform 1 0 16008 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1495_
timestamp 1649977179
transform -1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1496_
timestamp 1649977179
transform -1 0 16652 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1497_
timestamp 1649977179
transform -1 0 15824 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1498_
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1499_
timestamp 1649977179
transform 1 0 14168 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1500_
timestamp 1649977179
transform -1 0 19504 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1501_
timestamp 1649977179
transform -1 0 18768 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1502_
timestamp 1649977179
transform 1 0 19504 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1503_
timestamp 1649977179
transform -1 0 18492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1504_
timestamp 1649977179
transform 1 0 25944 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1505_
timestamp 1649977179
transform -1 0 27232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1506_
timestamp 1649977179
transform -1 0 30636 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1507_
timestamp 1649977179
transform 1 0 25576 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1508_
timestamp 1649977179
transform -1 0 30268 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1509_
timestamp 1649977179
transform 1 0 31096 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1510_
timestamp 1649977179
transform -1 0 30728 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1511_
timestamp 1649977179
transform -1 0 31096 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1512_
timestamp 1649977179
transform -1 0 30820 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1513_
timestamp 1649977179
transform -1 0 28244 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1514_
timestamp 1649977179
transform 1 0 26864 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1515_
timestamp 1649977179
transform -1 0 28796 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1516_
timestamp 1649977179
transform 1 0 27232 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1517_
timestamp 1649977179
transform -1 0 18768 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1518_
timestamp 1649977179
transform 1 0 11868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1519_
timestamp 1649977179
transform 1 0 17296 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1520_
timestamp 1649977179
transform -1 0 19964 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1521_
timestamp 1649977179
transform -1 0 19136 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1522_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9200 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1523_
timestamp 1649977179
transform -1 0 7912 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1524_
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1525_
timestamp 1649977179
transform -1 0 5888 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1526_
timestamp 1649977179
transform 1 0 5152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1527_
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _1528_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4b_2  _1529_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1530_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5060 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1531_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35880 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1532_
timestamp 1649977179
transform 1 0 22816 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1533_
timestamp 1649977179
transform 1 0 22448 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1534_
timestamp 1649977179
transform -1 0 30176 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1535_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 24932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1536_
timestamp 1649977179
transform 1 0 5244 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1537_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6624 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1538_
timestamp 1649977179
transform 1 0 9844 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1539_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1540_
timestamp 1649977179
transform -1 0 9568 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1541_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1542_
timestamp 1649977179
transform -1 0 35696 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1649977179
transform 1 0 22540 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1544_
timestamp 1649977179
transform 1 0 23092 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1545_
timestamp 1649977179
transform -1 0 30176 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1546_
timestamp 1649977179
transform -1 0 24196 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 1649977179
transform 1 0 4232 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1548_
timestamp 1649977179
transform 1 0 4968 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1549_
timestamp 1649977179
transform 1 0 9844 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1550_
timestamp 1649977179
transform -1 0 10672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1551_
timestamp 1649977179
transform -1 0 7820 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1552_
timestamp 1649977179
transform 1 0 6164 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1553_
timestamp 1649977179
transform -1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1554_
timestamp 1649977179
transform 1 0 6348 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1555_
timestamp 1649977179
transform -1 0 35696 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1556_
timestamp 1649977179
transform 1 0 21804 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1557_
timestamp 1649977179
transform 1 0 22080 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1558_
timestamp 1649977179
transform -1 0 28980 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1559_
timestamp 1649977179
transform -1 0 25116 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1560_
timestamp 1649977179
transform 1 0 4140 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1561_
timestamp 1649977179
transform 1 0 4876 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1562_
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1563_
timestamp 1649977179
transform 1 0 12880 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1564_
timestamp 1649977179
transform -1 0 6992 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1565_
timestamp 1649977179
transform 1 0 5152 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1566_
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1567_
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1568_
timestamp 1649977179
transform 1 0 35420 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1569_
timestamp 1649977179
transform 1 0 36248 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1570_
timestamp 1649977179
transform 1 0 35144 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1571_
timestamp 1649977179
transform 1 0 35880 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1572_
timestamp 1649977179
transform -1 0 36708 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1573_
timestamp 1649977179
transform 1 0 23460 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1574_
timestamp 1649977179
transform 1 0 29624 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1575_
timestamp 1649977179
transform -1 0 23092 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1576_
timestamp 1649977179
transform 1 0 29440 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1577_
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1578_
timestamp 1649977179
transform 1 0 21896 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1579_
timestamp 1649977179
transform 1 0 28244 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1580_
timestamp 1649977179
transform 1 0 21620 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1581_
timestamp 1649977179
transform 1 0 28152 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1649977179
transform 1 0 27140 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1583_
timestamp 1649977179
transform 1 0 31096 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1584_
timestamp 1649977179
transform -1 0 33856 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1585_
timestamp 1649977179
transform -1 0 31648 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1586_
timestamp 1649977179
transform -1 0 33856 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1587_
timestamp 1649977179
transform -1 0 31464 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1588_
timestamp 1649977179
transform -1 0 31096 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1589_
timestamp 1649977179
transform 1 0 12880 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1590_
timestamp 1649977179
transform -1 0 13616 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1591_
timestamp 1649977179
transform 1 0 11592 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1592_
timestamp 1649977179
transform -1 0 13432 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1593_
timestamp 1649977179
transform 1 0 6624 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1594_
timestamp 1649977179
transform 1 0 6808 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1595_
timestamp 1649977179
transform 1 0 19412 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1596_
timestamp 1649977179
transform 1 0 22172 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1597_
timestamp 1649977179
transform 1 0 18032 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1598_
timestamp 1649977179
transform 1 0 22448 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1599_
timestamp 1649977179
transform -1 0 14720 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1600_
timestamp 1649977179
transform -1 0 14536 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1601_
timestamp 1649977179
transform -1 0 8280 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1602_
timestamp 1649977179
transform 1 0 4784 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1603_
timestamp 1649977179
transform 1 0 7544 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _1604_
timestamp 1649977179
transform -1 0 7728 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1605_
timestamp 1649977179
transform -1 0 36616 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1606_
timestamp 1649977179
transform -1 0 31372 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1608_
timestamp 1649977179
transform -1 0 30820 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1609_
timestamp 1649977179
transform -1 0 30176 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1610_
timestamp 1649977179
transform -1 0 14444 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1611_
timestamp 1649977179
transform -1 0 13064 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1612_
timestamp 1649977179
transform 1 0 7820 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1613_
timestamp 1649977179
transform 1 0 8096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1614_
timestamp 1649977179
transform -1 0 20608 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1615_
timestamp 1649977179
transform -1 0 17204 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1616_
timestamp 1649977179
transform 1 0 14812 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1617_
timestamp 1649977179
transform 1 0 15364 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1618_
timestamp 1649977179
transform -1 0 9108 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1619_
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1620_
timestamp 1649977179
transform 1 0 7268 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1621_
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1622_
timestamp 1649977179
transform -1 0 35696 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1623_
timestamp 1649977179
transform 1 0 31004 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1624_
timestamp 1649977179
transform 1 0 32108 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1649977179
transform -1 0 33948 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1626_
timestamp 1649977179
transform -1 0 33304 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1627_
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1628_
timestamp 1649977179
transform 1 0 18032 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1629_
timestamp 1649977179
transform -1 0 22724 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1630_
timestamp 1649977179
transform -1 0 21528 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1631_
timestamp 1649977179
transform -1 0 20976 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1632_
timestamp 1649977179
transform 1 0 5152 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1633_
timestamp 1649977179
transform -1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1634_
timestamp 1649977179
transform -1 0 36432 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1635_
timestamp 1649977179
transform -1 0 34316 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1636_
timestamp 1649977179
transform 1 0 32292 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1637_
timestamp 1649977179
transform -1 0 34960 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1638_
timestamp 1649977179
transform -1 0 33764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1639_
timestamp 1649977179
transform 1 0 12972 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1640_
timestamp 1649977179
transform 1 0 17112 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1641_
timestamp 1649977179
transform -1 0 23368 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1642_
timestamp 1649977179
transform -1 0 22632 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1643_
timestamp 1649977179
transform -1 0 19688 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1644_
timestamp 1649977179
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1645_
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1646_
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1647_
timestamp 1649977179
transform -1 0 36432 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1648_
timestamp 1649977179
transform 1 0 31924 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1649_
timestamp 1649977179
transform 1 0 33120 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1650_
timestamp 1649977179
transform -1 0 34224 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1651_
timestamp 1649977179
transform -1 0 33488 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1652_
timestamp 1649977179
transform 1 0 13156 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1653_
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1654_
timestamp 1649977179
transform -1 0 23460 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1655_
timestamp 1649977179
transform -1 0 23092 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1656_
timestamp 1649977179
transform -1 0 22264 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1657_
timestamp 1649977179
transform 1 0 4968 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a21bo_1  _1658_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1659_
timestamp 1649977179
transform -1 0 12328 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1660_
timestamp 1649977179
transform -1 0 37904 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1662_
timestamp 1649977179
transform 1 0 28428 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1663_
timestamp 1649977179
transform -1 0 35328 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1664_
timestamp 1649977179
transform -1 0 30084 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1665_
timestamp 1649977179
transform 1 0 13340 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1666_
timestamp 1649977179
transform 1 0 18768 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1667_
timestamp 1649977179
transform 1 0 22172 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1668_
timestamp 1649977179
transform -1 0 23092 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1669_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22632 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1670_
timestamp 1649977179
transform 1 0 4508 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1671_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1672_
timestamp 1649977179
transform -1 0 38180 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1673_
timestamp 1649977179
transform 1 0 28428 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1674_
timestamp 1649977179
transform 1 0 28336 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp 1649977179
transform -1 0 34592 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1676_
timestamp 1649977179
transform -1 0 30728 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1677_
timestamp 1649977179
transform 1 0 12512 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1678_
timestamp 1649977179
transform 1 0 16192 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1679_
timestamp 1649977179
transform -1 0 22816 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1680_
timestamp 1649977179
transform -1 0 19688 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1681_
timestamp 1649977179
transform -1 0 18032 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1682_
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1683_
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1684_
timestamp 1649977179
transform -1 0 37904 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1685_
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1686_
timestamp 1649977179
transform 1 0 22448 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1687_
timestamp 1649977179
transform -1 0 33396 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1688_
timestamp 1649977179
transform -1 0 25300 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1689_
timestamp 1649977179
transform 1 0 12604 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1690_
timestamp 1649977179
transform 1 0 15088 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1691_
timestamp 1649977179
transform 1 0 19228 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1692_
timestamp 1649977179
transform 1 0 19688 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _1693_
timestamp 1649977179
transform -1 0 20148 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1694_
timestamp 1649977179
transform -1 0 4600 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1695_
timestamp 1649977179
transform -1 0 4324 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1696_
timestamp 1649977179
transform -1 0 37352 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1697_
timestamp 1649977179
transform 1 0 25208 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1698_
timestamp 1649977179
transform 1 0 25392 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1699_
timestamp 1649977179
transform -1 0 33028 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1700_
timestamp 1649977179
transform -1 0 27508 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1701_
timestamp 1649977179
transform 1 0 12420 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1702_
timestamp 1649977179
transform 1 0 13524 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1703_
timestamp 1649977179
transform -1 0 21896 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1704_
timestamp 1649977179
transform -1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1705_
timestamp 1649977179
transform -1 0 15272 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1706_
timestamp 1649977179
transform 1 0 7544 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1707_
timestamp 1649977179
transform -1 0 10396 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1708_
timestamp 1649977179
transform -1 0 4968 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1709_
timestamp 1649977179
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1710_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1840 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1649977179
transform 1 0 2760 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1649977179
transform 1 0 2760 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1649977179
transform 1 0 1840 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1649977179
transform 1 0 2024 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1649977179
transform 1 0 2760 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 1649977179
transform 1 0 8832 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1649977179
transform 1 0 2300 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1649977179
transform -1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1649977179
transform 1 0 2116 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 1649977179
transform 1 0 6256 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1722_
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1723_
timestamp 1649977179
transform -1 0 3864 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1724_
timestamp 1649977179
transform 1 0 2392 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1725_
timestamp 1649977179
transform 1 0 5152 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1726_
timestamp 1649977179
transform 1 0 6072 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1727_
timestamp 1649977179
transform 1 0 10120 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1728_
timestamp 1649977179
transform -1 0 18124 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1729_
timestamp 1649977179
transform -1 0 17480 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1730_
timestamp 1649977179
transform -1 0 15456 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1731_
timestamp 1649977179
transform 1 0 11960 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1732_
timestamp 1649977179
transform 1 0 11408 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1733_
timestamp 1649977179
transform 1 0 12144 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1734_
timestamp 1649977179
transform 1 0 30084 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1735_
timestamp 1649977179
transform 1 0 27600 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1736_
timestamp 1649977179
transform 1 0 27600 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1737_
timestamp 1649977179
transform -1 0 32200 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1738_
timestamp 1649977179
transform -1 0 31188 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1739_
timestamp 1649977179
transform 1 0 37536 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1740_
timestamp 1649977179
transform 1 0 37904 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1741_
timestamp 1649977179
transform -1 0 40020 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1742_
timestamp 1649977179
transform -1 0 39376 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1743_
timestamp 1649977179
transform -1 0 38824 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1744_
timestamp 1649977179
transform -1 0 36156 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1745_
timestamp 1649977179
transform 1 0 32936 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1746_
timestamp 1649977179
transform 1 0 27600 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1747_
timestamp 1649977179
transform 1 0 27324 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1748_
timestamp 1649977179
transform 1 0 27140 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1749_
timestamp 1649977179
transform -1 0 32292 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1750_
timestamp 1649977179
transform 1 0 30912 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1751_
timestamp 1649977179
transform 1 0 32660 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1752_
timestamp 1649977179
transform -1 0 36340 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1753_
timestamp 1649977179
transform -1 0 36432 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1754_
timestamp 1649977179
transform 1 0 35052 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1755_
timestamp 1649977179
transform 1 0 34776 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1756_
timestamp 1649977179
transform 1 0 31924 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1649977179
transform 1 0 32292 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1649977179
transform -1 0 7820 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1649977179
transform -1 0 7820 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1649977179
transform -1 0 22080 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1649977179
transform -1 0 19688 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1649977179
transform -1 0 20700 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1649977179
transform -1 0 22172 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1767_
timestamp 1649977179
transform 1 0 19320 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1649977179
transform 1 0 14812 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1649977179
transform -1 0 16192 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1770_
timestamp 1649977179
transform 1 0 8280 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1649977179
transform -1 0 10396 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1649977179
transform 1 0 10948 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1649977179
transform 1 0 12788 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1649977179
transform 1 0 14444 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1649977179
transform 1 0 24196 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1649977179
transform -1 0 27140 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1649977179
transform -1 0 26588 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1649977179
transform -1 0 25576 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1649977179
transform -1 0 27600 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1649977179
transform -1 0 27232 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1649977179
transform -1 0 23920 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1649977179
transform -1 0 25208 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1649977179
transform -1 0 23920 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1649977179
transform 1 0 25300 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1649977179
transform 1 0 25024 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1649977179
transform -1 0 33580 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1788_
timestamp 1649977179
transform -1 0 34224 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1789_
timestamp 1649977179
transform 1 0 31096 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1649977179
transform -1 0 33948 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1649977179
transform -1 0 31004 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1649977179
transform 1 0 21620 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1649977179
transform 1 0 25024 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1649977179
transform -1 0 15548 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1649977179
transform -1 0 14628 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1649977179
transform -1 0 18584 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1649977179
transform -1 0 18400 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1649977179
transform -1 0 30268 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1800_
timestamp 1649977179
transform -1 0 32752 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1649977179
transform -1 0 29992 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1649977179
transform 1 0 27600 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1649977179
transform -1 0 26680 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1649977179
transform -1 0 21344 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1649977179
transform -1 0 23276 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1806_
timestamp 1649977179
transform 1 0 35236 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1649977179
transform 1 0 38272 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1808_
timestamp 1649977179
transform 1 0 37444 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1809_
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1810_
timestamp 1649977179
transform 1 0 38548 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1811_
timestamp 1649977179
transform 1 0 35880 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1649977179
transform -1 0 40112 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1649977179
transform -1 0 40204 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1649977179
transform -1 0 39744 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1649977179
transform 1 0 40296 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1649977179
transform -1 0 40296 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1649977179
transform 1 0 35420 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1649977179
transform 1 0 34868 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1649977179
transform 1 0 34776 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1649977179
transform 1 0 37904 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1649977179
transform 1 0 38456 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1649977179
transform -1 0 37168 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1649977179
transform -1 0 40020 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1649977179
transform -1 0 39376 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1649977179
transform -1 0 40020 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1649977179
transform -1 0 40204 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1649977179
transform 1 0 38824 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1649977179
transform 1 0 35972 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1649977179
transform -1 0 26864 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1649977179
transform -1 0 31004 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1833_
timestamp 1649977179
transform -1 0 31096 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1834_
timestamp 1649977179
transform -1 0 31004 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1835_
timestamp 1649977179
transform 1 0 32844 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1649977179
transform -1 0 36156 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1649977179
transform -1 0 34132 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1649977179
transform -1 0 34960 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1649977179
transform -1 0 34132 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1649977179
transform -1 0 27324 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1649977179
transform 1 0 24840 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1649977179
transform 1 0 2392 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1649977179
transform 1 0 1840 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1649977179
transform -1 0 7820 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1649977179
transform 1 0 6624 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1649977179
transform 1 0 20792 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1649977179
transform 1 0 23828 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1649977179
transform 1 0 21712 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1649977179
transform 1 0 17664 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1649977179
transform 1 0 19504 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1649977179
transform 1 0 16836 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1649977179
transform 1 0 15088 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1858_
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1859_
timestamp 1649977179
transform 1 0 25392 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1860_
timestamp 1649977179
transform 1 0 25024 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1861_
timestamp 1649977179
transform 1 0 27876 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1862_
timestamp 1649977179
transform 1 0 26496 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1863_
timestamp 1649977179
transform 1 0 25576 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1864_
timestamp 1649977179
transform -1 0 23644 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1865_
timestamp 1649977179
transform 1 0 23092 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1866_
timestamp 1649977179
transform -1 0 7820 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1867_
timestamp 1649977179
transform 1 0 2576 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1868_
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1869_
timestamp 1649977179
transform 1 0 6348 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1870_
timestamp 1649977179
transform 1 0 6808 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1871_
timestamp 1649977179
transform 1 0 14076 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1872_
timestamp 1649977179
transform 1 0 15640 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1873_
timestamp 1649977179
transform -1 0 20700 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1874_
timestamp 1649977179
transform 1 0 17296 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1875_
timestamp 1649977179
transform -1 0 17020 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1876_
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1877_
timestamp 1649977179
transform 1 0 10580 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1878_
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1879_
timestamp 1649977179
transform 1 0 2392 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1880_
timestamp 1649977179
transform 1 0 2208 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1881_
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1882_
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1883_
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1884_
timestamp 1649977179
transform 1 0 9292 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1885_
timestamp 1649977179
transform 1 0 9292 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1886_
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1887_
timestamp 1649977179
transform 1 0 9936 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1888_
timestamp 1649977179
transform 1 0 9292 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1889_
timestamp 1649977179
transform 1 0 7820 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1890_
timestamp 1649977179
transform 1 0 10212 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1891_
timestamp 1649977179
transform 1 0 9384 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1892_
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1893_
timestamp 1649977179
transform -1 0 15548 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1894_
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1895_
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1896_
timestamp 1649977179
transform 1 0 18952 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1897_
timestamp 1649977179
transform -1 0 23092 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1898_
timestamp 1649977179
transform -1 0 24104 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1899_
timestamp 1649977179
transform 1 0 17112 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1900_
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1901_
timestamp 1649977179
transform 1 0 18676 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1902_
timestamp 1649977179
transform 1 0 15364 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1903_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1904_
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1905_
timestamp 1649977179
transform 1 0 19412 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1906_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1907_
timestamp 1649977179
transform 1 0 29900 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1908_
timestamp 1649977179
transform 1 0 31004 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1909_
timestamp 1649977179
transform 1 0 31280 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1910_
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1911_
timestamp 1649977179
transform 1 0 27232 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1912_
timestamp 1649977179
transform 1 0 17296 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1913_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1914_
timestamp 1649977179
transform -1 0 5336 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1915_
timestamp 1649977179
transform -1 0 8832 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1916_
timestamp 1649977179
transform -1 0 7820 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1917_
timestamp 1649977179
transform -1 0 8280 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1918_
timestamp 1649977179
transform -1 0 8740 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1919_
timestamp 1649977179
transform -1 0 9200 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1920_
timestamp 1649977179
transform 1 0 9660 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1921_
timestamp 1649977179
transform -1 0 12604 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1922_
timestamp 1649977179
transform 1 0 9384 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1923_
timestamp 1649977179
transform 1 0 12052 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1924_
timestamp 1649977179
transform 1 0 2392 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1925_
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1926_
timestamp 1649977179
transform 1 0 1840 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _2167_
timestamp 1649977179
transform -1 0 45816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2168_
timestamp 1649977179
transform -1 0 25852 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2169_
timestamp 1649977179
transform -1 0 45172 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2170_
timestamp 1649977179
transform 1 0 18492 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2171_
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2172_
timestamp 1649977179
transform 1 0 17848 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2173_
timestamp 1649977179
transform 1 0 18308 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2174_
timestamp 1649977179
transform 1 0 20424 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2175_
timestamp 1649977179
transform 1 0 19780 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2176_
timestamp 1649977179
transform -1 0 25208 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2177_
timestamp 1649977179
transform -1 0 34224 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2178_
timestamp 1649977179
transform -1 0 32384 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2179_
timestamp 1649977179
transform -1 0 29900 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2180_
timestamp 1649977179
transform -1 0 27416 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2181_
timestamp 1649977179
transform -1 0 26128 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2182_
timestamp 1649977179
transform -1 0 26496 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2183_
timestamp 1649977179
transform -1 0 26496 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2184_
timestamp 1649977179
transform -1 0 24196 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2185_
timestamp 1649977179
transform -1 0 22908 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2186_
timestamp 1649977179
transform -1 0 21344 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2187_
timestamp 1649977179
transform -1 0 19412 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2188_
timestamp 1649977179
transform -1 0 18768 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2189_
timestamp 1649977179
transform -1 0 17480 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2190_
timestamp 1649977179
transform 1 0 16836 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2191_
timestamp 1649977179
transform 1 0 15916 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2192_
timestamp 1649977179
transform 1 0 13524 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2193_
timestamp 1649977179
transform 1 0 19688 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2194_
timestamp 1649977179
transform -1 0 22264 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2195_
timestamp 1649977179
transform -1 0 31648 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2196_
timestamp 1649977179
transform -1 0 36064 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20792 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1649977179
transform -1 0 9660 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1649977179
transform 1 0 10396 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1649977179
transform 1 0 28612 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1649977179
transform 1 0 28612 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_wb_clk_i
timestamp 1649977179
transform -1 0 17204 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_wb_clk_i
timestamp 1649977179
transform 1 0 10304 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_wb_clk_i
timestamp 1649977179
transform -1 0 5980 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_wb_clk_i
timestamp 1649977179
transform 1 0 5704 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_wb_clk_i
timestamp 1649977179
transform -1 0 5980 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_wb_clk_i
timestamp 1649977179
transform 1 0 9016 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_wb_clk_i
timestamp 1649977179
transform 1 0 11776 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_wb_clk_i
timestamp 1649977179
transform -1 0 20148 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_wb_clk_i
timestamp 1649977179
transform 1 0 17112 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_wb_clk_i
timestamp 1649977179
transform 1 0 20792 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_wb_clk_i
timestamp 1649977179
transform -1 0 28796 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_wb_clk_i
timestamp 1649977179
transform -1 0 25668 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_wb_clk_i
timestamp 1649977179
transform 1 0 27876 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_wb_clk_i
timestamp 1649977179
transform 1 0 32384 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_wb_clk_i
timestamp 1649977179
transform 1 0 34960 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_wb_clk_i
timestamp 1649977179
transform 1 0 39100 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_wb_clk_i
timestamp 1649977179
transform 1 0 33948 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_wb_clk_i
timestamp 1649977179
transform 1 0 27692 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_wb_clk_i
timestamp 1649977179
transform -1 0 27508 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_wb_clk_i
timestamp 1649977179
transform -1 0 34316 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_wb_clk_i
timestamp 1649977179
transform 1 0 38088 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_wb_clk_i
timestamp 1649977179
transform 1 0 37168 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_wb_clk_i
timestamp 1649977179
transform 1 0 37076 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_wb_clk_i
timestamp 1649977179
transform 1 0 34132 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_wb_clk_i
timestamp 1649977179
transform 1 0 29900 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_wb_clk_i
timestamp 1649977179
transform 1 0 24656 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_wb_clk_i
timestamp 1649977179
transform 1 0 24472 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_wb_clk_i
timestamp 1649977179
transform -1 0 24012 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_28_wb_clk_i
timestamp 1649977179
transform 1 0 15824 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_29_wb_clk_i
timestamp 1649977179
transform 1 0 17296 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_30_wb_clk_i
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_31_wb_clk_i
timestamp 1649977179
transform 1 0 3220 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_32_wb_clk_i
timestamp 1649977179
transform 1 0 5888 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_33_wb_clk_i
timestamp 1649977179
transform -1 0 4416 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_34_wb_clk_i
timestamp 1649977179
transform 1 0 9200 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1649977179
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1649977179
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1649977179
transform -1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1649977179
transform -1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1649977179
transform -1 0 19136 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1649977179
transform -1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1649977179
transform -1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1649977179
transform 1 0 20056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1649977179
transform -1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1649977179
transform -1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1649977179
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1649977179
transform -1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1649977179
transform -1 0 20608 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1649977179
transform -1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform -1 0 22080 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1649977179
transform -1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 22080 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1649977179
transform -1 0 22264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input20
timestamp 1649977179
transform 1 0 22816 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1649977179
transform -1 0 23000 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1649977179
transform 1 0 23368 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input24
timestamp 1649977179
transform 1 0 13248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1649977179
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1649977179
transform -1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1649977179
transform 1 0 16836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input28
timestamp 1649977179
transform -1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1649977179
transform 1 0 17572 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1649977179
transform -1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 13616 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform -1 0 8188 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 3680 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform -1 0 1840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1649977179
transform 1 0 6256 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input46
timestamp 1649977179
transform 1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1649977179
transform 1 0 10304 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform 1 0 6992 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input50
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input51
timestamp 1649977179
transform 1 0 8280 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input52
timestamp 1649977179
transform -1 0 6900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input53
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input54
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input55
timestamp 1649977179
transform 1 0 9476 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform -1 0 4140 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform -1 0 4600 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform -1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 47564 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 40940 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 45632 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 10028 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 8464 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 6900 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform -1 0 5336 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 4140 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 2208 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 37812 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 36248 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 34684 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 33120 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 32108 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 29992 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform 1 0 28428 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 26956 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 25300 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 24380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 22172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 20608 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 19228 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 17480 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 17020 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 14720 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 13156 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 11868 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 42504 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 44068 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 39836 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 12236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 6256 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 5152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 10672 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 11868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_103 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 58236 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_104
timestamp 1649977179
transform -1 0 56856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_105
timestamp 1649977179
transform -1 0 55568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_106
timestamp 1649977179
transform -1 0 53728 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_107
timestamp 1649977179
transform -1 0 52164 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_108
timestamp 1649977179
transform -1 0 49036 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_109
timestamp 1649977179
transform -1 0 50600 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_110
timestamp 1649977179
transform 1 0 57960 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_111
timestamp 1649977179
transform 1 0 57960 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_112
timestamp 1649977179
transform 1 0 57316 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_113
timestamp 1649977179
transform 1 0 57960 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_114
timestamp 1649977179
transform -1 0 52992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_115
timestamp 1649977179
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_116
timestamp 1649977179
transform -1 0 51428 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_117
timestamp 1649977179
transform -1 0 52440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_118
timestamp 1649977179
transform -1 0 54280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_119
timestamp 1649977179
transform -1 0 52072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_120
timestamp 1649977179
transform -1 0 53084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_121
timestamp 1649977179
transform -1 0 53636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_122
timestamp 1649977179
transform -1 0 53728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_123
timestamp 1649977179
transform -1 0 54280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_124
timestamp 1649977179
transform -1 0 52992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_125
timestamp 1649977179
transform -1 0 54924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_126
timestamp 1649977179
transform -1 0 55568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_127
timestamp 1649977179
transform -1 0 52440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_128
timestamp 1649977179
transform -1 0 53084 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_129
timestamp 1649977179
transform -1 0 54372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_130
timestamp 1649977179
transform -1 0 56212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_131
timestamp 1649977179
transform -1 0 53636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_132
timestamp 1649977179
transform -1 0 55568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_133
timestamp 1649977179
transform -1 0 53728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_134
timestamp 1649977179
transform -1 0 54280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_135
timestamp 1649977179
transform -1 0 54924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_136
timestamp 1649977179
transform -1 0 56856 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_137
timestamp 1649977179
transform -1 0 55568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_138
timestamp 1649977179
transform -1 0 56212 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_139
timestamp 1649977179
transform -1 0 54372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_140
timestamp 1649977179
transform -1 0 56212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_141
timestamp 1649977179
transform -1 0 56856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_142
timestamp 1649977179
transform -1 0 55568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_143
timestamp 1649977179
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_144
timestamp 1649977179
transform -1 0 54004 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_145
timestamp 1649977179
transform -1 0 54648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_146
timestamp 1649977179
transform -1 0 56856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_147
timestamp 1649977179
transform -1 0 55568 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_148
timestamp 1649977179
transform -1 0 56212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_149
timestamp 1649977179
transform -1 0 55292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_150
timestamp 1649977179
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_151
timestamp 1649977179
transform -1 0 56212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_152
timestamp 1649977179
transform 1 0 57960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_153
timestamp 1649977179
transform 1 0 57316 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_154
timestamp 1649977179
transform 1 0 57960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_155
timestamp 1649977179
transform 1 0 57960 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_156
timestamp 1649977179
transform 1 0 57960 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_157
timestamp 1649977179
transform 1 0 57960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_158
timestamp 1649977179
transform 1 0 57960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_159
timestamp 1649977179
transform 1 0 57960 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_160
timestamp 1649977179
transform 1 0 57960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_161
timestamp 1649977179
transform 1 0 57960 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_162
timestamp 1649977179
transform 1 0 57960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_163
timestamp 1649977179
transform 1 0 57960 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_164
timestamp 1649977179
transform 1 0 57960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_165
timestamp 1649977179
transform 1 0 57960 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_166
timestamp 1649977179
transform 1 0 57960 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_167
timestamp 1649977179
transform 1 0 57960 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_168
timestamp 1649977179
transform 1 0 57960 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_169
timestamp 1649977179
transform 1 0 57960 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_170
timestamp 1649977179
transform 1 0 57960 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_171
timestamp 1649977179
transform 1 0 57960 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_172
timestamp 1649977179
transform 1 0 57960 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_173
timestamp 1649977179
transform 1 0 57960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_174
timestamp 1649977179
transform 1 0 57960 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_175
timestamp 1649977179
transform 1 0 57960 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_176
timestamp 1649977179
transform 1 0 57960 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_177
timestamp 1649977179
transform 1 0 57960 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_178
timestamp 1649977179
transform 1 0 57960 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_179
timestamp 1649977179
transform 1 0 57960 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_180
timestamp 1649977179
transform 1 0 57960 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_181
timestamp 1649977179
transform 1 0 57960 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_182
timestamp 1649977179
transform 1 0 57960 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_183
timestamp 1649977179
transform 1 0 57960 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_184
timestamp 1649977179
transform 1 0 57960 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_185
timestamp 1649977179
transform 1 0 57960 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_186
timestamp 1649977179
transform 1 0 57960 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_187
timestamp 1649977179
transform 1 0 57960 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_188
timestamp 1649977179
transform 1 0 57960 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_189
timestamp 1649977179
transform 1 0 57960 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_190
timestamp 1649977179
transform -1 0 51704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_191
timestamp 1649977179
transform -1 0 51796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_192
timestamp 1649977179
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_193
timestamp 1649977179
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_194
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_195
timestamp 1649977179
transform 1 0 15272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_196
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_197
timestamp 1649977179
transform 1 0 13064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_198
timestamp 1649977179
transform 1 0 15916 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_199
timestamp 1649977179
transform 1 0 15272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_200
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_201
timestamp 1649977179
transform 1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_202
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_203
timestamp 1649977179
transform 1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_204
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_205
timestamp 1649977179
transform 1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_206
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_207
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_208
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_209
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_210
timestamp 1649977179
transform -1 0 20424 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_211
timestamp 1649977179
transform 1 0 18768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_212
timestamp 1649977179
transform 1 0 19872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_213
timestamp 1649977179
transform -1 0 21252 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_214
timestamp 1649977179
transform 1 0 20516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_215
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_216
timestamp 1649977179
transform -1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_217
timestamp 1649977179
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_218
timestamp 1649977179
transform 1 0 21804 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_219
timestamp 1649977179
transform -1 0 22908 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_220
timestamp 1649977179
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_221
timestamp 1649977179
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_222
timestamp 1649977179
transform -1 0 23736 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_223
timestamp 1649977179
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_224
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_225
timestamp 1649977179
transform -1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_226
timestamp 1649977179
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_227
timestamp 1649977179
transform -1 0 24932 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_228
timestamp 1649977179
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_229
timestamp 1649977179
transform -1 0 25668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_230
timestamp 1649977179
transform 1 0 25300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_231
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_232
timestamp 1649977179
transform 1 0 25944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_233
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_234
timestamp 1649977179
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_235
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_236
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_237
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_238
timestamp 1649977179
transform 1 0 27416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_239
timestamp 1649977179
transform -1 0 28336 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_240
timestamp 1649977179
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_241
timestamp 1649977179
transform -1 0 28980 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_242
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_243
timestamp 1649977179
transform 1 0 28704 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_244
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_245
timestamp 1649977179
transform 1 0 29348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_246
timestamp 1649977179
transform -1 0 30268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_247
timestamp 1649977179
transform 1 0 29900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_248
timestamp 1649977179
transform -1 0 30912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_249
timestamp 1649977179
transform 1 0 30544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_250
timestamp 1649977179
transform -1 0 31464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_251
timestamp 1649977179
transform -1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_252
timestamp 1649977179
transform -1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_253
timestamp 1649977179
transform -1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_254
timestamp 1649977179
transform -1 0 33028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_255
timestamp 1649977179
transform -1 0 33672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_256
timestamp 1649977179
transform -1 0 33672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_257
timestamp 1649977179
transform -1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_258
timestamp 1649977179
transform -1 0 34316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_259
timestamp 1649977179
transform -1 0 35604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_260
timestamp 1649977179
transform -1 0 34960 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_261
timestamp 1649977179
transform -1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_262
timestamp 1649977179
transform -1 0 35604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_263
timestamp 1649977179
transform -1 0 35052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_264
timestamp 1649977179
transform -1 0 35696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_265
timestamp 1649977179
transform -1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_266
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_267
timestamp 1649977179
transform -1 0 36340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_268
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_269
timestamp 1649977179
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_270
timestamp 1649977179
transform -1 0 36984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_271
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_272
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_273
timestamp 1649977179
transform -1 0 37812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_274
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_275
timestamp 1649977179
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_276
timestamp 1649977179
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_277
timestamp 1649977179
transform -1 0 38916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_278
timestamp 1649977179
transform -1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_279
timestamp 1649977179
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_280
timestamp 1649977179
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_281
timestamp 1649977179
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_282
timestamp 1649977179
transform -1 0 40296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_283
timestamp 1649977179
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_284
timestamp 1649977179
transform -1 0 40940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_285
timestamp 1649977179
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_286
timestamp 1649977179
transform -1 0 41584 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_287
timestamp 1649977179
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_288
timestamp 1649977179
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_289
timestamp 1649977179
transform -1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_290
timestamp 1649977179
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_291
timestamp 1649977179
transform -1 0 42780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_292
timestamp 1649977179
transform -1 0 43424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_293
timestamp 1649977179
transform -1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_294
timestamp 1649977179
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_295
timestamp 1649977179
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_296
timestamp 1649977179
transform -1 0 45908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_297
timestamp 1649977179
transform -1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_298
timestamp 1649977179
transform -1 0 45264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_299
timestamp 1649977179
transform -1 0 46552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_300
timestamp 1649977179
transform -1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_301
timestamp 1649977179
transform -1 0 45908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_302
timestamp 1649977179
transform -1 0 46552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_303
timestamp 1649977179
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_304
timestamp 1649977179
transform -1 0 46552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_305
timestamp 1649977179
transform -1 0 47196 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_306
timestamp 1649977179
transform -1 0 48484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_307
timestamp 1649977179
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_308
timestamp 1649977179
transform -1 0 49128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_309
timestamp 1649977179
transform -1 0 48484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_310
timestamp 1649977179
transform -1 0 48024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_311
timestamp 1649977179
transform -1 0 49128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_312
timestamp 1649977179
transform -1 0 48668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_313
timestamp 1649977179
transform -1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_314
timestamp 1649977179
transform -1 0 49772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_315
timestamp 1649977179
transform -1 0 51060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_316
timestamp 1649977179
transform -1 0 50416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_317
timestamp 1649977179
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_318
timestamp 1649977179
transform -1 0 51060 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_319
timestamp 1649977179
transform -1 0 50508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_320
timestamp 1649977179
transform -1 0 51152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_321
timestamp 1649977179
transform 1 0 57960 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_322
timestamp 1649977179
transform 1 0 57960 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_323
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_324
timestamp 1649977179
transform 1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_325
timestamp 1649977179
transform -1 0 11040 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_326
timestamp 1649977179
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_327
timestamp 1649977179
transform 1 0 9476 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_328
timestamp 1649977179
transform 1 0 10580 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_329
timestamp 1649977179
transform -1 0 11868 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_330
timestamp 1649977179
transform 1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_331
timestamp 1649977179
transform -1 0 12512 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_332
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_333
timestamp 1649977179
transform -1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_334
timestamp 1649977179
transform -1 0 13340 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_335
timestamp 1649977179
transform -1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_336
timestamp 1649977179
transform 1 0 12696 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_337
timestamp 1649977179
transform 1 0 13524 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_338
timestamp 1649977179
transform -1 0 14444 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_339
timestamp 1649977179
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_340
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_341
timestamp 1649977179
transform 1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_342
timestamp 1649977179
transform 1 0 13984 0 -1 4352
box -38 -48 314 592
<< labels >>
flabel metal2 s 47122 59200 47178 60000 0 FreeSans 224 90 0 0 CMP_out_c
port 0 nsew signal tristate
flabel metal2 s 40866 59200 40922 60000 0 FreeSans 224 90 0 0 OTA_out_c
port 1 nsew signal tristate
flabel metal2 s 45558 59200 45614 60000 0 FreeSans 224 90 0 0 OTA_sh_c
port 2 nsew signal tristate
flabel metal2 s 9586 59200 9642 60000 0 FreeSans 224 90 0 0 Pd10_a
port 3 nsew signal tristate
flabel metal2 s 8022 59200 8078 60000 0 FreeSans 224 90 0 0 Pd10_b
port 4 nsew signal tristate
flabel metal2 s 6458 59200 6514 60000 0 FreeSans 224 90 0 0 Pd11_a
port 5 nsew signal tristate
flabel metal2 s 4894 59200 4950 60000 0 FreeSans 224 90 0 0 Pd11_b
port 6 nsew signal tristate
flabel metal2 s 3330 59200 3386 60000 0 FreeSans 224 90 0 0 Pd12_a
port 7 nsew signal tristate
flabel metal2 s 1766 59200 1822 60000 0 FreeSans 224 90 0 0 Pd12_b
port 8 nsew signal tristate
flabel metal2 s 37738 59200 37794 60000 0 FreeSans 224 90 0 0 Pd1_a
port 9 nsew signal tristate
flabel metal2 s 36174 59200 36230 60000 0 FreeSans 224 90 0 0 Pd1_b
port 10 nsew signal tristate
flabel metal2 s 34610 59200 34666 60000 0 FreeSans 224 90 0 0 Pd2_a
port 11 nsew signal tristate
flabel metal2 s 33046 59200 33102 60000 0 FreeSans 224 90 0 0 Pd2_b
port 12 nsew signal tristate
flabel metal2 s 31482 59200 31538 60000 0 FreeSans 224 90 0 0 Pd3_a
port 13 nsew signal tristate
flabel metal2 s 29918 59200 29974 60000 0 FreeSans 224 90 0 0 Pd3_b
port 14 nsew signal tristate
flabel metal2 s 28354 59200 28410 60000 0 FreeSans 224 90 0 0 Pd4_a
port 15 nsew signal tristate
flabel metal2 s 26790 59200 26846 60000 0 FreeSans 224 90 0 0 Pd4_b
port 16 nsew signal tristate
flabel metal2 s 25226 59200 25282 60000 0 FreeSans 224 90 0 0 Pd5_a
port 17 nsew signal tristate
flabel metal2 s 23662 59200 23718 60000 0 FreeSans 224 90 0 0 Pd5_b
port 18 nsew signal tristate
flabel metal2 s 22098 59200 22154 60000 0 FreeSans 224 90 0 0 Pd6_a
port 19 nsew signal tristate
flabel metal2 s 20534 59200 20590 60000 0 FreeSans 224 90 0 0 Pd6_b
port 20 nsew signal tristate
flabel metal2 s 18970 59200 19026 60000 0 FreeSans 224 90 0 0 Pd7_a
port 21 nsew signal tristate
flabel metal2 s 17406 59200 17462 60000 0 FreeSans 224 90 0 0 Pd7_b
port 22 nsew signal tristate
flabel metal2 s 15842 59200 15898 60000 0 FreeSans 224 90 0 0 Pd8_a
port 23 nsew signal tristate
flabel metal2 s 14278 59200 14334 60000 0 FreeSans 224 90 0 0 Pd8_b
port 24 nsew signal tristate
flabel metal2 s 12714 59200 12770 60000 0 FreeSans 224 90 0 0 Pd9_a
port 25 nsew signal tristate
flabel metal2 s 11150 59200 11206 60000 0 FreeSans 224 90 0 0 Pd9_b
port 26 nsew signal tristate
flabel metal2 s 42430 59200 42486 60000 0 FreeSans 224 90 0 0 SH_out_c
port 27 nsew signal tristate
flabel metal2 s 58070 59200 58126 60000 0 FreeSans 224 90 0 0 Sh
port 28 nsew signal tristate
flabel metal2 s 56506 59200 56562 60000 0 FreeSans 224 90 0 0 Sh_cmp
port 29 nsew signal tristate
flabel metal2 s 54942 59200 54998 60000 0 FreeSans 224 90 0 0 Sh_rst
port 30 nsew signal tristate
flabel metal2 s 53378 59200 53434 60000 0 FreeSans 224 90 0 0 Sw1
port 31 nsew signal tristate
flabel metal2 s 51814 59200 51870 60000 0 FreeSans 224 90 0 0 Sw2
port 32 nsew signal tristate
flabel metal2 s 48686 59200 48742 60000 0 FreeSans 224 90 0 0 Vd1
port 33 nsew signal tristate
flabel metal2 s 50250 59200 50306 60000 0 FreeSans 224 90 0 0 Vd2
port 34 nsew signal tristate
flabel metal2 s 43994 59200 44050 60000 0 FreeSans 224 90 0 0 Vref_cmp_c
port 35 nsew signal tristate
flabel metal2 s 39302 59200 39358 60000 0 FreeSans 224 90 0 0 Vref_sel_c
port 36 nsew signal tristate
flabel metal3 s 59200 52368 60000 52488 0 FreeSans 480 0 0 0 clk_o
port 37 nsew signal tristate
flabel metal3 s 59200 59168 60000 59288 0 FreeSans 480 0 0 0 counter_rst
port 38 nsew signal tristate
flabel metal3 s 59200 57808 60000 57928 0 FreeSans 480 0 0 0 data_o
port 39 nsew signal tristate
flabel metal3 s 59200 55088 60000 55208 0 FreeSans 480 0 0 0 done_o
port 40 nsew signal tristate
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 io_in[0]
port 41 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 io_in[10]
port 42 nsew signal input
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 io_in[11]
port 43 nsew signal input
flabel metal3 s 0 20136 800 20256 0 FreeSans 480 0 0 0 io_in[12]
port 44 nsew signal input
flabel metal3 s 0 21632 800 21752 0 FreeSans 480 0 0 0 io_in[13]
port 45 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 io_in[14]
port 46 nsew signal input
flabel metal3 s 0 24624 800 24744 0 FreeSans 480 0 0 0 io_in[15]
port 47 nsew signal input
flabel metal3 s 0 26120 800 26240 0 FreeSans 480 0 0 0 io_in[16]
port 48 nsew signal input
flabel metal3 s 0 27616 800 27736 0 FreeSans 480 0 0 0 io_in[17]
port 49 nsew signal input
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 io_in[18]
port 50 nsew signal input
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 io_in[19]
port 51 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 io_in[1]
port 52 nsew signal input
flabel metal3 s 0 32104 800 32224 0 FreeSans 480 0 0 0 io_in[20]
port 53 nsew signal input
flabel metal3 s 0 33600 800 33720 0 FreeSans 480 0 0 0 io_in[21]
port 54 nsew signal input
flabel metal3 s 0 35096 800 35216 0 FreeSans 480 0 0 0 io_in[22]
port 55 nsew signal input
flabel metal3 s 0 36592 800 36712 0 FreeSans 480 0 0 0 io_in[23]
port 56 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 io_in[24]
port 57 nsew signal input
flabel metal3 s 0 39584 800 39704 0 FreeSans 480 0 0 0 io_in[25]
port 58 nsew signal input
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 io_in[26]
port 59 nsew signal input
flabel metal3 s 0 42576 800 42696 0 FreeSans 480 0 0 0 io_in[27]
port 60 nsew signal input
flabel metal3 s 0 44072 800 44192 0 FreeSans 480 0 0 0 io_in[28]
port 61 nsew signal input
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 io_in[29]
port 62 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 io_in[2]
port 63 nsew signal input
flabel metal3 s 0 47064 800 47184 0 FreeSans 480 0 0 0 io_in[30]
port 64 nsew signal input
flabel metal3 s 0 48560 800 48680 0 FreeSans 480 0 0 0 io_in[31]
port 65 nsew signal input
flabel metal3 s 0 50056 800 50176 0 FreeSans 480 0 0 0 io_in[32]
port 66 nsew signal input
flabel metal3 s 0 51552 800 51672 0 FreeSans 480 0 0 0 io_in[33]
port 67 nsew signal input
flabel metal3 s 0 53048 800 53168 0 FreeSans 480 0 0 0 io_in[34]
port 68 nsew signal input
flabel metal3 s 0 54544 800 54664 0 FreeSans 480 0 0 0 io_in[35]
port 69 nsew signal input
flabel metal3 s 0 56040 800 56160 0 FreeSans 480 0 0 0 io_in[36]
port 70 nsew signal input
flabel metal3 s 0 57536 800 57656 0 FreeSans 480 0 0 0 io_in[37]
port 71 nsew signal input
flabel metal3 s 0 6672 800 6792 0 FreeSans 480 0 0 0 io_in[3]
port 72 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 io_in[4]
port 73 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 io_in[5]
port 74 nsew signal input
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 io_in[6]
port 75 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 io_in[7]
port 76 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 io_in[8]
port 77 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 io_in[9]
port 78 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 79 nsew signal tristate
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 io_oeb[10]
port 80 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 io_oeb[11]
port 81 nsew signal tristate
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 io_oeb[12]
port 82 nsew signal tristate
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 io_oeb[13]
port 83 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 io_oeb[14]
port 84 nsew signal tristate
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 io_oeb[15]
port 85 nsew signal tristate
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 io_oeb[16]
port 86 nsew signal tristate
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 io_oeb[17]
port 87 nsew signal tristate
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 io_oeb[18]
port 88 nsew signal tristate
flabel metal2 s 52642 0 52698 800 0 FreeSans 224 90 0 0 io_oeb[19]
port 89 nsew signal tristate
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 io_oeb[1]
port 90 nsew signal tristate
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 io_oeb[20]
port 91 nsew signal tristate
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 io_oeb[21]
port 92 nsew signal tristate
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 io_oeb[22]
port 93 nsew signal tristate
flabel metal2 s 53010 0 53066 800 0 FreeSans 224 90 0 0 io_oeb[23]
port 94 nsew signal tristate
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 io_oeb[24]
port 95 nsew signal tristate
flabel metal2 s 53194 0 53250 800 0 FreeSans 224 90 0 0 io_oeb[25]
port 96 nsew signal tristate
flabel metal2 s 53286 0 53342 800 0 FreeSans 224 90 0 0 io_oeb[26]
port 97 nsew signal tristate
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 io_oeb[27]
port 98 nsew signal tristate
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 io_oeb[28]
port 99 nsew signal tristate
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 io_oeb[29]
port 100 nsew signal tristate
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 io_oeb[2]
port 101 nsew signal tristate
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 io_oeb[30]
port 102 nsew signal tristate
flabel metal2 s 53746 0 53802 800 0 FreeSans 224 90 0 0 io_oeb[31]
port 103 nsew signal tristate
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 io_oeb[32]
port 104 nsew signal tristate
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 io_oeb[33]
port 105 nsew signal tristate
flabel metal2 s 54022 0 54078 800 0 FreeSans 224 90 0 0 io_oeb[34]
port 106 nsew signal tristate
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 io_oeb[35]
port 107 nsew signal tristate
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 io_oeb[36]
port 108 nsew signal tristate
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 io_oeb[37]
port 109 nsew signal tristate
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 io_oeb[3]
port 110 nsew signal tristate
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 io_oeb[4]
port 111 nsew signal tristate
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 io_oeb[5]
port 112 nsew signal tristate
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 io_oeb[6]
port 113 nsew signal tristate
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 io_oeb[7]
port 114 nsew signal tristate
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 io_oeb[8]
port 115 nsew signal tristate
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 io_oeb[9]
port 116 nsew signal tristate
flabel metal3 s 59200 688 60000 808 0 FreeSans 480 0 0 0 io_out[0]
port 117 nsew signal tristate
flabel metal3 s 59200 14288 60000 14408 0 FreeSans 480 0 0 0 io_out[10]
port 118 nsew signal tristate
flabel metal3 s 59200 15648 60000 15768 0 FreeSans 480 0 0 0 io_out[11]
port 119 nsew signal tristate
flabel metal3 s 59200 17008 60000 17128 0 FreeSans 480 0 0 0 io_out[12]
port 120 nsew signal tristate
flabel metal3 s 59200 18368 60000 18488 0 FreeSans 480 0 0 0 io_out[13]
port 121 nsew signal tristate
flabel metal3 s 59200 19728 60000 19848 0 FreeSans 480 0 0 0 io_out[14]
port 122 nsew signal tristate
flabel metal3 s 59200 21088 60000 21208 0 FreeSans 480 0 0 0 io_out[15]
port 123 nsew signal tristate
flabel metal3 s 59200 22448 60000 22568 0 FreeSans 480 0 0 0 io_out[16]
port 124 nsew signal tristate
flabel metal3 s 59200 23808 60000 23928 0 FreeSans 480 0 0 0 io_out[17]
port 125 nsew signal tristate
flabel metal3 s 59200 25168 60000 25288 0 FreeSans 480 0 0 0 io_out[18]
port 126 nsew signal tristate
flabel metal3 s 59200 26528 60000 26648 0 FreeSans 480 0 0 0 io_out[19]
port 127 nsew signal tristate
flabel metal3 s 59200 2048 60000 2168 0 FreeSans 480 0 0 0 io_out[1]
port 128 nsew signal tristate
flabel metal3 s 59200 27888 60000 28008 0 FreeSans 480 0 0 0 io_out[20]
port 129 nsew signal tristate
flabel metal3 s 59200 29248 60000 29368 0 FreeSans 480 0 0 0 io_out[21]
port 130 nsew signal tristate
flabel metal3 s 59200 30608 60000 30728 0 FreeSans 480 0 0 0 io_out[22]
port 131 nsew signal tristate
flabel metal3 s 59200 31968 60000 32088 0 FreeSans 480 0 0 0 io_out[23]
port 132 nsew signal tristate
flabel metal3 s 59200 33328 60000 33448 0 FreeSans 480 0 0 0 io_out[24]
port 133 nsew signal tristate
flabel metal3 s 59200 34688 60000 34808 0 FreeSans 480 0 0 0 io_out[25]
port 134 nsew signal tristate
flabel metal3 s 59200 36048 60000 36168 0 FreeSans 480 0 0 0 io_out[26]
port 135 nsew signal tristate
flabel metal3 s 59200 37408 60000 37528 0 FreeSans 480 0 0 0 io_out[27]
port 136 nsew signal tristate
flabel metal3 s 59200 38768 60000 38888 0 FreeSans 480 0 0 0 io_out[28]
port 137 nsew signal tristate
flabel metal3 s 59200 40128 60000 40248 0 FreeSans 480 0 0 0 io_out[29]
port 138 nsew signal tristate
flabel metal3 s 59200 3408 60000 3528 0 FreeSans 480 0 0 0 io_out[2]
port 139 nsew signal tristate
flabel metal3 s 59200 41488 60000 41608 0 FreeSans 480 0 0 0 io_out[30]
port 140 nsew signal tristate
flabel metal3 s 59200 42848 60000 42968 0 FreeSans 480 0 0 0 io_out[31]
port 141 nsew signal tristate
flabel metal3 s 59200 44208 60000 44328 0 FreeSans 480 0 0 0 io_out[32]
port 142 nsew signal tristate
flabel metal3 s 59200 45568 60000 45688 0 FreeSans 480 0 0 0 io_out[33]
port 143 nsew signal tristate
flabel metal3 s 59200 46928 60000 47048 0 FreeSans 480 0 0 0 io_out[34]
port 144 nsew signal tristate
flabel metal3 s 59200 48288 60000 48408 0 FreeSans 480 0 0 0 io_out[35]
port 145 nsew signal tristate
flabel metal3 s 59200 49648 60000 49768 0 FreeSans 480 0 0 0 io_out[36]
port 146 nsew signal tristate
flabel metal3 s 59200 51008 60000 51128 0 FreeSans 480 0 0 0 io_out[37]
port 147 nsew signal tristate
flabel metal3 s 59200 4768 60000 4888 0 FreeSans 480 0 0 0 io_out[3]
port 148 nsew signal tristate
flabel metal3 s 59200 6128 60000 6248 0 FreeSans 480 0 0 0 io_out[4]
port 149 nsew signal tristate
flabel metal3 s 59200 7488 60000 7608 0 FreeSans 480 0 0 0 io_out[5]
port 150 nsew signal tristate
flabel metal3 s 59200 8848 60000 8968 0 FreeSans 480 0 0 0 io_out[6]
port 151 nsew signal tristate
flabel metal3 s 59200 10208 60000 10328 0 FreeSans 480 0 0 0 io_out[7]
port 152 nsew signal tristate
flabel metal3 s 59200 11568 60000 11688 0 FreeSans 480 0 0 0 io_out[8]
port 153 nsew signal tristate
flabel metal3 s 59200 12928 60000 13048 0 FreeSans 480 0 0 0 io_out[9]
port 154 nsew signal tristate
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 irq[0]
port 155 nsew signal tristate
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 irq[1]
port 156 nsew signal tristate
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 irq[2]
port 157 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 158 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 159 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 160 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 161 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 162 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 163 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 164 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 165 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 166 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 167 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 168 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 169 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 170 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 171 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 172 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 173 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 174 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 175 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 176 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 177 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 178 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 179 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 180 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 181 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 182 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 183 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 184 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 185 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 186 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 187 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 188 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 189 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 190 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 191 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 192 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 193 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 194 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 195 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 196 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 197 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 198 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 199 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 200 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 201 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 202 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 203 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 204 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 205 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 206 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 207 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 208 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 209 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 210 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 211 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 212 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 213 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 214 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 215 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 216 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 217 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 218 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 219 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 220 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 221 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 222 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 223 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 224 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 225 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 226 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 227 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 228 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 229 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 230 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 231 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 232 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 233 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 234 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 235 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 236 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 237 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 238 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 239 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 240 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 241 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 242 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 243 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 244 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 245 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 246 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 247 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 248 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 249 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 250 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 251 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 252 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 253 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 254 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 255 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 256 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 257 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 258 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 259 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 260 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 261 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 262 nsew signal input
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 263 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 264 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 265 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 266 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 267 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 268 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 269 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 270 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 271 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 272 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 273 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 274 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 275 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 276 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 277 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 278 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 279 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 280 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 281 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 282 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 283 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 284 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 285 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 286 nsew signal tristate
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 287 nsew signal tristate
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 288 nsew signal tristate
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 289 nsew signal tristate
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 290 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 291 nsew signal tristate
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 292 nsew signal tristate
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 293 nsew signal tristate
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 294 nsew signal tristate
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 295 nsew signal tristate
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 296 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 297 nsew signal tristate
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 298 nsew signal tristate
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 299 nsew signal tristate
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 300 nsew signal tristate
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 301 nsew signal tristate
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 302 nsew signal tristate
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 303 nsew signal tristate
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 304 nsew signal tristate
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 305 nsew signal tristate
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 306 nsew signal tristate
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 307 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 308 nsew signal tristate
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 309 nsew signal tristate
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 310 nsew signal tristate
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 311 nsew signal tristate
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 312 nsew signal tristate
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 313 nsew signal tristate
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 314 nsew signal tristate
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 315 nsew signal tristate
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 316 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 317 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 318 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 319 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 320 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 321 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 322 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 323 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 324 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 325 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 326 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 327 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 328 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 329 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 330 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 331 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 332 nsew signal tristate
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 333 nsew signal tristate
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 334 nsew signal tristate
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 335 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 336 nsew signal tristate
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 337 nsew signal tristate
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 338 nsew signal tristate
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 339 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 340 nsew signal tristate
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 341 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 342 nsew signal tristate
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 343 nsew signal tristate
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 344 nsew signal tristate
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 345 nsew signal tristate
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 346 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 347 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 348 nsew signal tristate
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 349 nsew signal tristate
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 350 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 351 nsew signal tristate
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 352 nsew signal tristate
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 353 nsew signal tristate
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 354 nsew signal tristate
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 355 nsew signal tristate
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 356 nsew signal tristate
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 357 nsew signal tristate
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 358 nsew signal tristate
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 359 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 360 nsew signal tristate
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 361 nsew signal tristate
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 362 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 363 nsew signal tristate
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 364 nsew signal tristate
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 365 nsew signal tristate
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 366 nsew signal tristate
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 367 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 368 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 369 nsew signal tristate
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 370 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 371 nsew signal tristate
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 372 nsew signal tristate
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 373 nsew signal tristate
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 374 nsew signal tristate
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 375 nsew signal tristate
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 376 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 377 nsew signal tristate
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 378 nsew signal tristate
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 379 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 380 nsew signal tristate
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 381 nsew signal tristate
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 382 nsew signal tristate
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 383 nsew signal tristate
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 384 nsew signal tristate
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 385 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 386 nsew signal tristate
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 387 nsew signal tristate
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 388 nsew signal tristate
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 389 nsew signal tristate
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 390 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 391 nsew signal tristate
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 392 nsew signal tristate
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 393 nsew signal tristate
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 394 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 395 nsew signal tristate
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 396 nsew signal tristate
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 397 nsew signal tristate
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 398 nsew signal tristate
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 399 nsew signal tristate
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 400 nsew signal tristate
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 401 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 402 nsew signal tristate
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 403 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 404 nsew signal tristate
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 405 nsew signal tristate
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 406 nsew signal tristate
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 407 nsew signal tristate
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 408 nsew signal tristate
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 409 nsew signal tristate
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 410 nsew signal tristate
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 411 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 412 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 413 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 414 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 415 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 416 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 417 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 418 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 419 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 420 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 421 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 422 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 423 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 424 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 425 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 426 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 427 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 428 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 429 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 430 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 431 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 432 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 433 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 434 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 435 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 436 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 437 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 438 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 439 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 440 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 441 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 442 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 443 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 444 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 445 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 446 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 447 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 448 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 449 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 450 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 451 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 452 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 453 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 454 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 455 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 456 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 457 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 458 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 459 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 460 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 461 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 462 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 463 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 464 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 465 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 466 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 467 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 468 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 469 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 470 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 471 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 472 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 473 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 474 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 475 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 476 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 477 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 478 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 479 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 480 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 481 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 482 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 483 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 484 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 485 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 486 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 487 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 488 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 489 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 490 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 491 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 492 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 493 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 494 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 495 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 496 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 497 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 498 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 499 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 500 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 501 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 502 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 503 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 504 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 505 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 506 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 507 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 508 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 509 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 510 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 511 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 512 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 513 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 514 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 515 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 516 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 517 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 518 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 519 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 520 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 521 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 522 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 523 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 524 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 525 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 526 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 527 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 528 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 529 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 530 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 531 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 532 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 533 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 534 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 535 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 536 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 537 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 538 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 539 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 540 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 541 nsew signal input
flabel metal3 s 59200 53728 60000 53848 0 FreeSans 480 0 0 0 rst_o
port 542 nsew signal tristate
flabel metal3 s 59200 56448 60000 56568 0 FreeSans 480 0 0 0 start_o
port 543 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 544 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 544 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 545 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 545 nsew ground bidirectional
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 wb_clk_i
port 546 nsew signal input
flabel metal2 s 5630 0 5686 800 0 FreeSans 224 90 0 0 wb_rst_i
port 547 nsew signal input
flabel metal2 s 5722 0 5778 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 548 nsew signal tristate
flabel metal2 s 6090 0 6146 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 549 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 550 nsew signal input
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 551 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 552 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 553 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 554 nsew signal input
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 555 nsew signal input
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 556 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 557 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 558 nsew signal input
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 559 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 560 nsew signal input
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 561 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 562 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 563 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 564 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 565 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 566 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 567 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 568 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 569 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 570 nsew signal input
flabel metal2 s 6826 0 6882 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 571 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 572 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 573 nsew signal input
flabel metal2 s 7194 0 7250 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 574 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 575 nsew signal input
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 576 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 577 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 578 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 579 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 580 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 581 nsew signal input
flabel metal2 s 6182 0 6238 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 582 nsew signal input
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 583 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 584 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 585 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 586 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 587 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 588 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 589 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 590 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 591 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 592 nsew signal input
flabel metal2 s 6550 0 6606 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 593 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 594 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 595 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 596 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 597 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 598 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 599 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 600 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 601 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 602 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 603 nsew signal input
flabel metal2 s 6918 0 6974 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 604 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 605 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 606 nsew signal input
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 607 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 608 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 609 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 610 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 611 nsew signal input
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 612 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 613 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 614 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 615 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 616 nsew signal tristate
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 617 nsew signal tristate
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 618 nsew signal tristate
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 619 nsew signal tristate
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 620 nsew signal tristate
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 621 nsew signal tristate
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 622 nsew signal tristate
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 623 nsew signal tristate
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 624 nsew signal tristate
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 625 nsew signal tristate
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 626 nsew signal tristate
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 627 nsew signal tristate
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 628 nsew signal tristate
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 629 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 630 nsew signal tristate
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 631 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 632 nsew signal tristate
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 633 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 634 nsew signal tristate
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 635 nsew signal tristate
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 636 nsew signal tristate
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 637 nsew signal tristate
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 638 nsew signal tristate
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 639 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 640 nsew signal tristate
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 641 nsew signal tristate
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 642 nsew signal tristate
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 643 nsew signal tristate
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 644 nsew signal tristate
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 645 nsew signal tristate
flabel metal2 s 6366 0 6422 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 646 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 647 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 648 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 649 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 650 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 wbs_we_i
port 651 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
