VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO muler
  CLASS BLOCK ;
  FOREIGN muler ;
  ORIGIN 2.700 14.500 ;
  SIZE 13.700 BY 22.500 ;
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 1.875 -4.700 2.100 -4.100 ;
        RECT 3.550 -4.700 3.775 -4.100 ;
        RECT 4.700 -4.700 4.925 -4.100 ;
        RECT 1.425 -4.875 5.625 -4.700 ;
      LAYER mcon ;
        RECT 1.650 -4.875 1.825 -4.700 ;
        RECT 2.125 -4.875 2.300 -4.700 ;
        RECT 2.600 -4.875 2.775 -4.700 ;
        RECT 3.075 -4.875 3.250 -4.700 ;
        RECT 3.550 -4.875 3.725 -4.700 ;
        RECT 4.025 -4.875 4.200 -4.700 ;
        RECT 4.500 -4.875 4.675 -4.700 ;
        RECT 4.975 -4.875 5.150 -4.700 ;
      LAYER met1 ;
        RECT 1.425 -5.025 5.625 -4.550 ;
        RECT 1.500 -8.530 2.500 -5.025 ;
      LAYER via ;
        RECT 1.500 -8.500 2.500 -7.500 ;
      LAYER met2 ;
        RECT 1.000 -9.000 3.000 -7.000 ;
      LAYER via2 ;
        RECT 1.500 -8.500 2.500 -7.500 ;
      LAYER met3 ;
        RECT 1.000 -9.000 3.000 -7.000 ;
      LAYER via3 ;
        RECT 1.475 -8.525 2.525 -7.475 ;
      LAYER met4 ;
        RECT 1.470 -8.530 2.530 -7.470 ;
        RECT 1.500 -11.000 2.500 -8.530 ;
        RECT -0.500 -14.500 11.000 -11.000 ;
    END
  END VSS
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.425 -2.150 5.625 -1.975 ;
        RECT 1.850 -3.050 2.125 -2.150 ;
        RECT 3.500 -3.075 3.775 -2.150 ;
        RECT 4.650 -3.075 4.925 -2.150 ;
      LAYER mcon ;
        RECT 1.650 -2.150 1.825 -1.975 ;
        RECT 2.125 -2.150 2.300 -1.975 ;
        RECT 2.600 -2.150 2.775 -1.975 ;
        RECT 3.075 -2.150 3.250 -1.975 ;
        RECT 3.550 -2.150 3.725 -1.975 ;
        RECT 4.025 -2.150 4.200 -1.975 ;
        RECT 4.500 -2.150 4.675 -1.975 ;
        RECT 4.975 -2.150 5.150 -1.975 ;
      LAYER met1 ;
        RECT 1.520 -1.000 2.495 2.015 ;
        RECT 1.500 -1.825 2.500 -1.000 ;
        RECT 1.375 -2.300 5.625 -1.825 ;
      LAYER via ;
        RECT 1.520 1.010 2.495 1.985 ;
      LAYER met2 ;
        RECT 1.000 0.500 3.000 2.500 ;
      LAYER via2 ;
        RECT 1.520 1.010 2.495 1.985 ;
      LAYER met3 ;
        RECT 1.000 0.500 3.000 2.500 ;
      LAYER via3 ;
        RECT 1.495 0.985 2.520 2.010 ;
      LAYER met4 ;
        RECT -0.500 4.500 11.000 8.000 ;
        RECT 1.520 2.015 2.495 4.500 ;
        RECT 1.490 0.980 2.525 2.015 ;
    END
  END VDD
  PIN M
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.116250 ;
    PORT
      LAYER li1 ;
        RECT 2.000 -3.550 2.375 -3.250 ;
      LAYER mcon ;
        RECT 2.075 -3.500 2.275 -3.325 ;
      LAYER met1 ;
        RECT -2.700 -2.725 -0.600 -2.450 ;
        RECT -2.700 -2.975 1.725 -2.725 ;
        RECT -2.700 -3.250 -0.600 -2.975 ;
        RECT 1.475 -3.050 1.725 -2.975 ;
        RECT 1.475 -3.250 2.250 -3.050 ;
        RECT 1.475 -3.300 2.375 -3.250 ;
        RECT 2.000 -3.550 2.375 -3.300 ;
    END
  END M
  PIN P
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT -2.700 -3.650 -0.600 -3.450 ;
        RECT 1.425 -3.650 1.800 -3.625 ;
        RECT -2.700 -3.900 1.800 -3.650 ;
        RECT -2.700 -4.250 -0.600 -3.900 ;
        RECT 1.425 -3.925 1.800 -3.900 ;
    END
  END P
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.195000 ;
    PORT
      LAYER li1 ;
        RECT 2.600 -3.875 2.875 -3.500 ;
      LAYER mcon ;
        RECT 2.650 -3.775 2.825 -3.600 ;
      LAYER met1 ;
        RECT 2.600 -3.700 2.875 -3.500 ;
        RECT 2.600 -4.000 2.900 -3.700 ;
        RECT 2.600 -4.135 2.825 -4.000 ;
        RECT 0.040 -4.360 2.825 -4.135 ;
        RECT -2.700 -5.335 -0.600 -5.050 ;
        RECT 0.040 -5.335 0.265 -4.360 ;
        RECT -2.700 -5.560 0.265 -5.335 ;
        RECT -2.700 -5.850 -0.600 -5.560 ;
    END
  END C
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.195000 ;
    ANTENNADIFFAREA 0.780000 ;
    PORT
      LAYER li1 ;
        RECT 2.850 -3.075 3.125 -2.325 ;
        RECT 5.125 -2.350 5.400 -2.325 ;
        RECT 5.125 -3.075 5.500 -2.350 ;
        RECT 2.850 -3.275 3.275 -3.075 ;
        RECT 3.100 -3.450 3.275 -3.275 ;
        RECT 3.700 -3.450 3.975 -3.325 ;
        RECT 3.100 -3.675 3.975 -3.450 ;
        RECT 3.100 -4.050 3.275 -3.675 ;
        RECT 3.700 -3.700 3.975 -3.675 ;
        RECT 5.325 -3.875 5.500 -3.075 ;
        RECT 2.850 -4.275 3.275 -4.050 ;
        RECT 5.175 -4.150 5.550 -3.875 ;
        RECT 2.850 -4.500 3.150 -4.275 ;
        RECT 5.175 -4.500 5.400 -4.150 ;
      LAYER mcon ;
        RECT 3.750 -3.600 3.925 -3.425 ;
        RECT 5.275 -4.100 5.450 -3.925 ;
      LAYER met1 ;
        RECT 3.700 -3.525 3.975 -3.325 ;
        RECT 3.700 -3.700 4.250 -3.525 ;
        RECT 4.100 -3.950 4.250 -3.700 ;
        RECT 5.175 -3.950 5.550 -3.875 ;
        RECT 6.100 -3.950 8.200 -3.600 ;
        RECT 4.100 -4.100 8.200 -3.950 ;
        RECT 5.175 -4.150 5.550 -4.100 ;
        RECT 6.100 -4.400 8.200 -4.100 ;
    END
  END OUT
  OBS
      LAYER nwell ;
        RECT 1.425 -3.500 5.625 -1.875 ;
      LAYER pwell ;
        RECT 1.600 -3.925 5.625 -3.900 ;
        RECT 1.425 -4.875 5.625 -3.925 ;
      LAYER li1 ;
        RECT 3.975 -2.350 4.250 -2.325 ;
        RECT 3.975 -3.075 4.350 -2.350 ;
        RECT 4.175 -3.500 4.350 -3.075 ;
        RECT 4.850 -3.500 5.125 -3.325 ;
        RECT 1.425 -3.925 1.800 -3.625 ;
        RECT 4.175 -3.700 5.125 -3.500 ;
        RECT 4.175 -3.900 4.350 -3.700 ;
        RECT 4.025 -4.100 4.350 -3.900 ;
        RECT 4.025 -4.500 4.250 -4.100 ;
  END
END muler
END LIBRARY

