magic
tech sky130B
magscale 1 2
timestamp 1667927669
<< viali >>
rect 4353 57409 4387 57443
rect 4997 57409 5031 57443
rect 5825 57409 5859 57443
rect 6653 57409 6687 57443
rect 7573 57409 7607 57443
rect 8217 57409 8251 57443
rect 9321 57409 9355 57443
rect 9965 57409 9999 57443
rect 10977 57409 11011 57443
rect 11621 57409 11655 57443
rect 12633 57409 12667 57443
rect 13277 57409 13311 57443
rect 14289 57409 14323 57443
rect 14933 57409 14967 57443
rect 15945 57409 15979 57443
rect 17601 57409 17635 57443
rect 18245 57409 18279 57443
rect 19257 57409 19291 57443
rect 19901 57409 19935 57443
rect 21005 57409 21039 57443
rect 21833 57409 21867 57443
rect 22569 57409 22603 57443
rect 23213 57409 23247 57443
rect 24869 57409 24903 57443
rect 25789 57409 25823 57443
rect 26433 57409 26467 57443
rect 27537 57409 27571 57443
rect 28181 57409 28215 57443
rect 29009 57409 29043 57443
rect 29837 57409 29871 57443
rect 30757 57409 30791 57443
rect 31401 57409 31435 57443
rect 32505 57409 32539 57443
rect 33149 57409 33183 57443
rect 34161 57409 34195 57443
rect 34805 57409 34839 57443
rect 36553 57409 36587 57443
rect 37565 57409 37599 57443
rect 38209 57409 38243 57443
rect 39865 57409 39899 57443
rect 40509 57409 40543 57443
rect 41153 57409 41187 57443
rect 42533 57409 42567 57443
rect 43177 57409 43211 57443
rect 44189 57409 44223 57443
rect 45017 57409 45051 57443
rect 45845 57409 45879 57443
rect 46489 57409 46523 57443
rect 47593 57409 47627 57443
rect 48237 57409 48271 57443
rect 49157 57409 49191 57443
rect 50169 57409 50203 57443
rect 50813 57409 50847 57443
rect 51457 57409 51491 57443
rect 52745 57409 52779 57443
rect 53389 57409 53423 57443
rect 54125 57409 54159 57443
rect 55965 57409 55999 57443
rect 56609 57409 56643 57443
rect 57897 57409 57931 57443
rect 58541 57409 58575 57443
rect 59185 57409 59219 57443
rect 60473 57409 60507 57443
rect 61117 57409 61151 57443
rect 61761 57409 61795 57443
rect 63049 57409 63083 57443
rect 64337 57409 64371 57443
rect 65717 57409 65751 57443
rect 66361 57409 66395 57443
rect 16681 57341 16715 57375
rect 35909 57341 35943 57375
rect 63693 57341 63727 57375
rect 55321 57273 55355 57307
rect 24409 57001 24443 57035
rect 41429 57001 41463 57035
rect 64613 57001 64647 57035
rect 67373 56321 67407 56355
rect 67557 56117 67591 56151
rect 67373 48705 67407 48739
rect 67557 48569 67591 48603
rect 66637 45441 66671 45475
rect 67189 45441 67223 45475
rect 67373 45305 67407 45339
rect 67833 41565 67867 41599
rect 67281 41429 67315 41463
rect 68017 41429 68051 41463
rect 67373 39593 67407 39627
rect 67189 39389 67223 39423
rect 67833 39389 67867 39423
rect 27629 34357 27663 34391
rect 27721 34017 27755 34051
rect 28181 34017 28215 34051
rect 26709 33949 26743 33983
rect 26985 33949 27019 33983
rect 27813 33949 27847 33983
rect 67833 33949 67867 33983
rect 26801 33881 26835 33915
rect 13185 33813 13219 33847
rect 27169 33813 27203 33847
rect 28825 33813 28859 33847
rect 68017 33813 68051 33847
rect 13185 33609 13219 33643
rect 28181 33541 28215 33575
rect 28917 33541 28951 33575
rect 8769 33473 8803 33507
rect 13001 33473 13035 33507
rect 13277 33473 13311 33507
rect 13921 33473 13955 33507
rect 14565 33473 14599 33507
rect 14749 33473 14783 33507
rect 24041 33473 24075 33507
rect 24685 33473 24719 33507
rect 25973 33473 26007 33507
rect 27169 33473 27203 33507
rect 27813 33473 27847 33507
rect 27951 33473 27985 33507
rect 28089 33473 28123 33507
rect 28297 33473 28331 33507
rect 29101 33473 29135 33507
rect 35173 33473 35207 33507
rect 35357 33473 35391 33507
rect 8861 33405 8895 33439
rect 13737 33405 13771 33439
rect 24593 33405 24627 33439
rect 26065 33405 26099 33439
rect 26985 33405 27019 33439
rect 29377 33405 29411 33439
rect 37289 33405 37323 33439
rect 9137 33337 9171 33371
rect 14565 33337 14599 33371
rect 25053 33337 25087 33371
rect 26341 33337 26375 33371
rect 27353 33337 27387 33371
rect 28457 33337 28491 33371
rect 35909 33337 35943 33371
rect 12817 33269 12851 33303
rect 14105 33269 14139 33303
rect 15301 33269 15335 33303
rect 29285 33269 29319 33303
rect 34621 33269 34655 33303
rect 35357 33269 35391 33303
rect 16221 33065 16255 33099
rect 26065 33065 26099 33099
rect 26801 33065 26835 33099
rect 34069 33065 34103 33099
rect 12541 32997 12575 33031
rect 19349 32997 19383 33031
rect 27813 32997 27847 33031
rect 9781 32929 9815 32963
rect 13001 32929 13035 32963
rect 15117 32929 15151 32963
rect 16589 32929 16623 32963
rect 27353 32929 27387 32963
rect 28825 32929 28859 32963
rect 35081 32929 35115 32963
rect 36277 32929 36311 32963
rect 37105 32929 37139 32963
rect 38485 32929 38519 32963
rect 9689 32861 9723 32895
rect 12909 32861 12943 32895
rect 14289 32861 14323 32895
rect 14473 32861 14507 32895
rect 14565 32861 14599 32895
rect 15025 32861 15059 32895
rect 15209 32861 15243 32895
rect 16405 32861 16439 32895
rect 17141 32861 17175 32895
rect 18061 32861 18095 32895
rect 22201 32861 22235 32895
rect 24685 32861 24719 32895
rect 25145 32861 25179 32895
rect 25329 32861 25363 32895
rect 25973 32861 26007 32895
rect 26617 32861 26651 32895
rect 26801 32861 26835 32895
rect 27445 32861 27479 32895
rect 28273 32861 28307 32895
rect 28365 32861 28399 32895
rect 28549 32861 28583 32895
rect 28641 32861 28675 32895
rect 29561 32861 29595 32895
rect 29745 32861 29779 32895
rect 32413 32861 32447 32895
rect 35265 32861 35299 32895
rect 36185 32861 36219 32895
rect 37013 32861 37047 32895
rect 37197 32861 37231 32895
rect 38301 32861 38335 32895
rect 25513 32793 25547 32827
rect 29653 32793 29687 32827
rect 35449 32793 35483 32827
rect 10057 32725 10091 32759
rect 14105 32725 14139 32759
rect 15669 32725 15703 32759
rect 18245 32725 18279 32759
rect 21557 32725 21591 32759
rect 22477 32725 22511 32759
rect 32505 32725 32539 32759
rect 36553 32725 36587 32759
rect 38117 32725 38151 32759
rect 25421 32521 25455 32555
rect 28641 32521 28675 32555
rect 38669 32521 38703 32555
rect 14197 32453 14231 32487
rect 24869 32453 24903 32487
rect 34621 32453 34655 32487
rect 6561 32385 6595 32419
rect 9045 32385 9079 32419
rect 12725 32385 12759 32419
rect 13829 32385 13863 32419
rect 13922 32385 13956 32419
rect 14105 32385 14139 32419
rect 14335 32385 14369 32419
rect 15485 32385 15519 32419
rect 16037 32385 16071 32419
rect 18613 32385 18647 32419
rect 23213 32385 23247 32419
rect 25329 32385 25363 32419
rect 25513 32385 25547 32419
rect 26433 32385 26467 32419
rect 27445 32385 27479 32419
rect 28825 32385 28859 32419
rect 29009 32385 29043 32419
rect 33517 32385 33551 32419
rect 34529 32385 34563 32419
rect 35725 32385 35759 32419
rect 36553 32385 36587 32419
rect 37473 32385 37507 32419
rect 37749 32385 37783 32419
rect 38577 32385 38611 32419
rect 38853 32385 38887 32419
rect 39865 32385 39899 32419
rect 9137 32317 9171 32351
rect 12817 32317 12851 32351
rect 17693 32317 17727 32351
rect 17969 32317 18003 32351
rect 34805 32317 34839 32351
rect 35541 32317 35575 32351
rect 35633 32317 35667 32351
rect 39957 32317 39991 32351
rect 12357 32249 12391 32283
rect 19165 32249 19199 32283
rect 27629 32249 27663 32283
rect 34161 32249 34195 32283
rect 36645 32249 36679 32283
rect 37657 32249 37691 32283
rect 6377 32181 6411 32215
rect 9321 32181 9355 32215
rect 14473 32181 14507 32215
rect 15301 32181 15335 32215
rect 18429 32181 18463 32215
rect 23029 32181 23063 32215
rect 33701 32181 33735 32215
rect 36093 32181 36127 32215
rect 37289 32181 37323 32215
rect 39037 32181 39071 32215
rect 40141 32181 40175 32215
rect 7113 31977 7147 32011
rect 8401 31977 8435 32011
rect 13369 31977 13403 32011
rect 14197 31977 14231 32011
rect 16405 31977 16439 32011
rect 19349 31977 19383 32011
rect 22017 31977 22051 32011
rect 25789 31977 25823 32011
rect 36093 31977 36127 32011
rect 18705 31909 18739 31943
rect 23857 31909 23891 31943
rect 28365 31909 28399 31943
rect 37933 31909 37967 31943
rect 38945 31909 38979 31943
rect 57897 31909 57931 31943
rect 7665 31841 7699 31875
rect 27721 31841 27755 31875
rect 27905 31841 27939 31875
rect 38485 31841 38519 31875
rect 39957 31841 39991 31875
rect 41153 31841 41187 31875
rect 5273 31773 5307 31807
rect 7573 31773 7607 31807
rect 11989 31773 12023 31807
rect 14105 31773 14139 31807
rect 15025 31773 15059 31807
rect 17325 31773 17359 31807
rect 19441 31773 19475 31807
rect 20637 31773 20671 31807
rect 22477 31773 22511 31807
rect 24409 31773 24443 31807
rect 29009 31773 29043 31807
rect 31217 31773 31251 31807
rect 34713 31773 34747 31807
rect 37289 31773 37323 31807
rect 37437 31773 37471 31807
rect 37565 31773 37599 31807
rect 37754 31773 37788 31807
rect 38577 31773 38611 31807
rect 40049 31773 40083 31807
rect 41245 31773 41279 31807
rect 41889 31773 41923 31807
rect 57713 31773 57747 31807
rect 58357 31773 58391 31807
rect 5540 31705 5574 31739
rect 12256 31705 12290 31739
rect 15292 31705 15326 31739
rect 17592 31705 17626 31739
rect 20904 31705 20938 31739
rect 22744 31705 22778 31739
rect 24654 31705 24688 31739
rect 31484 31705 31518 31739
rect 34980 31705 35014 31739
rect 37657 31705 37691 31739
rect 6653 31637 6687 31671
rect 7481 31637 7515 31671
rect 19993 31637 20027 31671
rect 27169 31637 27203 31671
rect 27997 31637 28031 31671
rect 28825 31637 28859 31671
rect 32597 31637 32631 31671
rect 34069 31637 34103 31671
rect 36553 31637 36587 31671
rect 40417 31637 40451 31671
rect 40877 31637 40911 31671
rect 42073 31637 42107 31671
rect 5457 31433 5491 31467
rect 8217 31433 8251 31467
rect 12633 31433 12667 31467
rect 13277 31433 13311 31467
rect 13645 31433 13679 31467
rect 15393 31433 15427 31467
rect 15761 31433 15795 31467
rect 17325 31433 17359 31467
rect 19533 31433 19567 31467
rect 21005 31433 21039 31467
rect 21833 31433 21867 31467
rect 22293 31433 22327 31467
rect 23213 31433 23247 31467
rect 23673 31433 23707 31467
rect 24501 31433 24535 31467
rect 25145 31433 25179 31467
rect 25605 31433 25639 31467
rect 27537 31433 27571 31467
rect 29745 31433 29779 31467
rect 31401 31433 31435 31467
rect 32505 31433 32539 31467
rect 33425 31433 33459 31467
rect 35265 31433 35299 31467
rect 35725 31433 35759 31467
rect 41061 31433 41095 31467
rect 41521 31433 41555 31467
rect 6644 31365 6678 31399
rect 22201 31365 22235 31399
rect 28632 31365 28666 31399
rect 37534 31365 37568 31399
rect 40325 31365 40359 31399
rect 41153 31365 41187 31399
rect 8401 31297 8435 31331
rect 9137 31297 9171 31331
rect 9965 31297 9999 31331
rect 10241 31297 10275 31331
rect 12817 31297 12851 31331
rect 18153 31297 18187 31331
rect 18420 31297 18454 31331
rect 20177 31297 20211 31331
rect 21189 31297 21223 31331
rect 23581 31297 23615 31331
rect 24685 31297 24719 31331
rect 25513 31297 25547 31331
rect 27169 31297 27203 31331
rect 31585 31297 31619 31331
rect 34141 31297 34175 31331
rect 35909 31297 35943 31331
rect 36553 31297 36587 31331
rect 37289 31297 37323 31331
rect 42441 31297 42475 31331
rect 5549 31229 5583 31263
rect 5733 31229 5767 31263
rect 6377 31229 6411 31263
rect 9229 31229 9263 31263
rect 10057 31229 10091 31263
rect 13737 31229 13771 31263
rect 13829 31229 13863 31263
rect 15853 31229 15887 31263
rect 15945 31229 15979 31263
rect 17141 31229 17175 31263
rect 17233 31229 17267 31263
rect 22477 31229 22511 31263
rect 23765 31229 23799 31263
rect 25697 31229 25731 31263
rect 27077 31229 27111 31263
rect 28365 31229 28399 31263
rect 32597 31229 32631 31263
rect 32689 31229 32723 31263
rect 33885 31229 33919 31263
rect 40969 31229 41003 31263
rect 4629 31161 4663 31195
rect 7757 31161 7791 31195
rect 9505 31161 9539 31195
rect 20361 31161 20395 31195
rect 36737 31161 36771 31195
rect 5089 31093 5123 31127
rect 9965 31093 9999 31127
rect 10425 31093 10459 31127
rect 14933 31093 14967 31127
rect 17693 31093 17727 31127
rect 32137 31093 32171 31127
rect 38669 31093 38703 31127
rect 42625 31093 42659 31127
rect 5365 30889 5399 30923
rect 7205 30889 7239 30923
rect 8401 30889 8435 30923
rect 16589 30889 16623 30923
rect 17509 30889 17543 30923
rect 18705 30889 18739 30923
rect 19809 30889 19843 30923
rect 22477 30889 22511 30923
rect 36461 30889 36495 30923
rect 37013 30889 37047 30923
rect 41245 30889 41279 30923
rect 27077 30821 27111 30855
rect 31493 30821 31527 30855
rect 5825 30753 5859 30787
rect 7757 30753 7791 30787
rect 18153 30753 18187 30787
rect 25697 30753 25731 30787
rect 27997 30753 28031 30787
rect 28089 30753 28123 30787
rect 30205 30753 30239 30787
rect 37473 30753 37507 30787
rect 37565 30753 37599 30787
rect 5181 30685 5215 30719
rect 6092 30685 6126 30719
rect 8033 30685 8067 30719
rect 9045 30685 9079 30719
rect 12173 30685 12207 30719
rect 15485 30685 15519 30719
rect 17325 30685 17359 30719
rect 20637 30685 20671 30719
rect 24685 30685 24719 30719
rect 25237 30685 25271 30719
rect 29009 30685 29043 30719
rect 31309 30685 31343 30719
rect 31953 30685 31987 30719
rect 32209 30685 32243 30719
rect 42358 30685 42392 30719
rect 42625 30685 42659 30719
rect 7941 30617 7975 30651
rect 11906 30617 11940 30651
rect 14197 30617 14231 30651
rect 15025 30617 15059 30651
rect 16497 30617 16531 30651
rect 19717 30617 19751 30651
rect 20904 30617 20938 30651
rect 23121 30617 23155 30651
rect 25964 30617 25998 30651
rect 30021 30617 30055 30651
rect 35909 30617 35943 30651
rect 37381 30617 37415 30651
rect 10793 30549 10827 30583
rect 15669 30549 15703 30583
rect 18245 30549 18279 30583
rect 18337 30549 18371 30583
rect 22017 30549 22051 30583
rect 24501 30549 24535 30583
rect 27537 30549 27571 30583
rect 27905 30549 27939 30583
rect 29561 30549 29595 30583
rect 29929 30549 29963 30583
rect 33333 30549 33367 30583
rect 10333 30345 10367 30379
rect 11713 30345 11747 30379
rect 15393 30345 15427 30379
rect 18061 30345 18095 30379
rect 21097 30345 21131 30379
rect 25973 30345 26007 30379
rect 32137 30345 32171 30379
rect 41889 30345 41923 30379
rect 17325 30277 17359 30311
rect 17969 30277 18003 30311
rect 18613 30277 18647 30311
rect 24308 30277 24342 30311
rect 31493 30277 31527 30311
rect 32597 30277 32631 30311
rect 43554 30277 43588 30311
rect 10701 30209 10735 30243
rect 11529 30209 11563 30243
rect 15761 30209 15795 30243
rect 21281 30209 21315 30243
rect 22201 30209 22235 30243
rect 26157 30209 26191 30243
rect 28273 30209 28307 30243
rect 28540 30209 28574 30243
rect 30849 30209 30883 30243
rect 32505 30209 32539 30243
rect 36461 30209 36495 30243
rect 40417 30209 40451 30243
rect 40693 30209 40727 30243
rect 41521 30209 41555 30243
rect 43821 30209 43855 30243
rect 10793 30141 10827 30175
rect 14933 30141 14967 30175
rect 15853 30141 15887 30175
rect 15945 30141 15979 30175
rect 22293 30141 22327 30175
rect 22477 30141 22511 30175
rect 24041 30141 24075 30175
rect 27353 30141 27387 30175
rect 32689 30141 32723 30175
rect 40601 30141 40635 30175
rect 41337 30141 41371 30175
rect 41429 30141 41463 30175
rect 19441 30073 19475 30107
rect 21833 30073 21867 30107
rect 42441 30073 42475 30107
rect 16865 30005 16899 30039
rect 20085 30005 20119 30039
rect 25421 30005 25455 30039
rect 29653 30005 29687 30039
rect 30665 30005 30699 30039
rect 36277 30005 36311 30039
rect 40233 30005 40267 30039
rect 40693 30005 40727 30039
rect 11805 29801 11839 29835
rect 16681 29801 16715 29835
rect 24777 29801 24811 29835
rect 28825 29801 28859 29835
rect 37841 29801 37875 29835
rect 41337 29801 41371 29835
rect 67373 29801 67407 29835
rect 6285 29733 6319 29767
rect 7297 29733 7331 29767
rect 9505 29733 9539 29767
rect 40693 29733 40727 29767
rect 7021 29665 7055 29699
rect 9045 29665 9079 29699
rect 12357 29665 12391 29699
rect 25421 29665 25455 29699
rect 30481 29665 30515 29699
rect 36001 29665 36035 29699
rect 41521 29665 41555 29699
rect 4905 29597 4939 29631
rect 6929 29597 6963 29631
rect 9137 29597 9171 29631
rect 10977 29597 11011 29631
rect 11161 29597 11195 29631
rect 15301 29597 15335 29631
rect 15568 29597 15602 29631
rect 17509 29597 17543 29631
rect 17969 29597 18003 29631
rect 19441 29597 19475 29631
rect 20453 29597 20487 29631
rect 21649 29597 21683 29631
rect 29009 29597 29043 29631
rect 30748 29597 30782 29631
rect 35357 29597 35391 29631
rect 41613 29597 41647 29631
rect 67189 29597 67223 29631
rect 67833 29597 67867 29631
rect 5172 29529 5206 29563
rect 12173 29529 12207 29563
rect 17141 29529 17175 29563
rect 20269 29529 20303 29563
rect 25237 29529 25271 29563
rect 36246 29529 36280 29563
rect 11345 29461 11379 29495
rect 12265 29461 12299 29495
rect 13093 29461 13127 29495
rect 14749 29461 14783 29495
rect 19257 29461 19291 29495
rect 23857 29461 23891 29495
rect 25145 29461 25179 29495
rect 31861 29461 31895 29495
rect 35541 29461 35575 29495
rect 37381 29461 37415 29495
rect 43085 29461 43119 29495
rect 5273 29257 5307 29291
rect 6745 29257 6779 29291
rect 12909 29257 12943 29291
rect 37289 29257 37323 29291
rect 37657 29257 37691 29291
rect 40049 29257 40083 29291
rect 41061 29257 41095 29291
rect 45109 29257 45143 29291
rect 6837 29189 6871 29223
rect 7573 29189 7607 29223
rect 9321 29189 9355 29223
rect 10425 29189 10459 29223
rect 15945 29189 15979 29223
rect 35164 29189 35198 29223
rect 42809 29189 42843 29223
rect 5457 29121 5491 29155
rect 9137 29121 9171 29155
rect 10333 29121 10367 29155
rect 10609 29121 10643 29155
rect 11529 29121 11563 29155
rect 11713 29121 11747 29155
rect 12541 29121 12575 29155
rect 14381 29121 14415 29155
rect 15209 29121 15243 29155
rect 15761 29121 15795 29155
rect 16681 29121 16715 29155
rect 16865 29121 16899 29155
rect 19450 29121 19484 29155
rect 19717 29121 19751 29155
rect 22109 29121 22143 29155
rect 24593 29121 24627 29155
rect 31329 29121 31363 29155
rect 31585 29121 31619 29155
rect 32321 29121 32355 29155
rect 38669 29121 38703 29155
rect 39681 29121 39715 29155
rect 40693 29121 40727 29155
rect 43269 29121 43303 29155
rect 43361 29121 43395 29155
rect 43545 29121 43579 29155
rect 44465 29121 44499 29155
rect 44925 29121 44959 29155
rect 6929 29053 6963 29087
rect 8953 29053 8987 29087
rect 12633 29053 12667 29087
rect 14289 29053 14323 29087
rect 34897 29053 34931 29087
rect 37749 29053 37783 29087
rect 37841 29053 37875 29087
rect 38761 29053 38795 29087
rect 39589 29053 39623 29087
rect 40601 29053 40635 29087
rect 6377 28985 6411 29019
rect 10793 28985 10827 29019
rect 11897 28985 11931 29019
rect 14013 28985 14047 29019
rect 17417 28985 17451 29019
rect 32137 28985 32171 29019
rect 36277 28985 36311 29019
rect 39037 28985 39071 29019
rect 43729 28985 43763 29019
rect 16681 28917 16715 28951
rect 18337 28917 18371 28951
rect 21925 28917 21959 28951
rect 24777 28917 24811 28951
rect 30205 28917 30239 28951
rect 44281 28917 44315 28951
rect 8953 28713 8987 28747
rect 10149 28713 10183 28747
rect 10977 28713 11011 28747
rect 12725 28713 12759 28747
rect 14105 28713 14139 28747
rect 14565 28713 14599 28747
rect 19257 28713 19291 28747
rect 30849 28713 30883 28747
rect 38485 28645 38519 28679
rect 9137 28577 9171 28611
rect 14197 28577 14231 28611
rect 16497 28577 16531 28611
rect 19901 28577 19935 28611
rect 21741 28577 21775 28611
rect 27813 28577 27847 28611
rect 31401 28577 31435 28611
rect 32229 28577 32263 28611
rect 35081 28577 35115 28611
rect 36093 28577 36127 28611
rect 38025 28577 38059 28611
rect 45017 28577 45051 28611
rect 9229 28509 9263 28543
rect 11621 28509 11655 28543
rect 11714 28509 11748 28543
rect 11897 28509 11931 28543
rect 12086 28509 12120 28543
rect 12909 28509 12943 28543
rect 13185 28509 13219 28543
rect 14105 28509 14139 28543
rect 14381 28509 14415 28543
rect 15209 28509 15243 28543
rect 16037 28509 16071 28543
rect 16773 28509 16807 28543
rect 17785 28509 17819 28543
rect 19717 28509 19751 28543
rect 22008 28509 22042 28543
rect 24409 28509 24443 28543
rect 24676 28509 24710 28543
rect 27905 28509 27939 28543
rect 32321 28509 32355 28543
rect 35173 28509 35207 28543
rect 36360 28509 36394 28543
rect 38117 28509 38151 28543
rect 38945 28509 38979 28543
rect 42257 28509 42291 28543
rect 42809 28509 42843 28543
rect 42993 28509 43027 28543
rect 43453 28509 43487 28543
rect 43729 28509 43763 28543
rect 45293 28509 45327 28543
rect 46121 28509 46155 28543
rect 11989 28441 12023 28475
rect 13093 28441 13127 28475
rect 17049 28441 17083 28475
rect 19625 28441 19659 28475
rect 20545 28441 20579 28475
rect 21097 28441 21131 28475
rect 30389 28441 30423 28475
rect 31217 28441 31251 28475
rect 42901 28441 42935 28475
rect 9597 28373 9631 28407
rect 12265 28373 12299 28407
rect 16681 28373 16715 28407
rect 16865 28373 16899 28407
rect 17601 28373 17635 28407
rect 18429 28373 18463 28407
rect 21189 28373 21223 28407
rect 23121 28373 23155 28407
rect 25789 28373 25823 28407
rect 28273 28373 28307 28407
rect 31309 28373 31343 28407
rect 32689 28373 32723 28407
rect 35265 28373 35299 28407
rect 35633 28373 35667 28407
rect 37473 28373 37507 28407
rect 44465 28373 44499 28407
rect 6929 28169 6963 28203
rect 10425 28169 10459 28203
rect 11713 28169 11747 28203
rect 12633 28169 12667 28203
rect 14197 28169 14231 28203
rect 15577 28169 15611 28203
rect 20177 28169 20211 28203
rect 21281 28169 21315 28203
rect 22109 28169 22143 28203
rect 22569 28169 22603 28203
rect 23397 28169 23431 28203
rect 24409 28169 24443 28203
rect 24777 28169 24811 28203
rect 27353 28169 27387 28203
rect 31217 28169 31251 28203
rect 31585 28169 31619 28203
rect 32689 28169 32723 28203
rect 35081 28169 35115 28203
rect 36001 28169 36035 28203
rect 36461 28169 36495 28203
rect 37841 28169 37875 28203
rect 38117 28169 38151 28203
rect 45477 28169 45511 28203
rect 45937 28169 45971 28203
rect 33149 28101 33183 28135
rect 37289 28101 37323 28135
rect 38025 28101 38059 28135
rect 38577 28101 38611 28135
rect 44005 28101 44039 28135
rect 6561 28033 6595 28067
rect 7389 28033 7423 28067
rect 10793 28033 10827 28067
rect 11621 28033 11655 28067
rect 11897 28033 11931 28067
rect 12541 28033 12575 28067
rect 12725 28033 12759 28067
rect 14565 28033 14599 28067
rect 15393 28033 15427 28067
rect 15669 28033 15703 28067
rect 17785 28033 17819 28067
rect 18889 28033 18923 28067
rect 19349 28033 19383 28067
rect 20913 28033 20947 28067
rect 22477 28033 22511 28067
rect 24869 28033 24903 28067
rect 26249 28033 26283 28067
rect 28365 28033 28399 28067
rect 30021 28033 30055 28067
rect 31125 28033 31159 28067
rect 32321 28033 32355 28067
rect 33425 28033 33459 28067
rect 35265 28033 35299 28067
rect 36369 28033 36403 28067
rect 40877 28033 40911 28067
rect 43729 28033 43763 28067
rect 46121 28033 46155 28067
rect 6469 27965 6503 27999
rect 10701 27965 10735 27999
rect 14657 27965 14691 27999
rect 15209 27965 15243 27999
rect 20821 27965 20855 27999
rect 22753 27965 22787 27999
rect 24961 27965 24995 27999
rect 27445 27965 27479 27999
rect 27537 27965 27571 27999
rect 28273 27965 28307 27999
rect 29929 27965 29963 27999
rect 30941 27965 30975 27999
rect 32229 27965 32263 27999
rect 33241 27965 33275 27999
rect 36553 27965 36587 27999
rect 46305 27965 46339 27999
rect 19533 27897 19567 27931
rect 26985 27897 27019 27931
rect 30389 27897 30423 27931
rect 38577 27897 38611 27931
rect 8861 27829 8895 27863
rect 12081 27829 12115 27863
rect 13369 27829 13403 27863
rect 17233 27829 17267 27863
rect 18337 27829 18371 27863
rect 26065 27829 26099 27863
rect 28641 27829 28675 27863
rect 33149 27829 33183 27863
rect 33609 27829 33643 27863
rect 6469 27625 6503 27659
rect 11713 27625 11747 27659
rect 27905 27625 27939 27659
rect 35909 27625 35943 27659
rect 37933 27625 37967 27659
rect 9229 27557 9263 27591
rect 18613 27557 18647 27591
rect 20729 27557 20763 27591
rect 20913 27557 20947 27591
rect 30113 27557 30147 27591
rect 31677 27557 31711 27591
rect 40325 27557 40359 27591
rect 45017 27557 45051 27591
rect 45201 27557 45235 27591
rect 9965 27489 9999 27523
rect 15025 27489 15059 27523
rect 19809 27489 19843 27523
rect 21741 27489 21775 27523
rect 24593 27489 24627 27523
rect 25973 27489 26007 27523
rect 29653 27489 29687 27523
rect 31217 27489 31251 27523
rect 41153 27489 41187 27523
rect 43453 27489 43487 27523
rect 45477 27489 45511 27523
rect 4445 27421 4479 27455
rect 5089 27421 5123 27455
rect 7113 27421 7147 27455
rect 8953 27421 8987 27455
rect 9873 27421 9907 27455
rect 11529 27421 11563 27455
rect 11713 27421 11747 27455
rect 14749 27421 14783 27455
rect 14933 27421 14967 27455
rect 17233 27421 17267 27455
rect 19717 27421 19751 27455
rect 21649 27421 21683 27455
rect 22477 27421 22511 27455
rect 22661 27421 22695 27455
rect 24763 27421 24797 27455
rect 28089 27421 28123 27455
rect 28365 27421 28399 27455
rect 28825 27421 28859 27455
rect 29009 27421 29043 27455
rect 29745 27421 29779 27455
rect 31309 27421 31343 27455
rect 36645 27421 36679 27455
rect 36829 27421 36863 27455
rect 39129 27421 39163 27455
rect 39313 27421 39347 27455
rect 39865 27421 39899 27455
rect 40141 27421 40175 27455
rect 41429 27421 41463 27455
rect 42257 27421 42291 27455
rect 43729 27421 43763 27455
rect 5356 27353 5390 27387
rect 9229 27353 9263 27387
rect 12265 27353 12299 27387
rect 17478 27353 17512 27387
rect 19349 27353 19383 27387
rect 19441 27353 19475 27387
rect 20453 27353 20487 27387
rect 22569 27353 22603 27387
rect 26240 27353 26274 27387
rect 28273 27353 28307 27387
rect 37289 27353 37323 27387
rect 4629 27285 4663 27319
rect 6929 27285 6963 27319
rect 9045 27285 9079 27319
rect 10241 27285 10275 27319
rect 11069 27285 11103 27319
rect 12909 27285 12943 27319
rect 15577 27285 15611 27319
rect 19993 27285 20027 27319
rect 22017 27285 22051 27319
rect 23397 27285 23431 27319
rect 25053 27285 25087 27319
rect 27353 27285 27387 27319
rect 29009 27285 29043 27319
rect 36737 27285 36771 27319
rect 38669 27285 38703 27319
rect 39221 27285 39255 27319
rect 39957 27285 39991 27319
rect 41337 27285 41371 27319
rect 41797 27285 41831 27319
rect 42441 27285 42475 27319
rect 44465 27285 44499 27319
rect 7757 27081 7791 27115
rect 8769 27081 8803 27115
rect 12633 27081 12667 27115
rect 13645 27081 13679 27115
rect 17325 27081 17359 27115
rect 19441 27081 19475 27115
rect 20361 27081 20395 27115
rect 23213 27081 23247 27115
rect 24225 27081 24259 27115
rect 25421 27081 25455 27115
rect 27445 27081 27479 27115
rect 36277 27081 36311 27115
rect 39129 27081 39163 27115
rect 40693 27081 40727 27115
rect 45385 27081 45419 27115
rect 45937 27081 45971 27115
rect 6644 27013 6678 27047
rect 31217 27013 31251 27047
rect 39865 27013 39899 27047
rect 43913 27013 43947 27047
rect 4445 26945 4479 26979
rect 4712 26945 4746 26979
rect 8309 26945 8343 26979
rect 9413 26945 9447 26979
rect 10609 26945 10643 26979
rect 12357 26945 12391 26979
rect 13093 26945 13127 26979
rect 13185 26945 13219 26979
rect 13369 26945 13403 26979
rect 13461 26945 13495 26979
rect 17141 26945 17175 26979
rect 18328 26945 18362 26979
rect 20269 26945 20303 26979
rect 21097 26945 21131 26979
rect 22845 26945 22879 26979
rect 24317 26945 24351 26979
rect 25053 26945 25087 26979
rect 27537 26945 27571 26979
rect 30757 26945 30791 26979
rect 31401 26945 31435 26979
rect 32137 26945 32171 26979
rect 34529 26945 34563 26979
rect 35909 26945 35943 26979
rect 38853 26945 38887 26979
rect 38945 26945 38979 26979
rect 39589 26945 39623 26979
rect 39682 26945 39716 26979
rect 39957 26945 39991 26979
rect 40054 26945 40088 26979
rect 40877 26945 40911 26979
rect 41061 26945 41095 26979
rect 41153 26945 41187 26979
rect 43637 26945 43671 26979
rect 45845 26945 45879 26979
rect 6377 26877 6411 26911
rect 9321 26877 9355 26911
rect 10701 26877 10735 26911
rect 10885 26877 10919 26911
rect 11989 26877 12023 26911
rect 12081 26877 12115 26911
rect 12449 26877 12483 26911
rect 18061 26877 18095 26911
rect 20545 26877 20579 26911
rect 22937 26877 22971 26911
rect 24961 26877 24995 26911
rect 36001 26877 36035 26911
rect 25881 26809 25915 26843
rect 40233 26809 40267 26843
rect 5825 26741 5859 26775
rect 8401 26741 8435 26775
rect 9781 26741 9815 26775
rect 10241 26741 10275 26775
rect 14289 26741 14323 26775
rect 14841 26741 14875 26775
rect 15577 26741 15611 26775
rect 19901 26741 19935 26775
rect 32321 26741 32355 26775
rect 34713 26741 34747 26775
rect 35265 26741 35299 26775
rect 4813 26537 4847 26571
rect 6009 26537 6043 26571
rect 7389 26537 7423 26571
rect 9045 26537 9079 26571
rect 9965 26537 9999 26571
rect 11069 26537 11103 26571
rect 12265 26537 12299 26571
rect 12817 26537 12851 26571
rect 14749 26537 14783 26571
rect 21005 26537 21039 26571
rect 36737 26537 36771 26571
rect 38209 26537 38243 26571
rect 39313 26537 39347 26571
rect 40785 26537 40819 26571
rect 45109 26537 45143 26571
rect 9137 26469 9171 26503
rect 14565 26469 14599 26503
rect 17969 26469 18003 26503
rect 20821 26469 20855 26503
rect 31677 26469 31711 26503
rect 39865 26469 39899 26503
rect 41613 26469 41647 26503
rect 68017 26469 68051 26503
rect 5273 26401 5307 26435
rect 5457 26401 5491 26435
rect 6837 26401 6871 26435
rect 15393 26401 15427 26435
rect 19257 26401 19291 26435
rect 20545 26401 20579 26435
rect 23489 26401 23523 26435
rect 24961 26401 24995 26435
rect 28917 26401 28951 26435
rect 30113 26401 30147 26435
rect 31217 26401 31251 26435
rect 32229 26401 32263 26435
rect 42993 26401 43027 26435
rect 5181 26333 5215 26367
rect 6193 26333 6227 26367
rect 11897 26333 11931 26367
rect 12725 26333 12759 26367
rect 12909 26333 12943 26367
rect 19533 26333 19567 26367
rect 23673 26333 23707 26367
rect 25237 26333 25271 26367
rect 25697 26333 25731 26367
rect 29009 26333 29043 26367
rect 29561 26333 29595 26367
rect 29929 26333 29963 26367
rect 31309 26333 31343 26367
rect 32321 26333 32355 26367
rect 34713 26333 34747 26367
rect 34969 26333 35003 26367
rect 37933 26333 37967 26367
rect 38669 26333 38703 26367
rect 39037 26333 39071 26367
rect 39129 26333 39163 26367
rect 40049 26333 40083 26367
rect 40325 26333 40359 26367
rect 40969 26333 41003 26367
rect 41153 26333 41187 26367
rect 42726 26333 42760 26367
rect 45201 26333 45235 26367
rect 67833 26333 67867 26367
rect 6929 26265 6963 26299
rect 7021 26265 7055 26299
rect 9505 26265 9539 26299
rect 10609 26265 10643 26299
rect 12081 26265 12115 26299
rect 14289 26265 14323 26299
rect 15669 26265 15703 26299
rect 17417 26265 17451 26299
rect 29653 26265 29687 26299
rect 36645 26265 36679 26299
rect 38025 26265 38059 26299
rect 38209 26265 38243 26299
rect 23857 26197 23891 26231
rect 32689 26197 32723 26231
rect 36093 26197 36127 26231
rect 37381 26197 37415 26231
rect 40233 26197 40267 26231
rect 5733 25993 5767 26027
rect 7297 25993 7331 26027
rect 10609 25993 10643 26027
rect 15945 25993 15979 26027
rect 16957 25993 16991 26027
rect 17417 25993 17451 26027
rect 21925 25993 21959 26027
rect 32137 25993 32171 26027
rect 34713 25993 34747 26027
rect 37933 25993 37967 26027
rect 39497 25993 39531 26027
rect 40601 25993 40635 26027
rect 12633 25925 12667 25959
rect 17325 25925 17359 25959
rect 18245 25925 18279 25959
rect 19533 25925 19567 25959
rect 22753 25925 22787 25959
rect 23397 25925 23431 25959
rect 24593 25925 24627 25959
rect 33250 25925 33284 25959
rect 35081 25925 35115 25959
rect 4905 25857 4939 25891
rect 9229 25857 9263 25891
rect 9496 25857 9530 25891
rect 13369 25857 13403 25891
rect 15393 25857 15427 25891
rect 16129 25857 16163 25891
rect 19073 25857 19107 25891
rect 19717 25857 19751 25891
rect 19809 25857 19843 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 23305 25857 23339 25891
rect 23489 25857 23523 25891
rect 24225 25857 24259 25891
rect 24373 25857 24407 25891
rect 24501 25857 24535 25891
rect 24690 25857 24724 25891
rect 25513 25857 25547 25891
rect 30573 25857 30607 25891
rect 31217 25857 31251 25891
rect 39313 25857 39347 25891
rect 39497 25857 39531 25891
rect 40233 25857 40267 25891
rect 40417 25857 40451 25891
rect 14289 25789 14323 25823
rect 14749 25789 14783 25823
rect 17509 25789 17543 25823
rect 25421 25789 25455 25823
rect 31309 25789 31343 25823
rect 33517 25789 33551 25823
rect 35173 25789 35207 25823
rect 35357 25789 35391 25823
rect 37473 25789 37507 25823
rect 14565 25721 14599 25755
rect 19533 25721 19567 25755
rect 25881 25721 25915 25755
rect 37749 25721 37783 25755
rect 4721 25653 4755 25687
rect 15301 25653 15335 25687
rect 20361 25653 20395 25687
rect 24869 25653 24903 25687
rect 31493 25653 31527 25687
rect 36461 25653 36495 25687
rect 38761 25653 38795 25687
rect 6377 25449 6411 25483
rect 9689 25449 9723 25483
rect 12817 25449 12851 25483
rect 14381 25449 14415 25483
rect 16681 25449 16715 25483
rect 18245 25449 18279 25483
rect 22753 25449 22787 25483
rect 23305 25449 23339 25483
rect 24501 25449 24535 25483
rect 27169 25449 27203 25483
rect 32505 25449 32539 25483
rect 32965 25449 32999 25483
rect 37749 25449 37783 25483
rect 37933 25449 37967 25483
rect 7573 25381 7607 25415
rect 30757 25381 30791 25415
rect 6929 25313 6963 25347
rect 15209 25313 15243 25347
rect 30297 25313 30331 25347
rect 31861 25313 31895 25347
rect 32045 25313 32079 25347
rect 33149 25313 33183 25347
rect 4537 25245 4571 25279
rect 4804 25245 4838 25279
rect 6837 25245 6871 25279
rect 9873 25245 9907 25279
rect 17233 25245 17267 25279
rect 18429 25245 18463 25279
rect 19441 25245 19475 25279
rect 23305 25245 23339 25279
rect 23489 25245 23523 25279
rect 24685 25245 24719 25279
rect 24961 25245 24995 25279
rect 25421 25245 25455 25279
rect 25605 25245 25639 25279
rect 25881 25245 25915 25279
rect 26709 25245 26743 25279
rect 26985 25245 27019 25279
rect 30389 25245 30423 25279
rect 32965 25245 32999 25279
rect 33241 25245 33275 25279
rect 37473 25245 37507 25279
rect 60565 25245 60599 25279
rect 61209 25245 61243 25279
rect 7757 25177 7791 25211
rect 14473 25177 14507 25211
rect 17417 25177 17451 25211
rect 24869 25177 24903 25211
rect 32137 25177 32171 25211
rect 5917 25109 5951 25143
rect 6745 25109 6779 25143
rect 8401 25109 8435 25143
rect 11253 25109 11287 25143
rect 11805 25109 11839 25143
rect 13553 25109 13587 25143
rect 15301 25109 15335 25143
rect 15393 25109 15427 25143
rect 15761 25109 15795 25143
rect 19349 25109 19383 25143
rect 25789 25109 25823 25143
rect 26801 25109 26835 25143
rect 31217 25109 31251 25143
rect 33425 25109 33459 25143
rect 36921 25109 36955 25143
rect 60749 25109 60783 25143
rect 10149 24905 10183 24939
rect 10517 24905 10551 24939
rect 11529 24837 11563 24871
rect 4905 24769 4939 24803
rect 6920 24769 6954 24803
rect 8493 24769 8527 24803
rect 10609 24769 10643 24803
rect 12265 24769 12299 24803
rect 13093 24769 13127 24803
rect 13277 24769 13311 24803
rect 13369 24769 13403 24803
rect 14188 24769 14222 24803
rect 15945 24769 15979 24803
rect 17233 24769 17267 24803
rect 17417 24769 17451 24803
rect 21833 24769 21867 24803
rect 25973 24769 26007 24803
rect 28273 24769 28307 24803
rect 29101 24769 29135 24803
rect 29285 24769 29319 24803
rect 29745 24769 29779 24803
rect 32137 24769 32171 24803
rect 32321 24769 32355 24803
rect 32505 24769 32539 24803
rect 32597 24769 32631 24803
rect 34713 24769 34747 24803
rect 35541 24769 35575 24803
rect 36553 24769 36587 24803
rect 38025 24769 38059 24803
rect 38761 24769 38795 24803
rect 40601 24769 40635 24803
rect 44649 24769 44683 24803
rect 45569 24769 45603 24803
rect 4997 24701 5031 24735
rect 6653 24701 6687 24735
rect 10793 24701 10827 24735
rect 12449 24701 12483 24735
rect 13921 24701 13955 24735
rect 17877 24701 17911 24735
rect 18153 24701 18187 24735
rect 19625 24701 19659 24735
rect 25789 24701 25823 24735
rect 27629 24701 27663 24735
rect 28181 24701 28215 24735
rect 35265 24701 35299 24735
rect 35449 24701 35483 24735
rect 38853 24701 38887 24735
rect 40693 24701 40727 24735
rect 44925 24701 44959 24735
rect 15761 24633 15795 24667
rect 26157 24633 26191 24667
rect 28641 24633 28675 24667
rect 35909 24633 35943 24667
rect 39129 24633 39163 24667
rect 4629 24565 4663 24599
rect 8033 24565 8067 24599
rect 13093 24565 13127 24599
rect 15301 24565 15335 24599
rect 17049 24565 17083 24599
rect 20453 24565 20487 24599
rect 21925 24565 21959 24599
rect 22569 24565 22603 24599
rect 29101 24565 29135 24599
rect 36369 24565 36403 24599
rect 40325 24565 40359 24599
rect 43913 24565 43947 24599
rect 45477 24565 45511 24599
rect 16589 24361 16623 24395
rect 17969 24361 18003 24395
rect 37473 24361 37507 24395
rect 45017 24361 45051 24395
rect 23581 24293 23615 24327
rect 25237 24293 25271 24327
rect 29009 24293 29043 24327
rect 34805 24293 34839 24327
rect 47133 24293 47167 24327
rect 4721 24225 4755 24259
rect 7757 24225 7791 24259
rect 7941 24225 7975 24259
rect 14933 24225 14967 24259
rect 20177 24225 20211 24259
rect 20821 24225 20855 24259
rect 22845 24225 22879 24259
rect 24961 24225 24995 24259
rect 25789 24225 25823 24259
rect 28549 24225 28583 24259
rect 33425 24225 33459 24259
rect 36093 24225 36127 24259
rect 42717 24225 42751 24259
rect 45201 24225 45235 24259
rect 4629 24157 4663 24191
rect 6101 24157 6135 24191
rect 6285 24157 6319 24191
rect 6561 24157 6595 24191
rect 7665 24157 7699 24191
rect 9137 24157 9171 24191
rect 9321 24157 9355 24191
rect 11161 24157 11195 24191
rect 12173 24157 12207 24191
rect 14657 24157 14691 24191
rect 15853 24157 15887 24191
rect 16773 24157 16807 24191
rect 16957 24157 16991 24191
rect 18061 24157 18095 24191
rect 18521 24157 18555 24191
rect 18705 24157 18739 24191
rect 19441 24157 19475 24191
rect 24869 24157 24903 24191
rect 25959 24157 25993 24191
rect 27997 24157 28031 24191
rect 28719 24157 28753 24191
rect 29561 24157 29595 24191
rect 29745 24157 29779 24191
rect 30297 24157 30331 24191
rect 40509 24157 40543 24191
rect 42993 24157 43027 24191
rect 43821 24157 43855 24191
rect 44281 24157 44315 24191
rect 45293 24157 45327 24191
rect 46213 24157 46247 24191
rect 46305 24157 46339 24191
rect 46489 24157 46523 24191
rect 46949 24157 46983 24191
rect 9873 24089 9907 24123
rect 12440 24089 12474 24123
rect 21097 24089 21131 24123
rect 23397 24089 23431 24123
rect 34161 24089 34195 24123
rect 36360 24089 36394 24123
rect 40785 24089 40819 24123
rect 4997 24021 5031 24055
rect 6469 24021 6503 24055
rect 7297 24021 7331 24055
rect 8953 24021 8987 24055
rect 11345 24021 11379 24055
rect 13553 24021 13587 24055
rect 15669 24021 15703 24055
rect 18613 24021 18647 24055
rect 26249 24021 26283 24055
rect 29653 24021 29687 24055
rect 32781 24021 32815 24055
rect 42257 24021 42291 24055
rect 44373 24021 44407 24055
rect 45661 24021 45695 24055
rect 7389 23817 7423 23851
rect 8125 23817 8159 23851
rect 9965 23817 9999 23851
rect 12909 23817 12943 23851
rect 13369 23817 13403 23851
rect 14105 23817 14139 23851
rect 20913 23817 20947 23851
rect 22845 23817 22879 23851
rect 24593 23817 24627 23851
rect 25697 23817 25731 23851
rect 28549 23817 28583 23851
rect 34161 23817 34195 23851
rect 35357 23817 35391 23851
rect 40785 23817 40819 23851
rect 41429 23817 41463 23851
rect 42533 23817 42567 23851
rect 5641 23749 5675 23783
rect 11774 23749 11808 23783
rect 17509 23749 17543 23783
rect 18613 23749 18647 23783
rect 22109 23749 22143 23783
rect 22753 23749 22787 23783
rect 28089 23749 28123 23783
rect 32321 23749 32355 23783
rect 33701 23749 33735 23783
rect 44189 23749 44223 23783
rect 4813 23681 4847 23715
rect 4997 23681 5031 23715
rect 5457 23681 5491 23715
rect 6745 23681 6779 23715
rect 7573 23681 7607 23715
rect 8033 23681 8067 23715
rect 8217 23681 8251 23715
rect 8677 23681 8711 23715
rect 8861 23681 8895 23715
rect 9781 23681 9815 23715
rect 9956 23671 9990 23705
rect 10701 23681 10735 23715
rect 10793 23681 10827 23715
rect 10885 23681 10919 23715
rect 13553 23681 13587 23715
rect 15761 23681 15795 23715
rect 16681 23681 16715 23715
rect 17417 23681 17451 23715
rect 17601 23681 17635 23715
rect 18521 23681 18555 23715
rect 18705 23681 18739 23715
rect 20545 23681 20579 23715
rect 22201 23681 22235 23715
rect 23673 23681 23707 23715
rect 25881 23681 25915 23715
rect 27169 23681 27203 23715
rect 28365 23681 28399 23715
rect 29009 23681 29043 23715
rect 29193 23681 29227 23715
rect 29929 23681 29963 23715
rect 30757 23681 30791 23715
rect 30849 23681 30883 23715
rect 32229 23681 32263 23715
rect 32413 23681 32447 23715
rect 32873 23681 32907 23715
rect 33057 23681 33091 23715
rect 33977 23681 34011 23715
rect 35449 23681 35483 23715
rect 36185 23681 36219 23715
rect 37657 23681 37691 23715
rect 39129 23681 39163 23715
rect 39313 23681 39347 23715
rect 40049 23681 40083 23715
rect 41245 23681 41279 23715
rect 42625 23681 42659 23715
rect 43269 23681 43303 23715
rect 43913 23681 43947 23715
rect 47869 23681 47903 23715
rect 48697 23681 48731 23715
rect 6377 23613 6411 23647
rect 6653 23613 6687 23647
rect 8769 23613 8803 23647
rect 10609 23613 10643 23647
rect 11529 23613 11563 23647
rect 15577 23613 15611 23647
rect 15669 23613 15703 23647
rect 20453 23613 20487 23647
rect 26065 23613 26099 23647
rect 27077 23613 27111 23647
rect 28181 23613 28215 23647
rect 29745 23613 29779 23647
rect 30573 23613 30607 23647
rect 33793 23613 33827 23647
rect 36093 23613 36127 23647
rect 37565 23613 37599 23647
rect 38669 23613 38703 23647
rect 39037 23613 39071 23647
rect 39773 23613 39807 23647
rect 46121 23613 46155 23647
rect 47593 23613 47627 23647
rect 4905 23545 4939 23579
rect 16129 23545 16163 23579
rect 27537 23545 27571 23579
rect 30113 23545 30147 23579
rect 30665 23545 30699 23579
rect 36553 23545 36587 23579
rect 45661 23545 45695 23579
rect 46489 23545 46523 23579
rect 5825 23477 5859 23511
rect 10425 23477 10459 23511
rect 23489 23477 23523 23511
rect 28273 23477 28307 23511
rect 29101 23477 29135 23511
rect 32965 23477 32999 23511
rect 33701 23477 33735 23511
rect 37381 23477 37415 23511
rect 43453 23477 43487 23511
rect 46581 23477 46615 23511
rect 8309 23273 8343 23307
rect 11161 23273 11195 23307
rect 14105 23273 14139 23307
rect 16773 23273 16807 23307
rect 19257 23273 19291 23307
rect 20453 23273 20487 23307
rect 28917 23273 28951 23307
rect 34897 23273 34931 23307
rect 41245 23273 41279 23307
rect 43913 23273 43947 23307
rect 6009 23205 6043 23239
rect 17877 23205 17911 23239
rect 23213 23205 23247 23239
rect 23765 23205 23799 23239
rect 26525 23205 26559 23239
rect 33333 23205 33367 23239
rect 35081 23205 35115 23239
rect 40049 23205 40083 23239
rect 41061 23205 41095 23239
rect 42809 23205 42843 23239
rect 44005 23205 44039 23239
rect 46581 23205 46615 23239
rect 11713 23137 11747 23171
rect 13093 23137 13127 23171
rect 14657 23137 14691 23171
rect 19625 23137 19659 23171
rect 21465 23137 21499 23171
rect 31401 23137 31435 23171
rect 32873 23137 32907 23171
rect 33885 23137 33919 23171
rect 38669 23137 38703 23171
rect 40325 23137 40359 23171
rect 42073 23137 42107 23171
rect 44373 23137 44407 23171
rect 46949 23137 46983 23171
rect 5365 23069 5399 23103
rect 5513 23069 5547 23103
rect 5733 23069 5767 23103
rect 5830 23069 5864 23103
rect 12357 23069 12391 23103
rect 15393 23069 15427 23103
rect 15660 23069 15694 23103
rect 17877 23069 17911 23103
rect 18061 23069 18095 23103
rect 19441 23069 19475 23103
rect 26433 23069 26467 23103
rect 26617 23069 26651 23103
rect 27721 23069 27755 23103
rect 27905 23069 27939 23103
rect 29561 23069 29595 23103
rect 29709 23069 29743 23103
rect 29929 23069 29963 23103
rect 30067 23069 30101 23103
rect 31493 23069 31527 23103
rect 32965 23069 32999 23103
rect 34713 23069 34747 23103
rect 34897 23069 34931 23103
rect 41889 23069 41923 23103
rect 45753 23069 45787 23103
rect 46029 23069 46063 23103
rect 47409 23069 47443 23103
rect 5641 23001 5675 23035
rect 11529 23001 11563 23035
rect 14473 23001 14507 23035
rect 20269 23001 20303 23035
rect 20485 23001 20519 23035
rect 21741 23001 21775 23035
rect 29837 23001 29871 23035
rect 37933 23001 37967 23035
rect 40785 23001 40819 23035
rect 42625 23001 42659 23035
rect 43269 23001 43303 23035
rect 11621 22933 11655 22967
rect 14565 22933 14599 22967
rect 20637 22933 20671 22967
rect 27169 22933 27203 22967
rect 27813 22933 27847 22967
rect 30205 22933 30239 22967
rect 31861 22933 31895 22967
rect 37473 22933 37507 22967
rect 39865 22933 39899 22967
rect 41705 22933 41739 22967
rect 45017 22933 45051 22967
rect 46489 22933 46523 22967
rect 47593 22933 47627 22967
rect 5549 22729 5583 22763
rect 6377 22729 6411 22763
rect 10425 22729 10459 22763
rect 12449 22729 12483 22763
rect 17141 22729 17175 22763
rect 17785 22729 17819 22763
rect 19533 22729 19567 22763
rect 23765 22729 23799 22763
rect 25789 22729 25823 22763
rect 26985 22729 27019 22763
rect 27353 22729 27387 22763
rect 27445 22729 27479 22763
rect 30021 22729 30055 22763
rect 31585 22729 31619 22763
rect 32137 22729 32171 22763
rect 33609 22729 33643 22763
rect 35449 22729 35483 22763
rect 45661 22729 45695 22763
rect 5181 22661 5215 22695
rect 13093 22661 13127 22695
rect 15025 22661 15059 22695
rect 16129 22661 16163 22695
rect 17049 22661 17083 22695
rect 20637 22661 20671 22695
rect 33149 22661 33183 22695
rect 36093 22661 36127 22695
rect 44189 22661 44223 22695
rect 4353 22593 4387 22627
rect 5365 22593 5399 22627
rect 6377 22593 6411 22627
rect 6561 22593 6595 22627
rect 11989 22593 12023 22627
rect 12633 22593 12667 22627
rect 12725 22593 12759 22627
rect 13829 22593 13863 22627
rect 17693 22593 17727 22627
rect 17969 22593 18003 22627
rect 18429 22593 18463 22627
rect 19625 22593 19659 22627
rect 20545 22593 20579 22627
rect 20821 22593 20855 22627
rect 22641 22593 22675 22627
rect 24593 22593 24627 22627
rect 26433 22593 26467 22627
rect 29929 22593 29963 22627
rect 30205 22593 30239 22627
rect 32597 22593 32631 22627
rect 33425 22593 33459 22627
rect 35633 22593 35667 22627
rect 35817 22593 35851 22627
rect 39129 22593 39163 22627
rect 40509 22593 40543 22627
rect 43913 22593 43947 22627
rect 46121 22593 46155 22627
rect 46305 22593 46339 22627
rect 4261 22525 4295 22559
rect 4721 22525 4755 22559
rect 13001 22525 13035 22559
rect 22385 22525 22419 22559
rect 27537 22525 27571 22559
rect 31125 22525 31159 22559
rect 33241 22525 33275 22559
rect 40233 22525 40267 22559
rect 14013 22457 14047 22491
rect 17969 22457 18003 22491
rect 24409 22457 24443 22491
rect 25145 22457 25179 22491
rect 31493 22457 31527 22491
rect 32229 22457 32263 22491
rect 39313 22457 39347 22491
rect 18521 22389 18555 22423
rect 20821 22389 20855 22423
rect 26249 22389 26283 22423
rect 30389 22389 30423 22423
rect 33425 22389 33459 22423
rect 34897 22389 34931 22423
rect 35817 22389 35851 22423
rect 41245 22389 41279 22423
rect 46121 22389 46155 22423
rect 4353 22185 4387 22219
rect 10793 22185 10827 22219
rect 17969 22185 18003 22219
rect 20913 22185 20947 22219
rect 21557 22185 21591 22219
rect 25237 22185 25271 22219
rect 27445 22185 27479 22219
rect 32505 22185 32539 22219
rect 34713 22185 34747 22219
rect 34897 22185 34931 22219
rect 40049 22185 40083 22219
rect 40864 22185 40898 22219
rect 42349 22185 42383 22219
rect 36277 22117 36311 22151
rect 36829 22117 36863 22151
rect 5733 22049 5767 22083
rect 16129 22049 16163 22083
rect 19901 22049 19935 22083
rect 26065 22049 26099 22083
rect 29561 22049 29595 22083
rect 29929 22049 29963 22083
rect 30021 22049 30055 22083
rect 30941 22049 30975 22083
rect 36369 22049 36403 22083
rect 40601 22049 40635 22083
rect 6377 21981 6411 22015
rect 10057 21981 10091 22015
rect 10241 21981 10275 22015
rect 12541 21981 12575 22015
rect 12725 21981 12759 22015
rect 20729 21981 20763 22015
rect 20913 21981 20947 22015
rect 21373 21981 21407 22015
rect 22017 21981 22051 22015
rect 22845 21981 22879 22015
rect 22937 21981 22971 22015
rect 25145 21981 25179 22015
rect 26332 21981 26366 22015
rect 29745 21981 29779 22015
rect 29837 21981 29871 22015
rect 31953 21981 31987 22015
rect 32045 21981 32079 22015
rect 32229 21981 32263 22015
rect 32321 21981 32355 22015
rect 34897 21981 34931 22015
rect 35265 21981 35299 22015
rect 37565 21981 37599 22015
rect 37841 21981 37875 22015
rect 39865 21981 39899 22015
rect 5488 21913 5522 21947
rect 12633 21913 12667 21947
rect 16313 21913 16347 21947
rect 17785 21913 17819 21947
rect 17985 21913 18019 21947
rect 19717 21913 19751 21947
rect 22201 21913 22235 21947
rect 31493 21913 31527 21947
rect 35909 21913 35943 21947
rect 6193 21845 6227 21879
rect 10149 21845 10183 21879
rect 14197 21845 14231 21879
rect 15577 21845 15611 21879
rect 16405 21845 16439 21879
rect 16773 21845 16807 21879
rect 18153 21845 18187 21879
rect 18613 21845 18647 21879
rect 24593 21845 24627 21879
rect 25605 21845 25639 21879
rect 34069 21845 34103 21879
rect 37381 21845 37415 21879
rect 37749 21845 37783 21879
rect 5457 21641 5491 21675
rect 5825 21641 5859 21675
rect 8033 21641 8067 21675
rect 10977 21641 11011 21675
rect 20913 21641 20947 21675
rect 21281 21641 21315 21675
rect 24593 21641 24627 21675
rect 26433 21641 26467 21675
rect 30113 21641 30147 21675
rect 11774 21573 11808 21607
rect 22753 21573 22787 21607
rect 34713 21573 34747 21607
rect 35541 21573 35575 21607
rect 7113 21505 7147 21539
rect 7941 21505 7975 21539
rect 8217 21505 8251 21539
rect 9137 21505 9171 21539
rect 10057 21505 10091 21539
rect 10241 21505 10275 21539
rect 10793 21505 10827 21539
rect 11529 21505 11563 21539
rect 13369 21505 13403 21539
rect 14197 21505 14231 21539
rect 15117 21505 15151 21539
rect 16681 21505 16715 21539
rect 17509 21505 17543 21539
rect 22937 21505 22971 21539
rect 24133 21505 24167 21539
rect 26157 21505 26191 21539
rect 26249 21505 26283 21539
rect 28825 21505 28859 21539
rect 29653 21505 29687 21539
rect 29745 21505 29779 21539
rect 29929 21505 29963 21539
rect 30573 21505 30607 21539
rect 30757 21505 30791 21539
rect 32321 21505 32355 21539
rect 32413 21505 32447 21539
rect 36553 21505 36587 21539
rect 36737 21505 36771 21539
rect 37289 21505 37323 21539
rect 38025 21505 38059 21539
rect 44281 21505 44315 21539
rect 45753 21505 45787 21539
rect 46029 21505 46063 21539
rect 46857 21505 46891 21539
rect 5273 21437 5307 21471
rect 5365 21437 5399 21471
rect 6377 21437 6411 21471
rect 7205 21437 7239 21471
rect 8953 21437 8987 21471
rect 13921 21437 13955 21471
rect 17785 21437 17819 21471
rect 20729 21437 20763 21471
rect 20821 21437 20855 21471
rect 25789 21437 25823 21471
rect 32689 21437 32723 21471
rect 32781 21437 32815 21471
rect 35265 21437 35299 21471
rect 35449 21437 35483 21471
rect 37933 21437 37967 21471
rect 44097 21437 44131 21471
rect 9321 21369 9355 21403
rect 12909 21369 12943 21403
rect 28457 21369 28491 21403
rect 32137 21369 32171 21403
rect 33333 21369 33367 21403
rect 7389 21301 7423 21335
rect 8401 21301 8435 21335
rect 10149 21301 10183 21335
rect 14933 21301 14967 21335
rect 16865 21301 16899 21335
rect 19257 21301 19291 21335
rect 19901 21301 19935 21335
rect 21833 21301 21867 21335
rect 24409 21301 24443 21335
rect 25053 21301 25087 21335
rect 27813 21301 27847 21335
rect 28365 21301 28399 21335
rect 30665 21301 30699 21335
rect 35909 21301 35943 21335
rect 36737 21301 36771 21335
rect 38301 21301 38335 21335
rect 44465 21301 44499 21335
rect 10517 21097 10551 21131
rect 11437 21097 11471 21131
rect 16589 21097 16623 21131
rect 18429 21097 18463 21131
rect 23581 21097 23615 21131
rect 25697 21097 25731 21131
rect 28457 21097 28491 21131
rect 30849 21097 30883 21131
rect 32137 21097 32171 21131
rect 35725 21097 35759 21131
rect 39957 21097 39991 21131
rect 41797 21097 41831 21131
rect 25053 21029 25087 21063
rect 27905 21029 27939 21063
rect 28825 21029 28859 21063
rect 29837 21029 29871 21063
rect 35633 21029 35667 21063
rect 36185 21029 36219 21063
rect 40325 21029 40359 21063
rect 6561 20961 6595 20995
rect 7481 20961 7515 20995
rect 7573 20961 7607 20995
rect 10885 20961 10919 20995
rect 11897 20961 11931 20995
rect 12081 20961 12115 20995
rect 14473 20961 14507 20995
rect 19257 20961 19291 20995
rect 19533 20961 19567 20995
rect 20545 20961 20579 20995
rect 30021 20961 30055 20995
rect 33517 20961 33551 20995
rect 34805 20961 34839 20995
rect 35265 20961 35299 20995
rect 38301 20961 38335 20995
rect 39957 20961 39991 20995
rect 9275 20893 9309 20927
rect 9413 20893 9447 20927
rect 9633 20893 9667 20927
rect 9781 20893 9815 20927
rect 10793 20893 10827 20927
rect 11805 20893 11839 20927
rect 14740 20893 14774 20927
rect 17702 20893 17736 20927
rect 17969 20893 18003 20927
rect 18613 20893 18647 20927
rect 20821 20893 20855 20927
rect 22201 20893 22235 20927
rect 25881 20893 25915 20927
rect 25973 20893 26007 20927
rect 27629 20893 27663 20927
rect 28365 20893 28399 20927
rect 30481 20893 30515 20927
rect 30665 20893 30699 20927
rect 32045 20893 32079 20927
rect 32229 20893 32263 20927
rect 32689 20893 32723 20927
rect 37565 20893 37599 20927
rect 38393 20893 38427 20927
rect 39865 20893 39899 20927
rect 40141 20893 40175 20927
rect 41889 20893 41923 20927
rect 42533 20893 42567 20927
rect 42717 20893 42751 20927
rect 43177 20893 43211 20927
rect 43453 20893 43487 20927
rect 45017 20893 45051 20927
rect 45661 20893 45695 20927
rect 6294 20825 6328 20859
rect 7389 20825 7423 20859
rect 9505 20825 9539 20859
rect 22468 20825 22502 20859
rect 24777 20825 24811 20859
rect 25697 20825 25731 20859
rect 27905 20825 27939 20859
rect 29561 20825 29595 20859
rect 37298 20825 37332 20859
rect 42625 20825 42659 20859
rect 5181 20757 5215 20791
rect 7021 20757 7055 20791
rect 9137 20757 9171 20791
rect 12725 20757 12759 20791
rect 15853 20757 15887 20791
rect 25237 20757 25271 20791
rect 26433 20757 26467 20791
rect 27721 20757 27755 20791
rect 38025 20757 38059 20791
rect 40969 20757 41003 20791
rect 44189 20757 44223 20791
rect 45201 20757 45235 20791
rect 45845 20757 45879 20791
rect 6377 20553 6411 20587
rect 9413 20553 9447 20587
rect 11529 20553 11563 20587
rect 17141 20553 17175 20587
rect 21189 20553 21223 20587
rect 22661 20553 22695 20587
rect 22753 20553 22787 20587
rect 25973 20553 26007 20587
rect 28273 20553 28307 20587
rect 29377 20553 29411 20587
rect 30021 20553 30055 20587
rect 32873 20553 32907 20587
rect 33977 20553 34011 20587
rect 36461 20553 36495 20587
rect 40601 20553 40635 20587
rect 41245 20553 41279 20587
rect 41337 20553 41371 20587
rect 42533 20553 42567 20587
rect 14381 20485 14415 20519
rect 15669 20485 15703 20519
rect 18061 20485 18095 20519
rect 18705 20485 18739 20519
rect 20453 20485 20487 20519
rect 32689 20485 32723 20519
rect 34682 20485 34716 20519
rect 37657 20485 37691 20519
rect 38117 20485 38151 20519
rect 41797 20485 41831 20519
rect 43913 20485 43947 20519
rect 6561 20417 6595 20451
rect 7481 20417 7515 20451
rect 8953 20417 8987 20451
rect 9045 20417 9079 20451
rect 9229 20417 9263 20451
rect 10333 20417 10367 20451
rect 10977 20417 11011 20451
rect 14473 20417 14507 20451
rect 17049 20417 17083 20451
rect 17969 20417 18003 20451
rect 18613 20417 18647 20451
rect 18981 20417 19015 20451
rect 19717 20417 19751 20451
rect 19901 20417 19935 20451
rect 24593 20417 24627 20451
rect 25513 20417 25547 20451
rect 27905 20417 27939 20451
rect 29745 20417 29779 20451
rect 32505 20417 32539 20451
rect 33793 20417 33827 20451
rect 36277 20417 36311 20451
rect 40049 20417 40083 20451
rect 40141 20417 40175 20451
rect 40325 20417 40359 20451
rect 40417 20417 40451 20451
rect 42441 20417 42475 20451
rect 42717 20417 42751 20451
rect 45845 20417 45879 20451
rect 46121 20417 46155 20451
rect 7389 20349 7423 20383
rect 9873 20349 9907 20383
rect 12081 20349 12115 20383
rect 14289 20349 14323 20383
rect 15761 20349 15795 20383
rect 15853 20349 15887 20383
rect 17233 20349 17267 20383
rect 19073 20349 19107 20383
rect 22845 20349 22879 20383
rect 25053 20349 25087 20383
rect 27813 20349 27847 20383
rect 29837 20349 29871 20383
rect 34437 20349 34471 20383
rect 38945 20349 38979 20383
rect 43637 20349 43671 20383
rect 45385 20349 45419 20383
rect 7849 20281 7883 20315
rect 15301 20281 15335 20315
rect 41797 20281 41831 20315
rect 5549 20213 5583 20247
rect 10241 20213 10275 20247
rect 10793 20213 10827 20247
rect 14841 20213 14875 20247
rect 16681 20213 16715 20247
rect 19257 20213 19291 20247
rect 19717 20213 19751 20247
rect 22293 20213 22327 20247
rect 24041 20213 24075 20247
rect 24777 20213 24811 20247
rect 25789 20213 25823 20247
rect 28733 20213 28767 20247
rect 35817 20213 35851 20247
rect 41061 20213 41095 20247
rect 42901 20213 42935 20247
rect 46857 20213 46891 20247
rect 6193 20009 6227 20043
rect 7665 20009 7699 20043
rect 11989 20009 12023 20043
rect 22477 20009 22511 20043
rect 23305 20009 23339 20043
rect 27353 20009 27387 20043
rect 31769 20009 31803 20043
rect 34897 20009 34931 20043
rect 40049 20009 40083 20043
rect 41429 20009 41463 20043
rect 41613 20009 41647 20043
rect 45477 20009 45511 20043
rect 14197 19941 14231 19975
rect 16681 19941 16715 19975
rect 17141 19941 17175 19975
rect 18061 19941 18095 19975
rect 21189 19941 21223 19975
rect 26065 19941 26099 19975
rect 30481 19941 30515 19975
rect 37841 19941 37875 19975
rect 45293 19941 45327 19975
rect 5089 19873 5123 19907
rect 8953 19873 8987 19907
rect 12541 19873 12575 19907
rect 15301 19873 15335 19907
rect 19625 19873 19659 19907
rect 25789 19873 25823 19907
rect 27169 19873 27203 19907
rect 30021 19873 30055 19907
rect 32137 19873 32171 19907
rect 35449 19873 35483 19907
rect 37565 19873 37599 19907
rect 40233 19873 40267 19907
rect 42809 19873 42843 19907
rect 45017 19873 45051 19907
rect 4997 19805 5031 19839
rect 6101 19805 6135 19839
rect 7849 19805 7883 19839
rect 8033 19805 8067 19839
rect 8125 19805 8159 19839
rect 9137 19805 9171 19839
rect 10149 19805 10183 19839
rect 12449 19805 12483 19839
rect 14841 19805 14875 19839
rect 18521 19805 18555 19839
rect 18705 19805 18739 19839
rect 19717 19805 19751 19839
rect 20085 19805 20119 19839
rect 20545 19805 20579 19839
rect 20729 19805 20763 19839
rect 22293 19805 22327 19839
rect 23121 19805 23155 19839
rect 25697 19805 25731 19839
rect 27077 19805 27111 19839
rect 30113 19805 30147 19839
rect 31677 19805 31711 19839
rect 32781 19805 32815 19839
rect 35357 19805 35391 19839
rect 37473 19805 37507 19839
rect 40325 19805 40359 19839
rect 43085 19805 43119 19839
rect 10416 19737 10450 19771
rect 15568 19737 15602 19771
rect 19993 19737 20027 19771
rect 34161 19737 34195 19771
rect 35265 19737 35299 19771
rect 40601 19737 40635 19771
rect 40693 19737 40727 19771
rect 41245 19737 41279 19771
rect 41461 19737 41495 19771
rect 5365 19669 5399 19703
rect 6561 19669 6595 19703
rect 7113 19669 7147 19703
rect 9321 19669 9355 19703
rect 11529 19669 11563 19703
rect 12357 19669 12391 19703
rect 14657 19669 14691 19703
rect 18705 19669 18739 19703
rect 19441 19669 19475 19703
rect 20637 19669 20671 19703
rect 31125 19669 31159 19703
rect 32597 19669 32631 19703
rect 43821 19669 43855 19703
rect 3893 19465 3927 19499
rect 5733 19465 5767 19499
rect 6837 19465 6871 19499
rect 15485 19465 15519 19499
rect 15945 19465 15979 19499
rect 31585 19465 31619 19499
rect 33609 19465 33643 19499
rect 40877 19465 40911 19499
rect 45109 19465 45143 19499
rect 4598 19397 4632 19431
rect 6377 19397 6411 19431
rect 7573 19397 7607 19431
rect 14372 19397 14406 19431
rect 20913 19397 20947 19431
rect 22477 19397 22511 19431
rect 43637 19397 43671 19431
rect 3709 19329 3743 19363
rect 4353 19329 4387 19363
rect 7297 19329 7331 19363
rect 7389 19329 7423 19363
rect 10517 19329 10551 19363
rect 14105 19329 14139 19363
rect 16129 19329 16163 19363
rect 18797 19329 18831 19363
rect 19533 19329 19567 19363
rect 19625 19329 19659 19363
rect 19809 19329 19843 19363
rect 19901 19329 19935 19363
rect 21833 19329 21867 19363
rect 23397 19329 23431 19363
rect 24409 19329 24443 19363
rect 24676 19329 24710 19363
rect 31401 19329 31435 19363
rect 32229 19329 32263 19363
rect 32496 19329 32530 19363
rect 39681 19329 39715 19363
rect 40509 19329 40543 19363
rect 40693 19329 40727 19363
rect 43361 19329 43395 19363
rect 9689 19261 9723 19295
rect 10609 19261 10643 19295
rect 11621 19261 11655 19295
rect 16773 19261 16807 19295
rect 19073 19261 19107 19295
rect 21005 19261 21039 19295
rect 21097 19261 21131 19295
rect 23121 19261 23155 19295
rect 39773 19261 39807 19295
rect 40049 19261 40083 19295
rect 6653 19193 6687 19227
rect 7573 19193 7607 19227
rect 22661 19193 22695 19227
rect 18889 19125 18923 19159
rect 18981 19125 19015 19159
rect 20085 19125 20119 19159
rect 20545 19125 20579 19159
rect 25789 19125 25823 19159
rect 26249 19125 26283 19159
rect 34805 19125 34839 19159
rect 4997 18921 5031 18955
rect 17877 18921 17911 18955
rect 19349 18921 19383 18955
rect 23581 18921 23615 18955
rect 24685 18921 24719 18955
rect 28641 18921 28675 18955
rect 29009 18921 29043 18955
rect 32873 18921 32907 18955
rect 33333 18921 33367 18955
rect 40233 18921 40267 18955
rect 44281 18921 44315 18955
rect 45109 18921 45143 18955
rect 10609 18853 10643 18887
rect 12633 18853 12667 18887
rect 25329 18853 25363 18887
rect 26985 18853 27019 18887
rect 28089 18853 28123 18887
rect 5641 18785 5675 18819
rect 7021 18785 7055 18819
rect 19533 18785 19567 18819
rect 25789 18785 25823 18819
rect 25973 18785 26007 18819
rect 27813 18785 27847 18819
rect 33793 18785 33827 18819
rect 33885 18785 33919 18819
rect 39313 18785 39347 18819
rect 5365 18717 5399 18751
rect 11805 18717 11839 18751
rect 16957 18717 16991 18751
rect 17785 18717 17819 18751
rect 19257 18717 19291 18751
rect 20545 18717 20579 18751
rect 21189 18717 21223 18751
rect 24869 18717 24903 18751
rect 27721 18717 27755 18751
rect 28549 18717 28583 18751
rect 31493 18717 31527 18751
rect 40141 18717 40175 18751
rect 40325 18717 40359 18751
rect 44189 18717 44223 18751
rect 45017 18717 45051 18751
rect 67833 18717 67867 18751
rect 10793 18649 10827 18683
rect 12265 18649 12299 18683
rect 21434 18649 21468 18683
rect 23305 18649 23339 18683
rect 29561 18649 29595 18683
rect 31760 18649 31794 18683
rect 33701 18649 33735 18683
rect 39046 18649 39080 18683
rect 5457 18581 5491 18615
rect 6285 18581 6319 18615
rect 7757 18581 7791 18615
rect 11621 18581 11655 18615
rect 12725 18581 12759 18615
rect 13277 18581 13311 18615
rect 17141 18581 17175 18615
rect 19809 18581 19843 18615
rect 20729 18581 20763 18615
rect 22569 18581 22603 18615
rect 25697 18581 25731 18615
rect 37933 18581 37967 18615
rect 68017 18581 68051 18615
rect 7205 18377 7239 18411
rect 8493 18377 8527 18411
rect 15761 18377 15795 18411
rect 18429 18377 18463 18411
rect 19257 18377 19291 18411
rect 19901 18377 19935 18411
rect 22845 18377 22879 18411
rect 25329 18377 25363 18411
rect 29193 18377 29227 18411
rect 32137 18377 32171 18411
rect 32597 18377 32631 18411
rect 33701 18377 33735 18411
rect 37933 18377 37967 18411
rect 38025 18377 38059 18411
rect 38393 18377 38427 18411
rect 38853 18377 38887 18411
rect 11774 18309 11808 18343
rect 7665 18241 7699 18275
rect 8309 18241 8343 18275
rect 11529 18241 11563 18275
rect 15669 18241 15703 18275
rect 17305 18241 17339 18275
rect 19073 18241 19107 18275
rect 19349 18241 19383 18275
rect 20453 18241 20487 18275
rect 23949 18241 23983 18275
rect 24961 18241 24995 18275
rect 29377 18241 29411 18275
rect 30757 18241 30791 18275
rect 31217 18241 31251 18275
rect 32505 18241 32539 18275
rect 33793 18241 33827 18275
rect 34529 18241 34563 18275
rect 39037 18241 39071 18275
rect 8125 18173 8159 18207
rect 13829 18173 13863 18207
rect 15945 18173 15979 18207
rect 17049 18173 17083 18207
rect 25053 18173 25087 18207
rect 26985 18173 27019 18207
rect 31585 18173 31619 18207
rect 32689 18173 32723 18207
rect 37841 18173 37875 18207
rect 13369 18105 13403 18139
rect 13553 18105 13587 18139
rect 14381 18105 14415 18139
rect 22293 18105 22327 18139
rect 24409 18105 24443 18139
rect 7481 18037 7515 18071
rect 12909 18037 12943 18071
rect 15301 18037 15335 18071
rect 18889 18037 18923 18071
rect 20683 18037 20717 18071
rect 23397 18037 23431 18071
rect 24961 18037 24995 18071
rect 25881 18037 25915 18071
rect 34713 18037 34747 18071
rect 43545 18037 43579 18071
rect 11989 17833 12023 17867
rect 16405 17833 16439 17867
rect 17049 17833 17083 17867
rect 26157 17833 26191 17867
rect 33517 17833 33551 17867
rect 36829 17833 36863 17867
rect 19901 17765 19935 17799
rect 23029 17765 23063 17799
rect 27353 17765 27387 17799
rect 31493 17765 31527 17799
rect 5457 17697 5491 17731
rect 7297 17697 7331 17731
rect 7665 17697 7699 17731
rect 12541 17697 12575 17731
rect 17601 17697 17635 17731
rect 32413 17697 32447 17731
rect 32597 17697 32631 17731
rect 44281 17697 44315 17731
rect 5365 17629 5399 17663
rect 7757 17629 7791 17663
rect 11069 17629 11103 17663
rect 11345 17629 11379 17663
rect 12357 17629 12391 17663
rect 15025 17629 15059 17663
rect 17417 17629 17451 17663
rect 19717 17629 19751 17663
rect 20637 17629 20671 17663
rect 20821 17629 20855 17663
rect 21281 17629 21315 17663
rect 23673 17629 23707 17663
rect 24869 17629 24903 17663
rect 30113 17629 30147 17663
rect 35826 17629 35860 17663
rect 36093 17629 36127 17663
rect 37565 17629 37599 17663
rect 40049 17629 40083 17663
rect 43085 17629 43119 17663
rect 55321 17629 55355 17663
rect 55965 17629 55999 17663
rect 13277 17561 13311 17595
rect 13461 17561 13495 17595
rect 15292 17561 15326 17595
rect 20729 17561 20763 17595
rect 21557 17561 21591 17595
rect 27169 17561 27203 17595
rect 30380 17561 30414 17595
rect 32321 17561 32355 17595
rect 36737 17561 36771 17595
rect 37810 17561 37844 17595
rect 44097 17561 44131 17595
rect 5733 17493 5767 17527
rect 7941 17493 7975 17527
rect 11161 17493 11195 17527
rect 11529 17493 11563 17527
rect 12449 17493 12483 17527
rect 14197 17493 14231 17527
rect 17509 17493 17543 17527
rect 18245 17493 18279 17527
rect 23489 17493 23523 17527
rect 31953 17493 31987 17527
rect 34713 17493 34747 17527
rect 38945 17493 38979 17527
rect 39865 17493 39899 17527
rect 42073 17493 42107 17527
rect 43269 17493 43303 17527
rect 43729 17493 43763 17527
rect 44189 17493 44223 17527
rect 55505 17493 55539 17527
rect 4629 17289 4663 17323
rect 5089 17289 5123 17323
rect 6469 17289 6503 17323
rect 7665 17289 7699 17323
rect 15209 17289 15243 17323
rect 20085 17289 20119 17323
rect 21925 17289 21959 17323
rect 22569 17289 22603 17323
rect 24409 17289 24443 17323
rect 27905 17289 27939 17323
rect 34897 17289 34931 17323
rect 35541 17289 35575 17323
rect 37473 17289 37507 17323
rect 13277 17221 13311 17255
rect 19901 17221 19935 17255
rect 26188 17221 26222 17255
rect 32597 17221 32631 17255
rect 43882 17221 43916 17255
rect 3985 17153 4019 17187
rect 4997 17153 5031 17187
rect 7297 17153 7331 17187
rect 8125 17153 8159 17187
rect 10793 17153 10827 17187
rect 11897 17153 11931 17187
rect 12541 17153 12575 17187
rect 12725 17153 12759 17187
rect 15393 17153 15427 17187
rect 16865 17153 16899 17187
rect 18797 17153 18831 17187
rect 18981 17153 19015 17187
rect 19257 17153 19291 17187
rect 20177 17153 20211 17187
rect 20821 17153 20855 17187
rect 21005 17153 21039 17187
rect 21097 17153 21131 17187
rect 21833 17153 21867 17187
rect 22017 17153 22051 17187
rect 22661 17153 22695 17187
rect 23121 17153 23155 17187
rect 23305 17153 23339 17187
rect 24225 17153 24259 17187
rect 26985 17153 27019 17187
rect 28089 17153 28123 17187
rect 30941 17153 30975 17187
rect 33701 17153 33735 17187
rect 34529 17153 34563 17187
rect 35449 17153 35483 17187
rect 37289 17153 37323 17187
rect 37933 17153 37967 17187
rect 38200 17153 38234 17187
rect 41613 17153 41647 17187
rect 42625 17153 42659 17187
rect 43637 17153 43671 17187
rect 45661 17153 45695 17187
rect 5273 17085 5307 17119
rect 7389 17085 7423 17119
rect 10701 17085 10735 17119
rect 11805 17085 11839 17119
rect 17693 17085 17727 17119
rect 24593 17085 24627 17119
rect 26433 17085 26467 17119
rect 27077 17085 27111 17119
rect 28549 17085 28583 17119
rect 34253 17085 34287 17119
rect 34437 17085 34471 17119
rect 42533 17085 42567 17119
rect 45569 17085 45603 17119
rect 12541 17017 12575 17051
rect 17969 17017 18003 17051
rect 19441 17017 19475 17051
rect 23489 17017 23523 17051
rect 25053 17017 25087 17051
rect 30757 17017 30791 17051
rect 46029 17017 46063 17051
rect 4169 16949 4203 16983
rect 10517 16949 10551 16983
rect 11621 16949 11655 16983
rect 16681 16949 16715 16983
rect 18153 16949 18187 16983
rect 19901 16949 19935 16983
rect 23121 16949 23155 16983
rect 24041 16949 24075 16983
rect 26985 16949 27019 16983
rect 27353 16949 27387 16983
rect 32689 16949 32723 16983
rect 36461 16949 36495 16983
rect 39313 16949 39347 16983
rect 41797 16949 41831 16983
rect 42901 16949 42935 16983
rect 45017 16949 45051 16983
rect 5733 16745 5767 16779
rect 7297 16745 7331 16779
rect 8953 16745 8987 16779
rect 11529 16745 11563 16779
rect 12633 16745 12667 16779
rect 19257 16745 19291 16779
rect 23397 16745 23431 16779
rect 37289 16745 37323 16779
rect 42441 16745 42475 16779
rect 43269 16745 43303 16779
rect 17969 16677 18003 16711
rect 18153 16677 18187 16711
rect 20913 16677 20947 16711
rect 31861 16677 31895 16711
rect 34713 16677 34747 16711
rect 40417 16677 40451 16711
rect 41429 16677 41463 16711
rect 41889 16677 41923 16711
rect 45201 16677 45235 16711
rect 46029 16677 46063 16711
rect 4353 16609 4387 16643
rect 6929 16609 6963 16643
rect 8125 16609 8159 16643
rect 9045 16609 9079 16643
rect 11621 16609 11655 16643
rect 19349 16609 19383 16643
rect 22201 16609 22235 16643
rect 23305 16609 23339 16643
rect 25145 16609 25179 16643
rect 27537 16609 27571 16643
rect 30941 16609 30975 16643
rect 33517 16609 33551 16643
rect 33701 16609 33735 16643
rect 36093 16609 36127 16643
rect 37749 16609 37783 16643
rect 37933 16609 37967 16643
rect 38577 16609 38611 16643
rect 38761 16609 38795 16643
rect 40141 16609 40175 16643
rect 40969 16609 41003 16643
rect 43729 16609 43763 16643
rect 43821 16609 43855 16643
rect 45109 16609 45143 16643
rect 45293 16609 45327 16643
rect 45569 16609 45603 16643
rect 7021 16541 7055 16575
rect 8217 16541 8251 16575
rect 9229 16541 9263 16575
rect 11529 16541 11563 16575
rect 11805 16541 11839 16575
rect 15853 16541 15887 16575
rect 19533 16541 19567 16575
rect 21925 16541 21959 16575
rect 23581 16541 23615 16575
rect 24869 16541 24903 16575
rect 28181 16541 28215 16575
rect 28825 16541 28859 16575
rect 32321 16541 32355 16575
rect 33793 16541 33827 16575
rect 40049 16541 40083 16575
rect 41061 16541 41095 16575
rect 42073 16541 42107 16575
rect 42165 16541 42199 16575
rect 45385 16541 45419 16575
rect 46029 16541 46063 16575
rect 46213 16541 46247 16575
rect 46305 16541 46339 16575
rect 4620 16473 4654 16507
rect 8953 16473 8987 16507
rect 16120 16473 16154 16507
rect 17693 16473 17727 16507
rect 19257 16473 19291 16507
rect 27292 16473 27326 16507
rect 30674 16473 30708 16507
rect 35826 16473 35860 16507
rect 43637 16473 43671 16507
rect 45201 16473 45235 16507
rect 7849 16405 7883 16439
rect 9413 16405 9447 16439
rect 11989 16405 12023 16439
rect 17233 16405 17267 16439
rect 19717 16405 19751 16439
rect 23029 16405 23063 16439
rect 26157 16405 26191 16439
rect 27997 16405 28031 16439
rect 29009 16405 29043 16439
rect 29561 16405 29595 16439
rect 32505 16405 32539 16439
rect 34161 16405 34195 16439
rect 36737 16405 36771 16439
rect 37657 16405 37691 16439
rect 38853 16405 38887 16439
rect 39221 16405 39255 16439
rect 42257 16405 42291 16439
rect 5825 16201 5859 16235
rect 6745 16201 6779 16235
rect 8125 16201 8159 16235
rect 10977 16201 11011 16235
rect 14841 16201 14875 16235
rect 15761 16201 15795 16235
rect 18797 16201 18831 16235
rect 22201 16201 22235 16235
rect 22753 16201 22787 16235
rect 24685 16201 24719 16235
rect 27261 16201 27295 16235
rect 27721 16201 27755 16235
rect 29469 16201 29503 16235
rect 29929 16201 29963 16235
rect 32321 16201 32355 16235
rect 33977 16201 34011 16235
rect 42717 16201 42751 16235
rect 43453 16201 43487 16235
rect 45293 16201 45327 16235
rect 11989 16133 12023 16167
rect 12817 16133 12851 16167
rect 13369 16133 13403 16167
rect 17325 16133 17359 16167
rect 23305 16133 23339 16167
rect 31585 16133 31619 16167
rect 32689 16133 32723 16167
rect 44158 16133 44192 16167
rect 4445 16065 4479 16099
rect 4712 16065 4746 16099
rect 7757 16065 7791 16099
rect 10609 16065 10643 16099
rect 15669 16065 15703 16099
rect 24777 16065 24811 16099
rect 25605 16065 25639 16099
rect 27353 16065 27387 16099
rect 28181 16065 28215 16099
rect 29837 16065 29871 16099
rect 33793 16065 33827 16099
rect 34805 16065 34839 16099
rect 43269 16065 43303 16099
rect 6837 15997 6871 16031
rect 6929 15997 6963 16031
rect 7849 15997 7883 16031
rect 10517 15997 10551 16031
rect 15945 15997 15979 16031
rect 18153 15997 18187 16031
rect 23489 15997 23523 16031
rect 24501 15997 24535 16031
rect 27077 15997 27111 16031
rect 30113 15997 30147 16031
rect 32781 15997 32815 16031
rect 32873 15997 32907 16031
rect 34713 15997 34747 16031
rect 43913 15997 43947 16031
rect 6377 15929 6411 15963
rect 25145 15929 25179 15963
rect 8585 15861 8619 15895
rect 14197 15861 14231 15895
rect 15301 15861 15335 15895
rect 28273 15861 28307 15895
rect 28917 15861 28951 15895
rect 34437 15861 34471 15895
rect 5181 15657 5215 15691
rect 7205 15657 7239 15691
rect 16681 15657 16715 15691
rect 21833 15657 21867 15691
rect 28181 15657 28215 15691
rect 39221 15657 39255 15691
rect 42349 15657 42383 15691
rect 9505 15589 9539 15623
rect 40233 15589 40267 15623
rect 41797 15589 41831 15623
rect 42993 15589 43027 15623
rect 44465 15589 44499 15623
rect 5825 15521 5859 15555
rect 7665 15521 7699 15555
rect 10885 15521 10919 15555
rect 14749 15521 14783 15555
rect 17233 15521 17267 15555
rect 26709 15521 26743 15555
rect 28089 15521 28123 15555
rect 29837 15521 29871 15555
rect 41429 15521 41463 15555
rect 44005 15521 44039 15555
rect 5365 15453 5399 15487
rect 10609 15453 10643 15487
rect 12817 15453 12851 15487
rect 14105 15453 14139 15487
rect 17049 15453 17083 15487
rect 22293 15453 22327 15487
rect 22477 15453 22511 15487
rect 23673 15453 23707 15487
rect 26801 15453 26835 15487
rect 28365 15453 28399 15487
rect 29929 15453 29963 15487
rect 32137 15453 32171 15487
rect 41507 15453 41541 15487
rect 42993 15453 43027 15487
rect 43269 15453 43303 15487
rect 44097 15453 44131 15487
rect 6092 15385 6126 15419
rect 7849 15385 7883 15419
rect 9689 15385 9723 15419
rect 12550 15385 12584 15419
rect 14994 15385 15028 15419
rect 17141 15385 17175 15419
rect 17877 15385 17911 15419
rect 24685 15385 24719 15419
rect 32404 15385 32438 15419
rect 39865 15385 39899 15419
rect 10241 15317 10275 15351
rect 10701 15317 10735 15351
rect 11437 15317 11471 15351
rect 14289 15317 14323 15351
rect 16129 15317 16163 15351
rect 19349 15317 19383 15351
rect 22385 15317 22419 15351
rect 22937 15317 22971 15351
rect 23765 15317 23799 15351
rect 26065 15317 26099 15351
rect 27169 15317 27203 15351
rect 28549 15317 28583 15351
rect 29561 15317 29595 15351
rect 33517 15317 33551 15351
rect 40325 15317 40359 15351
rect 43177 15317 43211 15351
rect 7021 15113 7055 15147
rect 10609 15113 10643 15147
rect 11621 15113 11655 15147
rect 12541 15113 12575 15147
rect 13185 15113 13219 15147
rect 20545 15113 20579 15147
rect 22201 15113 22235 15147
rect 24409 15113 24443 15147
rect 24869 15113 24903 15147
rect 27261 15113 27295 15147
rect 27905 15113 27939 15147
rect 34161 15113 34195 15147
rect 38853 15113 38887 15147
rect 39773 15113 39807 15147
rect 40877 15113 40911 15147
rect 13645 15045 13679 15079
rect 17049 15045 17083 15079
rect 21833 15045 21867 15079
rect 22033 15045 22067 15079
rect 22937 15045 22971 15079
rect 34345 15045 34379 15079
rect 40049 15045 40083 15079
rect 40141 15045 40175 15079
rect 42901 15045 42935 15079
rect 43269 15045 43303 15079
rect 9229 14977 9263 15011
rect 9496 14977 9530 15011
rect 12357 14977 12391 15011
rect 13553 14977 13587 15011
rect 14381 14977 14415 15011
rect 14565 14977 14599 15011
rect 15485 14977 15519 15011
rect 17233 14977 17267 15011
rect 18420 14977 18454 15011
rect 20269 14977 20303 15011
rect 21097 14977 21131 15011
rect 22661 14977 22695 15011
rect 25982 14977 26016 15011
rect 26249 14977 26283 15011
rect 27169 14977 27203 15011
rect 28084 14977 28118 15011
rect 28181 14977 28215 15011
rect 28273 14977 28307 15011
rect 28456 14977 28490 15011
rect 28549 14977 28583 15011
rect 29469 14977 29503 15011
rect 30481 14977 30515 15011
rect 32597 14977 32631 15011
rect 32781 14977 32815 15011
rect 33149 14977 33183 15011
rect 33241 14977 33275 15011
rect 33609 14977 33643 15011
rect 34069 14977 34103 15011
rect 39911 14977 39945 15011
rect 40324 14977 40358 15011
rect 40417 14977 40451 15011
rect 41061 14977 41095 15011
rect 41330 14977 41364 15011
rect 41521 14977 41555 15011
rect 43085 14977 43119 15011
rect 43361 14977 43395 15011
rect 44088 14977 44122 15011
rect 7113 14909 7147 14943
rect 7297 14909 7331 14943
rect 13829 14909 13863 14943
rect 18153 14909 18187 14943
rect 29561 14909 29595 14943
rect 30573 14909 30607 14943
rect 32689 14909 32723 14943
rect 37289 14909 37323 14943
rect 38577 14909 38611 14943
rect 38761 14909 38795 14943
rect 43821 14909 43855 14943
rect 14381 14841 14415 14875
rect 29837 14841 29871 14875
rect 34345 14841 34379 14875
rect 37565 14841 37599 14875
rect 37749 14841 37783 14875
rect 6653 14773 6687 14807
rect 7941 14773 7975 14807
rect 15577 14773 15611 14807
rect 19533 14773 19567 14807
rect 22017 14773 22051 14807
rect 30757 14773 30791 14807
rect 36645 14773 36679 14807
rect 39221 14773 39255 14807
rect 45201 14773 45235 14807
rect 45661 14773 45695 14807
rect 6377 14569 6411 14603
rect 9965 14569 9999 14603
rect 12449 14569 12483 14603
rect 13461 14569 13495 14603
rect 17049 14569 17083 14603
rect 20545 14569 20579 14603
rect 22569 14569 22603 14603
rect 23305 14569 23339 14603
rect 26893 14569 26927 14603
rect 28549 14569 28583 14603
rect 29561 14569 29595 14603
rect 32321 14569 32355 14603
rect 37289 14569 37323 14603
rect 39221 14569 39255 14603
rect 40325 14569 40359 14603
rect 41337 14569 41371 14603
rect 16405 14501 16439 14535
rect 28641 14501 28675 14535
rect 40969 14501 41003 14535
rect 15761 14433 15795 14467
rect 18245 14433 18279 14467
rect 18705 14433 18739 14467
rect 19901 14433 19935 14467
rect 29009 14433 29043 14467
rect 31953 14433 31987 14467
rect 38301 14433 38335 14467
rect 39957 14433 39991 14467
rect 42717 14433 42751 14467
rect 43453 14433 43487 14467
rect 6561 14365 6595 14399
rect 8217 14365 8251 14399
rect 10149 14365 10183 14399
rect 16221 14365 16255 14399
rect 16405 14365 16439 14399
rect 16865 14365 16899 14399
rect 17509 14365 17543 14399
rect 18337 14365 18371 14399
rect 19625 14365 19659 14399
rect 19717 14365 19751 14399
rect 20729 14365 20763 14399
rect 21189 14365 21223 14399
rect 22293 14365 22327 14399
rect 23121 14365 23155 14399
rect 29561 14365 29595 14399
rect 29837 14365 29871 14399
rect 32045 14365 32079 14399
rect 33149 14365 33183 14399
rect 35909 14365 35943 14399
rect 39129 14365 39163 14399
rect 40049 14365 40083 14399
rect 40877 14365 40911 14399
rect 41153 14365 41187 14399
rect 42533 14365 42567 14399
rect 43637 14365 43671 14399
rect 45385 14365 45419 14399
rect 45661 14365 45695 14399
rect 15516 14297 15550 14331
rect 22569 14297 22603 14331
rect 36176 14297 36210 14331
rect 38209 14297 38243 14331
rect 45017 14297 45051 14331
rect 7113 14229 7147 14263
rect 8309 14229 8343 14263
rect 14381 14229 14415 14263
rect 17601 14229 17635 14263
rect 19257 14229 19291 14263
rect 21281 14229 21315 14263
rect 22385 14229 22419 14263
rect 26433 14229 26467 14263
rect 27445 14229 27479 14263
rect 29745 14229 29779 14263
rect 33333 14229 33367 14263
rect 37749 14229 37783 14263
rect 38117 14229 38151 14263
rect 42165 14229 42199 14263
rect 42625 14229 42659 14263
rect 43729 14229 43763 14263
rect 44097 14229 44131 14263
rect 11897 14025 11931 14059
rect 15025 14025 15059 14059
rect 16773 14025 16807 14059
rect 18889 14025 18923 14059
rect 20545 14025 20579 14059
rect 23305 14025 23339 14059
rect 23673 14025 23707 14059
rect 36185 14025 36219 14059
rect 39865 14025 39899 14059
rect 41889 14025 41923 14059
rect 44281 14025 44315 14059
rect 11989 13957 12023 13991
rect 13829 13957 13863 13991
rect 18153 13957 18187 13991
rect 20177 13957 20211 13991
rect 20269 13957 20303 13991
rect 26249 13957 26283 13991
rect 35725 13957 35759 13991
rect 42686 13957 42720 13991
rect 44741 13957 44775 13991
rect 4721 13889 4755 13923
rect 10793 13889 10827 13923
rect 12817 13889 12851 13923
rect 14013 13889 14047 13923
rect 14197 13889 14231 13923
rect 14933 13889 14967 13923
rect 19349 13889 19383 13923
rect 19533 13889 19567 13923
rect 19993 13889 20027 13923
rect 20361 13889 20395 13923
rect 21005 13889 21039 13923
rect 21189 13889 21223 13923
rect 22017 13889 22051 13923
rect 23213 13889 23247 13923
rect 25513 13889 25547 13923
rect 26433 13889 26467 13923
rect 33416 13889 33450 13923
rect 36369 13889 36403 13923
rect 37473 13889 37507 13923
rect 38485 13889 38519 13923
rect 38752 13889 38786 13923
rect 41705 13889 41739 13923
rect 6745 13821 6779 13855
rect 10517 13821 10551 13855
rect 12173 13821 12207 13855
rect 13369 13821 13403 13855
rect 14749 13821 14783 13855
rect 15945 13821 15979 13855
rect 18337 13821 18371 13855
rect 21097 13821 21131 13855
rect 23121 13821 23155 13855
rect 25697 13821 25731 13855
rect 27445 13821 27479 13855
rect 27721 13821 27755 13855
rect 33149 13821 33183 13855
rect 37565 13821 37599 13855
rect 37841 13821 37875 13855
rect 40693 13821 40727 13855
rect 42441 13821 42475 13855
rect 7113 13753 7147 13787
rect 7205 13753 7239 13787
rect 10241 13753 10275 13787
rect 15393 13753 15427 13787
rect 44373 13753 44407 13787
rect 45201 13753 45235 13787
rect 4905 13685 4939 13719
rect 7665 13685 7699 13719
rect 10425 13685 10459 13719
rect 11529 13685 11563 13719
rect 19349 13685 19383 13719
rect 21833 13685 21867 13719
rect 34529 13685 34563 13719
rect 43821 13685 43855 13719
rect 6837 13481 6871 13515
rect 11897 13481 11931 13515
rect 14565 13481 14599 13515
rect 16313 13481 16347 13515
rect 16957 13481 16991 13515
rect 18245 13481 18279 13515
rect 21005 13481 21039 13515
rect 29009 13481 29043 13515
rect 30113 13481 30147 13515
rect 32965 13481 32999 13515
rect 36645 13481 36679 13515
rect 37657 13481 37691 13515
rect 38393 13481 38427 13515
rect 38945 13481 38979 13515
rect 42533 13481 42567 13515
rect 43361 13481 43395 13515
rect 43545 13481 43579 13515
rect 44005 13481 44039 13515
rect 15669 13413 15703 13447
rect 23397 13413 23431 13447
rect 25697 13413 25731 13447
rect 32505 13413 32539 13447
rect 7021 13345 7055 13379
rect 19257 13345 19291 13379
rect 21557 13345 21591 13379
rect 27537 13345 27571 13379
rect 29653 13345 29687 13379
rect 32229 13345 32263 13379
rect 33609 13345 33643 13379
rect 39865 13345 39899 13379
rect 42349 13345 42383 13379
rect 4721 13277 4755 13311
rect 4988 13277 5022 13311
rect 6561 13277 6595 13311
rect 7481 13277 7515 13311
rect 7757 13277 7791 13311
rect 10517 13277 10551 13311
rect 13093 13277 13127 13311
rect 14657 13277 14691 13311
rect 15669 13277 15703 13311
rect 15853 13277 15887 13311
rect 16497 13277 16531 13311
rect 21824 13277 21858 13311
rect 28181 13277 28215 13311
rect 29745 13277 29779 13311
rect 32137 13277 32171 13311
rect 33425 13277 33459 13311
rect 38301 13277 38335 13311
rect 39129 13277 39163 13311
rect 42257 13277 42291 13311
rect 43085 13277 43119 13311
rect 44189 13277 44223 13311
rect 7573 13209 7607 13243
rect 10784 13209 10818 13243
rect 12357 13209 12391 13243
rect 19533 13209 19567 13243
rect 27292 13209 27326 13243
rect 36553 13209 36587 13243
rect 6101 13141 6135 13175
rect 7941 13141 7975 13175
rect 22937 13141 22971 13175
rect 26157 13141 26191 13175
rect 27997 13141 28031 13175
rect 33333 13141 33367 13175
rect 41521 13141 41555 13175
rect 4997 12937 5031 12971
rect 5365 12937 5399 12971
rect 11529 12937 11563 12971
rect 14197 12937 14231 12971
rect 20085 12937 20119 12971
rect 22017 12937 22051 12971
rect 22477 12937 22511 12971
rect 26341 12937 26375 12971
rect 27261 12937 27295 12971
rect 27721 12937 27755 12971
rect 43729 12937 43763 12971
rect 6469 12869 6503 12903
rect 12449 12869 12483 12903
rect 17969 12869 18003 12903
rect 19073 12869 19107 12903
rect 20637 12869 20671 12903
rect 32689 12869 32723 12903
rect 33517 12869 33551 12903
rect 35633 12869 35667 12903
rect 39497 12869 39531 12903
rect 48789 12869 48823 12903
rect 7573 12801 7607 12835
rect 8401 12801 8435 12835
rect 8585 12801 8619 12835
rect 10425 12801 10459 12835
rect 10609 12801 10643 12835
rect 11713 12801 11747 12835
rect 13645 12801 13679 12835
rect 14105 12801 14139 12835
rect 14289 12801 14323 12835
rect 15209 12801 15243 12835
rect 15945 12801 15979 12835
rect 17233 12801 17267 12835
rect 18889 12801 18923 12835
rect 19533 12801 19567 12835
rect 19625 12801 19659 12835
rect 19809 12801 19843 12835
rect 19901 12801 19935 12835
rect 20729 12801 20763 12835
rect 22385 12801 22419 12835
rect 25513 12801 25547 12835
rect 27353 12801 27387 12835
rect 28365 12801 28399 12835
rect 37841 12801 37875 12835
rect 38761 12801 38795 12835
rect 40325 12801 40359 12835
rect 43269 12801 43303 12835
rect 48605 12801 48639 12835
rect 48881 12801 48915 12835
rect 49341 12801 49375 12835
rect 4537 12733 4571 12767
rect 5457 12733 5491 12767
rect 5549 12733 5583 12767
rect 7665 12733 7699 12767
rect 9045 12733 9079 12767
rect 9689 12733 9723 12767
rect 15301 12733 15335 12767
rect 22661 12733 22695 12767
rect 25421 12733 25455 12767
rect 27077 12733 27111 12767
rect 28273 12733 28307 12767
rect 33609 12733 33643 12767
rect 33793 12733 33827 12767
rect 6745 12665 6779 12699
rect 6929 12665 6963 12699
rect 10425 12665 10459 12699
rect 12633 12665 12667 12699
rect 25881 12665 25915 12699
rect 28733 12665 28767 12699
rect 7849 12597 7883 12631
rect 8585 12597 8619 12631
rect 14933 12597 14967 12631
rect 16037 12597 16071 12631
rect 21281 12597 21315 12631
rect 24869 12597 24903 12631
rect 33149 12597 33183 12631
rect 37749 12597 37783 12631
rect 40141 12597 40175 12631
rect 48605 12597 48639 12631
rect 49433 12597 49467 12631
rect 9597 12393 9631 12427
rect 12725 12393 12759 12427
rect 13369 12393 13403 12427
rect 16129 12393 16163 12427
rect 19993 12393 20027 12427
rect 20177 12393 20211 12427
rect 21005 12393 21039 12427
rect 21925 12393 21959 12427
rect 26985 12393 27019 12427
rect 39865 12393 39899 12427
rect 48237 12393 48271 12427
rect 48881 12393 48915 12427
rect 8217 12325 8251 12359
rect 15577 12325 15611 12359
rect 38853 12325 38887 12359
rect 48697 12325 48731 12359
rect 4905 12257 4939 12291
rect 7389 12257 7423 12291
rect 9321 12257 9355 12291
rect 35449 12257 35483 12291
rect 36093 12257 36127 12291
rect 36185 12257 36219 12291
rect 36369 12257 36403 12291
rect 9597 12189 9631 12223
rect 9689 12189 9723 12223
rect 12173 12189 12207 12223
rect 16308 12189 16342 12223
rect 16405 12189 16439 12223
rect 16625 12189 16659 12223
rect 16773 12189 16807 12223
rect 19441 12189 19475 12223
rect 20177 12189 20211 12223
rect 20269 12189 20303 12223
rect 21097 12189 21131 12223
rect 24593 12189 24627 12223
rect 25237 12189 25271 12223
rect 25605 12189 25639 12223
rect 26157 12189 26191 12223
rect 26617 12189 26651 12223
rect 26801 12189 26835 12223
rect 31493 12189 31527 12223
rect 36277 12189 36311 12223
rect 37013 12189 37047 12223
rect 37289 12189 37323 12223
rect 38577 12189 38611 12223
rect 38669 12189 38703 12223
rect 40509 12189 40543 12223
rect 40969 12189 41003 12223
rect 45201 12189 45235 12223
rect 48053 12189 48087 12223
rect 5172 12121 5206 12155
rect 7113 12121 7147 12155
rect 7941 12121 7975 12155
rect 14565 12121 14599 12155
rect 16497 12121 16531 12155
rect 20453 12121 20487 12155
rect 32137 12121 32171 12155
rect 32965 12121 32999 12155
rect 48849 12121 48883 12155
rect 49065 12121 49099 12155
rect 6285 12053 6319 12087
rect 6745 12053 6779 12087
rect 7205 12053 7239 12087
rect 8401 12053 8435 12087
rect 9505 12053 9539 12087
rect 11069 12053 11103 12087
rect 11989 12053 12023 12087
rect 14657 12053 14691 12087
rect 18705 12053 18739 12087
rect 19257 12053 19291 12087
rect 24501 12053 24535 12087
rect 31677 12053 31711 12087
rect 33609 12053 33643 12087
rect 36553 12053 36587 12087
rect 38025 12053 38059 12087
rect 41153 12053 41187 12087
rect 45109 12053 45143 12087
rect 5273 11849 5307 11883
rect 8309 11849 8343 11883
rect 10425 11849 10459 11883
rect 16681 11849 16715 11883
rect 20453 11849 20487 11883
rect 24777 11849 24811 11883
rect 25421 11849 25455 11883
rect 32781 11849 32815 11883
rect 37473 11849 37507 11883
rect 42533 11849 42567 11883
rect 45661 11849 45695 11883
rect 50813 11849 50847 11883
rect 11888 11781 11922 11815
rect 26341 11781 26375 11815
rect 30573 11781 30607 11815
rect 33486 11781 33520 11815
rect 38301 11781 38335 11815
rect 40325 11781 40359 11815
rect 46213 11781 46247 11815
rect 49985 11781 50019 11815
rect 50169 11781 50203 11815
rect 5457 11713 5491 11747
rect 7849 11713 7883 11747
rect 8033 11713 8067 11747
rect 8769 11713 8803 11747
rect 8953 11713 8987 11747
rect 10609 11713 10643 11747
rect 14197 11713 14231 11747
rect 16865 11713 16899 11747
rect 18613 11713 18647 11747
rect 18880 11713 18914 11747
rect 20729 11713 20763 11747
rect 21005 11713 21039 11747
rect 23029 11713 23063 11747
rect 25605 11713 25639 11747
rect 26249 11713 26283 11747
rect 26985 11713 27019 11747
rect 27169 11713 27203 11747
rect 28917 11713 28951 11747
rect 30481 11713 30515 11747
rect 30665 11713 30699 11747
rect 30941 11713 30975 11747
rect 31125 11713 31159 11747
rect 31401 11713 31435 11747
rect 32597 11713 32631 11747
rect 36194 11713 36228 11747
rect 36461 11713 36495 11747
rect 37289 11713 37323 11747
rect 37565 11713 37599 11747
rect 38025 11713 38059 11747
rect 40417 11713 40451 11747
rect 46121 11713 46155 11747
rect 48329 11713 48363 11747
rect 48513 11713 48547 11747
rect 48605 11713 48639 11747
rect 49249 11713 49283 11747
rect 49433 11713 49467 11747
rect 49893 11713 49927 11747
rect 50629 11713 50663 11747
rect 67373 11713 67407 11747
rect 7941 11645 7975 11679
rect 8125 11645 8159 11679
rect 10701 11645 10735 11679
rect 10793 11645 10827 11679
rect 11621 11645 11655 11679
rect 14289 11645 14323 11679
rect 15669 11645 15703 11679
rect 17049 11645 17083 11679
rect 17141 11645 17175 11679
rect 17601 11645 17635 11679
rect 23305 11645 23339 11679
rect 25237 11645 25271 11679
rect 28825 11645 28859 11679
rect 33241 11645 33275 11679
rect 39773 11645 39807 11679
rect 43913 11645 43947 11679
rect 44189 11645 44223 11679
rect 13001 11577 13035 11611
rect 15945 11577 15979 11611
rect 27077 11577 27111 11611
rect 29285 11577 29319 11611
rect 50169 11577 50203 11611
rect 7297 11509 7331 11543
rect 8953 11509 8987 11543
rect 14473 11509 14507 11543
rect 15117 11509 15151 11543
rect 16129 11509 16163 11543
rect 19993 11509 20027 11543
rect 20729 11509 20763 11543
rect 25789 11509 25823 11543
rect 27721 11509 27755 11543
rect 34621 11509 34655 11543
rect 35081 11509 35115 11543
rect 37289 11509 37323 11543
rect 42993 11509 43027 11543
rect 48145 11509 48179 11543
rect 49065 11509 49099 11543
rect 67557 11509 67591 11543
rect 8309 11305 8343 11339
rect 11253 11305 11287 11339
rect 12265 11305 12299 11339
rect 13553 11305 13587 11339
rect 19257 11305 19291 11339
rect 20821 11305 20855 11339
rect 21649 11305 21683 11339
rect 23121 11305 23155 11339
rect 26433 11305 26467 11339
rect 29561 11305 29595 11339
rect 30021 11305 30055 11339
rect 31309 11305 31343 11339
rect 33793 11305 33827 11339
rect 36737 11305 36771 11339
rect 39865 11305 39899 11339
rect 43729 11305 43763 11339
rect 46765 11305 46799 11339
rect 48145 11305 48179 11339
rect 49065 11305 49099 11339
rect 50353 11305 50387 11339
rect 67373 11305 67407 11339
rect 6193 11237 6227 11271
rect 8125 11237 8159 11271
rect 14473 11237 14507 11271
rect 16497 11237 16531 11271
rect 18705 11237 18739 11271
rect 22385 11237 22419 11271
rect 25329 11237 25363 11271
rect 28273 11237 28307 11271
rect 28457 11237 28491 11271
rect 47225 11237 47259 11271
rect 4813 11169 4847 11203
rect 7849 11169 7883 11203
rect 9045 11169 9079 11203
rect 12725 11169 12759 11203
rect 12909 11169 12943 11203
rect 14749 11169 14783 11203
rect 16681 11169 16715 11203
rect 19717 11169 19751 11203
rect 19901 11169 19935 11203
rect 23305 11169 23339 11203
rect 26893 11169 26927 11203
rect 27997 11169 28031 11203
rect 29653 11169 29687 11203
rect 30757 11169 30791 11203
rect 38209 11169 38243 11203
rect 41337 11169 41371 11203
rect 41613 11169 41647 11203
rect 45017 11169 45051 11203
rect 45293 11169 45327 11203
rect 9137 11101 9171 11135
rect 12633 11101 12667 11135
rect 14841 11101 14875 11135
rect 17509 11101 17543 11135
rect 19625 11101 19659 11135
rect 20913 11101 20947 11135
rect 21833 11101 21867 11135
rect 23397 11101 23431 11135
rect 24869 11101 24903 11135
rect 24961 11101 24995 11135
rect 25145 11101 25179 11135
rect 26065 11101 26099 11135
rect 26249 11101 26283 11135
rect 29837 11101 29871 11135
rect 30941 11101 30975 11135
rect 32882 11101 32916 11135
rect 33149 11101 33183 11135
rect 33609 11101 33643 11135
rect 37289 11101 37323 11135
rect 37473 11101 37507 11135
rect 38485 11101 38519 11135
rect 39313 11101 39347 11135
rect 42165 11101 42199 11135
rect 42349 11101 42383 11135
rect 42901 11101 42935 11135
rect 43085 11101 43119 11135
rect 43545 11101 43579 11135
rect 44281 11101 44315 11135
rect 47409 11101 47443 11135
rect 48053 11101 48087 11135
rect 48237 11101 48271 11135
rect 48697 11101 48731 11135
rect 48881 11101 48915 11135
rect 67189 11101 67223 11135
rect 67833 11101 67867 11135
rect 5080 11033 5114 11067
rect 16221 11033 16255 11067
rect 17141 11033 17175 11067
rect 17325 11033 17359 11067
rect 29561 11033 29595 11067
rect 30849 11033 30883 11067
rect 36185 11033 36219 11067
rect 37381 11033 37415 11067
rect 44373 11033 44407 11067
rect 50169 11033 50203 11067
rect 9505 10965 9539 10999
rect 20453 10965 20487 10999
rect 21373 10965 21407 10999
rect 31769 10965 31803 10999
rect 50369 10965 50403 10999
rect 50537 10965 50571 10999
rect 5181 10761 5215 10795
rect 6377 10761 6411 10795
rect 6745 10761 6779 10795
rect 8953 10761 8987 10795
rect 13277 10761 13311 10795
rect 13737 10761 13771 10795
rect 16773 10761 16807 10795
rect 20361 10761 20395 10795
rect 21925 10761 21959 10795
rect 30573 10761 30607 10795
rect 32505 10761 32539 10795
rect 33517 10761 33551 10795
rect 33885 10761 33919 10795
rect 38577 10761 38611 10795
rect 40785 10761 40819 10795
rect 43177 10761 43211 10795
rect 47041 10761 47075 10795
rect 47593 10761 47627 10795
rect 8401 10693 8435 10727
rect 33425 10693 33459 10727
rect 39129 10693 39163 10727
rect 41337 10693 41371 10727
rect 44097 10693 44131 10727
rect 47777 10693 47811 10727
rect 48789 10693 48823 10727
rect 5365 10625 5399 10659
rect 8125 10625 8159 10659
rect 8217 10625 8251 10659
rect 12164 10625 12198 10659
rect 14105 10625 14139 10659
rect 15577 10625 15611 10659
rect 20821 10625 20855 10659
rect 25881 10625 25915 10659
rect 29285 10625 29319 10659
rect 30941 10625 30975 10659
rect 32137 10625 32171 10659
rect 32321 10625 32355 10659
rect 32597 10625 32631 10659
rect 37565 10625 37599 10659
rect 37841 10625 37875 10659
rect 40233 10625 40267 10659
rect 40877 10625 40911 10659
rect 42441 10625 42475 10659
rect 46857 10625 46891 10659
rect 47041 10625 47075 10659
rect 47961 10625 47995 10659
rect 48605 10625 48639 10659
rect 48881 10625 48915 10659
rect 50169 10625 50203 10659
rect 50629 10625 50663 10659
rect 50813 10625 50847 10659
rect 6837 10557 6871 10591
rect 6929 10557 6963 10591
rect 11897 10557 11931 10591
rect 14197 10557 14231 10591
rect 15209 10557 15243 10591
rect 15485 10557 15519 10591
rect 20545 10557 20579 10591
rect 20637 10557 20671 10591
rect 20729 10557 20763 10591
rect 25973 10557 26007 10591
rect 29193 10557 29227 10591
rect 30849 10557 30883 10591
rect 33333 10557 33367 10591
rect 43821 10557 43855 10591
rect 49893 10557 49927 10591
rect 8401 10489 8435 10523
rect 26249 10489 26283 10523
rect 40049 10489 40083 10523
rect 45569 10489 45603 10523
rect 7665 10421 7699 10455
rect 25053 10421 25087 10455
rect 29653 10421 29687 10455
rect 39221 10421 39255 10455
rect 42625 10421 42659 10455
rect 48421 10421 48455 10455
rect 50813 10421 50847 10455
rect 12081 10217 12115 10251
rect 16221 10217 16255 10251
rect 20821 10217 20855 10251
rect 21189 10217 21223 10251
rect 25973 10217 26007 10251
rect 26157 10217 26191 10251
rect 28365 10217 28399 10251
rect 30389 10217 30423 10251
rect 31217 10217 31251 10251
rect 33425 10217 33459 10251
rect 40509 10217 40543 10251
rect 44465 10217 44499 10251
rect 47409 10217 47443 10251
rect 49433 10217 49467 10251
rect 50169 10217 50203 10251
rect 9229 10149 9263 10183
rect 16129 10149 16163 10183
rect 17969 10149 18003 10183
rect 24961 10149 24995 10183
rect 49525 10149 49559 10183
rect 6561 10081 6595 10115
rect 7021 10081 7055 10115
rect 8953 10081 8987 10115
rect 9321 10081 9355 10115
rect 13093 10081 13127 10115
rect 15761 10081 15795 10115
rect 16865 10081 16899 10115
rect 17141 10081 17175 10115
rect 19993 10081 20027 10115
rect 24501 10081 24535 10115
rect 29929 10081 29963 10115
rect 32137 10081 32171 10115
rect 32781 10081 32815 10115
rect 48053 10081 48087 10115
rect 49341 10081 49375 10115
rect 50446 10081 50480 10115
rect 50629 10081 50663 10115
rect 6929 10013 6963 10047
rect 9045 10013 9079 10047
rect 9229 10013 9263 10047
rect 9413 10013 9447 10047
rect 11897 10013 11931 10047
rect 12909 10013 12943 10047
rect 17233 10013 17267 10047
rect 20361 10013 20395 10047
rect 21281 10013 21315 10047
rect 22109 10013 22143 10047
rect 22385 10013 22419 10047
rect 24593 10013 24627 10047
rect 25697 10013 25731 10047
rect 30389 10013 30423 10047
rect 30665 10013 30699 10047
rect 32229 10013 32263 10047
rect 37289 10013 37323 10047
rect 38209 10013 38243 10047
rect 40049 10013 40083 10047
rect 42717 10013 42751 10047
rect 45201 10013 45235 10047
rect 45661 10013 45695 10047
rect 47225 10013 47259 10047
rect 47409 10013 47443 10047
rect 48329 10013 48363 10047
rect 49617 10013 49651 10047
rect 50327 10013 50361 10047
rect 50537 10013 50571 10047
rect 51181 10013 51215 10047
rect 20269 9945 20303 9979
rect 27997 9945 28031 9979
rect 28181 9945 28215 9979
rect 30573 9945 30607 9979
rect 39037 9945 39071 9979
rect 42993 9945 43027 9979
rect 45753 9945 45787 9979
rect 12541 9877 12575 9911
rect 13001 9877 13035 9911
rect 14197 9877 14231 9911
rect 20085 9877 20119 9911
rect 20177 9877 20211 9911
rect 23489 9877 23523 9911
rect 33977 9877 34011 9911
rect 37197 9877 37231 9911
rect 39957 9877 39991 9911
rect 45109 9877 45143 9911
rect 47593 9877 47627 9911
rect 51273 9877 51307 9911
rect 8309 9673 8343 9707
rect 16129 9673 16163 9707
rect 20361 9673 20395 9707
rect 25973 9673 26007 9707
rect 32597 9673 32631 9707
rect 38117 9673 38151 9707
rect 50169 9673 50203 9707
rect 15761 9605 15795 9639
rect 16681 9605 16715 9639
rect 17233 9605 17267 9639
rect 30849 9605 30883 9639
rect 32137 9605 32171 9639
rect 34253 9605 34287 9639
rect 47593 9605 47627 9639
rect 6653 9537 6687 9571
rect 8217 9537 8251 9571
rect 8493 9537 8527 9571
rect 9321 9537 9355 9571
rect 13185 9537 13219 9571
rect 13461 9537 13495 9571
rect 15669 9537 15703 9571
rect 15945 9537 15979 9571
rect 16865 9537 16899 9571
rect 16957 9537 16991 9571
rect 17049 9537 17083 9571
rect 20545 9537 20579 9571
rect 20729 9537 20763 9571
rect 20821 9537 20855 9571
rect 22293 9537 22327 9571
rect 24041 9537 24075 9571
rect 26157 9537 26191 9571
rect 27721 9537 27755 9571
rect 29377 9537 29411 9571
rect 30757 9537 30791 9571
rect 35265 9537 35299 9571
rect 36001 9537 36035 9571
rect 40509 9537 40543 9571
rect 40969 9537 41003 9571
rect 47869 9537 47903 9571
rect 48881 9537 48915 9571
rect 49157 9537 49191 9571
rect 49801 9537 49835 9571
rect 50077 9537 50111 9571
rect 50905 9537 50939 9571
rect 51733 9537 51767 9571
rect 6561 9469 6595 9503
rect 8953 9469 8987 9503
rect 9413 9469 9447 9503
rect 13277 9469 13311 9503
rect 21833 9469 21867 9503
rect 24501 9469 24535 9503
rect 26433 9469 26467 9503
rect 27997 9469 28031 9503
rect 30941 9469 30975 9503
rect 33425 9469 33459 9503
rect 35725 9469 35759 9503
rect 40233 9469 40267 9503
rect 43637 9469 43671 9503
rect 43913 9469 43947 9503
rect 45385 9469 45419 9503
rect 47593 9469 47627 9503
rect 49617 9469 49651 9503
rect 49985 9469 50019 9503
rect 50997 9469 51031 9503
rect 7021 9401 7055 9435
rect 8493 9401 8527 9435
rect 13645 9401 13679 9435
rect 27077 9401 27111 9435
rect 29929 9401 29963 9435
rect 32413 9401 32447 9435
rect 35081 9401 35115 9435
rect 51825 9401 51859 9435
rect 13461 9333 13495 9367
rect 22201 9333 22235 9367
rect 24133 9333 24167 9367
rect 26341 9333 26375 9367
rect 30389 9333 30423 9367
rect 36737 9333 36771 9367
rect 38761 9333 38795 9367
rect 41061 9333 41095 9367
rect 47777 9333 47811 9367
rect 49893 9333 49927 9367
rect 51273 9333 51307 9367
rect 15761 9129 15795 9163
rect 20361 9129 20395 9163
rect 21557 9129 21591 9163
rect 21925 9129 21959 9163
rect 26985 9129 27019 9163
rect 29653 9129 29687 9163
rect 30021 9129 30055 9163
rect 31861 9129 31895 9163
rect 33425 9129 33459 9163
rect 48881 9129 48915 9163
rect 49341 9129 49375 9163
rect 50169 9129 50203 9163
rect 51273 9129 51307 9163
rect 9597 9061 9631 9095
rect 15853 9061 15887 9095
rect 9781 8993 9815 9027
rect 16957 8993 16991 9027
rect 20545 8993 20579 9027
rect 25329 8993 25363 9027
rect 26157 8993 26191 9027
rect 32873 8993 32907 9027
rect 37197 8993 37231 9027
rect 39957 8993 39991 9027
rect 47777 8993 47811 9027
rect 48973 8993 49007 9027
rect 49065 8993 49099 9027
rect 9597 8925 9631 8959
rect 14565 8925 14599 8959
rect 14749 8925 14783 8959
rect 15301 8925 15335 8959
rect 17049 8925 17083 8959
rect 20361 8925 20395 8959
rect 20637 8925 20671 8959
rect 22017 8925 22051 8959
rect 28365 8925 28399 8959
rect 29009 8925 29043 8959
rect 29561 8925 29595 8959
rect 30481 8925 30515 8959
rect 33333 8925 33367 8959
rect 33517 8925 33551 8959
rect 44189 8925 44223 8959
rect 47961 8925 47995 8959
rect 48605 8925 48639 8959
rect 48789 8925 48823 8959
rect 50353 8925 50387 8959
rect 50537 8925 50571 8959
rect 50629 8925 50663 8959
rect 9965 8857 9999 8891
rect 16221 8857 16255 8891
rect 28120 8857 28154 8891
rect 30726 8857 30760 8891
rect 32505 8857 32539 8891
rect 32689 8857 32723 8891
rect 33977 8857 34011 8891
rect 36921 8857 36955 8891
rect 40233 8857 40267 8891
rect 51241 8857 51275 8891
rect 51457 8857 51491 8891
rect 14565 8789 14599 8823
rect 16681 8789 16715 8823
rect 17785 8789 17819 8823
rect 20821 8789 20855 8823
rect 22477 8789 22511 8823
rect 28825 8789 28859 8823
rect 35449 8789 35483 8823
rect 41705 8789 41739 8823
rect 44281 8789 44315 8823
rect 48145 8789 48179 8823
rect 51089 8789 51123 8823
rect 6377 8585 6411 8619
rect 6745 8585 6779 8619
rect 6837 8585 6871 8619
rect 7573 8585 7607 8619
rect 8769 8585 8803 8619
rect 11621 8585 11655 8619
rect 21833 8585 21867 8619
rect 25789 8585 25823 8619
rect 26341 8585 26375 8619
rect 27629 8585 27663 8619
rect 28089 8585 28123 8619
rect 29745 8585 29779 8619
rect 30389 8585 30423 8619
rect 31217 8585 31251 8619
rect 32137 8585 32171 8619
rect 36093 8585 36127 8619
rect 40417 8585 40451 8619
rect 40877 8585 40911 8619
rect 43545 8585 43579 8619
rect 50169 8585 50203 8619
rect 50337 8585 50371 8619
rect 9781 8517 9815 8551
rect 14565 8517 14599 8551
rect 16129 8517 16163 8551
rect 20361 8517 20395 8551
rect 24869 8517 24903 8551
rect 49249 8517 49283 8551
rect 50537 8517 50571 8551
rect 5457 8449 5491 8483
rect 9137 8449 9171 8483
rect 10793 8449 10827 8483
rect 12357 8449 12391 8483
rect 13737 8449 13771 8483
rect 14197 8449 14231 8483
rect 14351 8449 14385 8483
rect 15393 8449 15427 8483
rect 16681 8449 16715 8483
rect 16948 8449 16982 8483
rect 22109 8449 22143 8483
rect 22661 8449 22695 8483
rect 22845 8449 22879 8483
rect 23305 8449 23339 8483
rect 23489 8449 23523 8483
rect 25329 8449 25363 8483
rect 26249 8449 26283 8483
rect 26433 8449 26467 8483
rect 27721 8449 27755 8483
rect 28811 8449 28845 8483
rect 29653 8449 29687 8483
rect 32351 8449 32385 8483
rect 32505 8449 32539 8483
rect 33149 8449 33183 8483
rect 34161 8449 34195 8483
rect 34437 8449 34471 8483
rect 34621 8449 34655 8483
rect 35357 8449 35391 8483
rect 39681 8449 39715 8483
rect 40141 8449 40175 8483
rect 41061 8449 41095 8483
rect 41337 8449 41371 8483
rect 42717 8449 42751 8483
rect 45293 8449 45327 8483
rect 48513 8449 48547 8483
rect 49433 8449 49467 8483
rect 49525 8449 49559 8483
rect 7021 8381 7055 8415
rect 9229 8381 9263 8415
rect 12265 8381 12299 8415
rect 12725 8381 12759 8415
rect 15485 8381 15519 8415
rect 19533 8381 19567 8415
rect 20453 8381 20487 8415
rect 20545 8381 20579 8415
rect 21833 8381 21867 8415
rect 23397 8381 23431 8415
rect 27537 8381 27571 8415
rect 28641 8381 28675 8415
rect 30941 8381 30975 8415
rect 31125 8381 31159 8415
rect 35081 8381 35115 8415
rect 40417 8381 40451 8415
rect 42625 8381 42659 8415
rect 45017 8381 45051 8415
rect 48789 8381 48823 8415
rect 15025 8313 15059 8347
rect 18061 8313 18095 8347
rect 19993 8313 20027 8347
rect 24317 8313 24351 8347
rect 29101 8313 29135 8347
rect 31585 8313 31619 8347
rect 40233 8313 40267 8347
rect 41153 8313 41187 8347
rect 41245 8313 41279 8347
rect 43085 8313 43119 8347
rect 48697 8313 48731 8347
rect 49709 8313 49743 8347
rect 5273 8245 5307 8279
rect 22017 8245 22051 8279
rect 22845 8245 22879 8279
rect 25421 8245 25455 8279
rect 32965 8245 32999 8279
rect 34253 8245 34287 8279
rect 39589 8245 39623 8279
rect 48605 8245 48639 8279
rect 49525 8245 49559 8279
rect 50353 8245 50387 8279
rect 6469 8041 6503 8075
rect 9597 8041 9631 8075
rect 9873 8041 9907 8075
rect 10425 8041 10459 8075
rect 15117 8041 15151 8075
rect 16405 8041 16439 8075
rect 17049 8041 17083 8075
rect 19441 8041 19475 8075
rect 21281 8041 21315 8075
rect 23213 8041 23247 8075
rect 24593 8041 24627 8075
rect 25329 8041 25363 8075
rect 25789 8041 25823 8075
rect 28457 8041 28491 8075
rect 29653 8041 29687 8075
rect 30573 8041 30607 8075
rect 33793 8041 33827 8075
rect 33931 8041 33965 8075
rect 35265 8041 35299 8075
rect 35725 8041 35759 8075
rect 39313 8041 39347 8075
rect 40509 8041 40543 8075
rect 41429 8041 41463 8075
rect 41705 8041 41739 8075
rect 49341 8041 49375 8075
rect 10977 7973 11011 8007
rect 12357 7973 12391 8007
rect 21741 7973 21775 8007
rect 26433 7973 26467 8007
rect 27813 7973 27847 8007
rect 31217 7973 31251 8007
rect 5089 7905 5123 7939
rect 12081 7905 12115 7939
rect 15761 7905 15795 7939
rect 19901 7905 19935 7939
rect 27353 7905 27387 7939
rect 32597 7905 32631 7939
rect 34897 7905 34931 7939
rect 49433 7905 49467 7939
rect 5356 7837 5390 7871
rect 8033 7837 8067 7871
rect 9413 7837 9447 7871
rect 11989 7837 12023 7871
rect 12817 7837 12851 7871
rect 13001 7837 13035 7871
rect 13553 7837 13587 7871
rect 14933 7837 14967 7871
rect 16865 7837 16899 7871
rect 18429 7837 18463 7871
rect 19257 7837 19291 7871
rect 21925 7837 21959 7871
rect 22017 7837 22051 7871
rect 22293 7837 22327 7871
rect 23397 7837 23431 7871
rect 23489 7837 23523 7871
rect 24409 7837 24443 7871
rect 27445 7837 27479 7871
rect 30389 7837 30423 7871
rect 32341 7837 32375 7871
rect 33609 7837 33643 7871
rect 34069 7837 34103 7871
rect 35081 7837 35115 7871
rect 35909 7837 35943 7871
rect 39037 7837 39071 7871
rect 39313 7837 39347 7871
rect 41613 7837 41647 7871
rect 41705 7837 41739 7871
rect 42073 7837 42107 7871
rect 43913 7837 43947 7871
rect 44189 7837 44223 7871
rect 45201 7837 45235 7871
rect 48329 7837 48363 7871
rect 48513 7837 48547 7871
rect 49157 7837 49191 7871
rect 50353 7837 50387 7871
rect 11161 7769 11195 7803
rect 11345 7769 11379 7803
rect 12909 7769 12943 7803
rect 14749 7769 14783 7803
rect 18245 7769 18279 7803
rect 20168 7769 20202 7803
rect 22109 7769 22143 7803
rect 26801 7769 26835 7803
rect 28365 7769 28399 7803
rect 40325 7769 40359 7803
rect 40525 7769 40559 7803
rect 48421 7769 48455 7803
rect 7849 7701 7883 7735
rect 14289 7701 14323 7735
rect 15945 7701 15979 7735
rect 16037 7701 16071 7735
rect 26341 7701 26375 7735
rect 33057 7701 33091 7735
rect 33701 7701 33735 7735
rect 39129 7701 39163 7735
rect 40693 7701 40727 7735
rect 43729 7701 43763 7735
rect 44097 7701 44131 7735
rect 45109 7701 45143 7735
rect 48973 7701 49007 7735
rect 50169 7701 50203 7735
rect 8769 7497 8803 7531
rect 9229 7497 9263 7531
rect 9597 7497 9631 7531
rect 11529 7497 11563 7531
rect 20637 7497 20671 7531
rect 21189 7497 21223 7531
rect 28273 7497 28307 7531
rect 28825 7497 28859 7531
rect 31401 7497 31435 7531
rect 35541 7497 35575 7531
rect 41061 7497 41095 7531
rect 41797 7497 41831 7531
rect 45477 7497 45511 7531
rect 7656 7429 7690 7463
rect 10977 7429 11011 7463
rect 11989 7429 12023 7463
rect 14289 7429 14323 7463
rect 18613 7429 18647 7463
rect 22109 7429 22143 7463
rect 22293 7429 22327 7463
rect 23029 7429 23063 7463
rect 25329 7429 25363 7463
rect 27353 7429 27387 7463
rect 44005 7429 44039 7463
rect 6561 7361 6595 7395
rect 15485 7361 15519 7395
rect 19257 7361 19291 7395
rect 19513 7361 19547 7395
rect 21097 7361 21131 7395
rect 25237 7361 25271 7395
rect 26433 7361 26467 7395
rect 27721 7361 27755 7395
rect 30757 7361 30791 7395
rect 31309 7361 31343 7395
rect 32413 7361 32447 7395
rect 34437 7361 34471 7395
rect 34713 7361 34747 7395
rect 35357 7361 35391 7395
rect 37289 7361 37323 7395
rect 38025 7361 38059 7395
rect 40509 7361 40543 7395
rect 40969 7361 41003 7395
rect 41153 7361 41187 7395
rect 41613 7361 41647 7395
rect 41797 7361 41831 7395
rect 43085 7361 43119 7395
rect 43269 7361 43303 7395
rect 48513 7361 48547 7395
rect 49709 7361 49743 7395
rect 49985 7361 50019 7395
rect 7389 7293 7423 7327
rect 9689 7293 9723 7327
rect 9781 7293 9815 7327
rect 13461 7293 13495 7327
rect 14381 7293 14415 7327
rect 14565 7293 14599 7327
rect 15209 7293 15243 7327
rect 15393 7293 15427 7327
rect 16681 7293 16715 7327
rect 22753 7293 22787 7327
rect 24777 7293 24811 7327
rect 32137 7293 32171 7327
rect 35173 7293 35207 7327
rect 40233 7293 40267 7327
rect 43729 7293 43763 7327
rect 11713 7225 11747 7259
rect 12909 7225 12943 7259
rect 15853 7225 15887 7259
rect 26249 7225 26283 7259
rect 48973 7225 49007 7259
rect 6377 7157 6411 7191
rect 13921 7157 13955 7191
rect 33701 7157 33735 7191
rect 37473 7157 37507 7191
rect 38761 7157 38795 7191
rect 43269 7157 43303 7191
rect 47869 7157 47903 7191
rect 48329 7157 48363 7191
rect 7205 6953 7239 6987
rect 22109 6953 22143 6987
rect 24593 6953 24627 6987
rect 34805 6953 34839 6987
rect 40417 6953 40451 6987
rect 23581 6885 23615 6919
rect 33057 6885 33091 6919
rect 5365 6817 5399 6851
rect 7849 6817 7883 6851
rect 11529 6817 11563 6851
rect 16037 6817 16071 6851
rect 20637 6817 20671 6851
rect 26525 6817 26559 6851
rect 26709 6817 26743 6851
rect 28365 6817 28399 6851
rect 40141 6817 40175 6851
rect 45109 6817 45143 6851
rect 49617 6817 49651 6851
rect 50813 6817 50847 6851
rect 5632 6749 5666 6783
rect 7573 6749 7607 6783
rect 10701 6749 10735 6783
rect 11805 6749 11839 6783
rect 13369 6749 13403 6783
rect 16681 6749 16715 6783
rect 18521 6749 18555 6783
rect 19257 6749 19291 6783
rect 20269 6749 20303 6783
rect 20453 6749 20487 6783
rect 21557 6749 21591 6783
rect 22201 6749 22235 6783
rect 22937 6749 22971 6783
rect 23121 6749 23155 6783
rect 23857 6749 23891 6783
rect 25237 6749 25271 6783
rect 26433 6749 26467 6783
rect 29745 6749 29779 6783
rect 34897 6749 34931 6783
rect 40049 6749 40083 6783
rect 43821 6749 43855 6783
rect 44005 6749 44039 6783
rect 44235 6749 44269 6783
rect 45201 6749 45235 6783
rect 45661 6749 45695 6783
rect 47961 6749 47995 6783
rect 49341 6749 49375 6783
rect 50353 6749 50387 6783
rect 11713 6681 11747 6715
rect 14197 6681 14231 6715
rect 15792 6681 15826 6715
rect 17141 6681 17175 6715
rect 23581 6681 23615 6715
rect 24777 6681 24811 6715
rect 27813 6681 27847 6715
rect 44097 6681 44131 6715
rect 48145 6681 48179 6715
rect 6745 6613 6779 6647
rect 7665 6613 7699 6647
rect 10057 6613 10091 6647
rect 10517 6613 10551 6647
rect 12173 6613 12207 6647
rect 12817 6613 12851 6647
rect 13553 6613 13587 6647
rect 14657 6613 14691 6647
rect 16497 6613 16531 6647
rect 18705 6613 18739 6647
rect 19441 6613 19475 6647
rect 23029 6613 23063 6647
rect 23765 6613 23799 6647
rect 24409 6613 24443 6647
rect 24577 6613 24611 6647
rect 25329 6613 25363 6647
rect 26065 6613 26099 6647
rect 27261 6613 27295 6647
rect 29929 6613 29963 6647
rect 30481 6613 30515 6647
rect 43361 6613 43395 6647
rect 44373 6613 44407 6647
rect 45753 6613 45787 6647
rect 47777 6613 47811 6647
rect 48605 6613 48639 6647
rect 50169 6613 50203 6647
rect 7297 6409 7331 6443
rect 9321 6409 9355 6443
rect 9413 6409 9447 6443
rect 10977 6409 11011 6443
rect 12909 6409 12943 6443
rect 14749 6409 14783 6443
rect 18061 6409 18095 6443
rect 25605 6409 25639 6443
rect 27629 6409 27663 6443
rect 29653 6409 29687 6443
rect 31585 6409 31619 6443
rect 34805 6409 34839 6443
rect 41889 6409 41923 6443
rect 45661 6409 45695 6443
rect 7389 6341 7423 6375
rect 8217 6341 8251 6375
rect 10609 6341 10643 6375
rect 21005 6341 21039 6375
rect 22201 6341 22235 6375
rect 24133 6341 24167 6375
rect 33333 6341 33367 6375
rect 44189 6341 44223 6375
rect 11785 6273 11819 6307
rect 13369 6273 13403 6307
rect 13636 6273 13670 6307
rect 15209 6273 15243 6307
rect 15485 6273 15519 6307
rect 17693 6273 17727 6307
rect 18521 6273 18555 6307
rect 19073 6273 19107 6307
rect 23305 6273 23339 6307
rect 29193 6273 29227 6307
rect 29285 6273 29319 6307
rect 30205 6273 30239 6307
rect 30461 6273 30495 6307
rect 33057 6273 33091 6307
rect 37473 6273 37507 6307
rect 40987 6273 41021 6307
rect 41245 6273 41279 6307
rect 48329 6273 48363 6307
rect 49065 6273 49099 6307
rect 49893 6273 49927 6307
rect 50169 6273 50203 6307
rect 50629 6273 50663 6307
rect 51457 6273 51491 6307
rect 7481 6205 7515 6239
rect 9137 6205 9171 6239
rect 10425 6205 10459 6239
rect 10517 6205 10551 6239
rect 11529 6205 11563 6239
rect 17417 6205 17451 6239
rect 17601 6205 17635 6239
rect 22845 6205 22879 6239
rect 23857 6205 23891 6239
rect 27445 6205 27479 6239
rect 27537 6205 27571 6239
rect 29009 6205 29043 6239
rect 40049 6205 40083 6239
rect 40233 6205 40267 6239
rect 41086 6205 41120 6239
rect 43913 6205 43947 6239
rect 46857 6205 46891 6239
rect 48605 6205 48639 6239
rect 40693 6137 40727 6171
rect 6929 6069 6963 6103
rect 9781 6069 9815 6103
rect 16681 6069 16715 6103
rect 19257 6069 19291 6103
rect 26341 6069 26375 6103
rect 27997 6069 28031 6103
rect 37381 6069 37415 6103
rect 47593 6069 47627 6103
rect 50813 6069 50847 6103
rect 51273 6069 51307 6103
rect 7757 5865 7791 5899
rect 11897 5865 11931 5899
rect 27813 5865 27847 5899
rect 28733 5865 28767 5899
rect 32781 5865 32815 5899
rect 33885 5865 33919 5899
rect 46121 5865 46155 5899
rect 49065 5865 49099 5899
rect 7205 5797 7239 5831
rect 11437 5797 11471 5831
rect 22109 5797 22143 5831
rect 24593 5797 24627 5831
rect 25973 5797 26007 5831
rect 5825 5729 5859 5763
rect 10057 5729 10091 5763
rect 15025 5729 15059 5763
rect 19809 5729 19843 5763
rect 19993 5729 20027 5763
rect 23121 5729 23155 5763
rect 30021 5729 30055 5763
rect 30297 5729 30331 5763
rect 31033 5729 31067 5763
rect 35541 5729 35575 5763
rect 38393 5729 38427 5763
rect 40877 5729 40911 5763
rect 41153 5729 41187 5763
rect 48605 5729 48639 5763
rect 9505 5661 9539 5695
rect 10324 5661 10358 5695
rect 12081 5661 12115 5695
rect 12725 5661 12759 5695
rect 13369 5661 13403 5695
rect 14105 5661 14139 5695
rect 17417 5661 17451 5695
rect 18061 5661 18095 5695
rect 18705 5661 18739 5695
rect 19717 5661 19751 5695
rect 22937 5661 22971 5695
rect 23029 5661 23063 5695
rect 25789 5661 25823 5695
rect 26433 5661 26467 5695
rect 29929 5661 29963 5695
rect 33793 5661 33827 5695
rect 39313 5661 39347 5695
rect 40417 5661 40451 5695
rect 46581 5661 46615 5695
rect 48329 5661 48363 5695
rect 50905 5661 50939 5695
rect 51181 5661 51215 5695
rect 6092 5593 6126 5627
rect 14841 5593 14875 5627
rect 15577 5593 15611 5627
rect 16129 5593 16163 5627
rect 23765 5593 23799 5627
rect 25053 5593 25087 5627
rect 26678 5593 26712 5627
rect 31309 5593 31343 5627
rect 35817 5593 35851 5627
rect 49249 5593 49283 5627
rect 49433 5593 49467 5627
rect 9321 5525 9355 5559
rect 12909 5525 12943 5559
rect 13553 5525 13587 5559
rect 14289 5525 14323 5559
rect 16221 5525 16255 5559
rect 19349 5525 19383 5559
rect 22569 5525 22603 5559
rect 37289 5525 37323 5559
rect 37749 5525 37783 5559
rect 38117 5525 38151 5559
rect 38209 5525 38243 5559
rect 40233 5525 40267 5559
rect 47593 5525 47627 5559
rect 50169 5525 50203 5559
rect 51641 5525 51675 5559
rect 6377 5321 6411 5355
rect 10517 5321 10551 5355
rect 18613 5321 18647 5355
rect 20453 5321 20487 5355
rect 24685 5321 24719 5355
rect 28917 5321 28951 5355
rect 31125 5321 31159 5355
rect 32781 5321 32815 5355
rect 36001 5321 36035 5355
rect 37657 5321 37691 5355
rect 40785 5321 40819 5355
rect 41153 5321 41187 5355
rect 19318 5253 19352 5287
rect 24593 5253 24627 5287
rect 41245 5253 41279 5287
rect 6561 5185 6595 5219
rect 9137 5185 9171 5219
rect 9404 5185 9438 5219
rect 12449 5185 12483 5219
rect 15025 5185 15059 5219
rect 15761 5185 15795 5219
rect 18429 5185 18463 5219
rect 22477 5185 22511 5219
rect 23489 5185 23523 5219
rect 27537 5185 27571 5219
rect 27804 5185 27838 5219
rect 32873 5185 32907 5219
rect 36185 5185 36219 5219
rect 37749 5185 37783 5219
rect 38669 5185 38703 5219
rect 39865 5185 39899 5219
rect 39957 5185 39991 5219
rect 42901 5185 42935 5219
rect 43453 5185 43487 5219
rect 49801 5185 49835 5219
rect 50077 5185 50111 5219
rect 51181 5185 51215 5219
rect 51825 5185 51859 5219
rect 52745 5185 52779 5219
rect 53389 5185 53423 5219
rect 14565 5117 14599 5151
rect 19073 5117 19107 5151
rect 23213 5117 23247 5151
rect 23397 5117 23431 5151
rect 24409 5117 24443 5151
rect 37933 5117 37967 5151
rect 39773 5117 39807 5151
rect 41337 5117 41371 5151
rect 43913 5117 43947 5151
rect 45293 5117 45327 5151
rect 13921 5049 13955 5083
rect 37289 5049 37323 5083
rect 40325 5049 40359 5083
rect 42625 5049 42659 5083
rect 48237 5049 48271 5083
rect 11989 4981 12023 5015
rect 12633 4981 12667 5015
rect 13277 4981 13311 5015
rect 15117 4981 15151 5015
rect 15853 4981 15887 5015
rect 17325 4981 17359 5015
rect 17969 4981 18003 5015
rect 21925 4981 21959 5015
rect 22661 4981 22695 5015
rect 23857 4981 23891 5015
rect 25053 4981 25087 5015
rect 30665 4981 30699 5015
rect 38577 4981 38611 5015
rect 42441 4981 42475 5015
rect 45753 4981 45787 5015
rect 46397 4981 46431 5015
rect 47593 4981 47627 5015
rect 49065 4981 49099 5015
rect 50537 4981 50571 5015
rect 51365 4981 51399 5015
rect 52929 4981 52963 5015
rect 9321 4777 9355 4811
rect 14933 4777 14967 4811
rect 15853 4777 15887 4811
rect 16037 4777 16071 4811
rect 17049 4777 17083 4811
rect 20637 4777 20671 4811
rect 23857 4777 23891 4811
rect 27721 4777 27755 4811
rect 40417 4777 40451 4811
rect 41613 4777 41647 4811
rect 50813 4777 50847 4811
rect 54033 4777 54067 4811
rect 54585 4777 54619 4811
rect 55321 4777 55355 4811
rect 9873 4709 9907 4743
rect 10425 4709 10459 4743
rect 11621 4709 11655 4743
rect 14473 4709 14507 4743
rect 18061 4709 18095 4743
rect 37565 4709 37599 4743
rect 48881 4709 48915 4743
rect 52745 4709 52779 4743
rect 10977 4641 11011 4675
rect 13553 4641 13587 4675
rect 16129 4641 16163 4675
rect 19257 4641 19291 4675
rect 22477 4641 22511 4675
rect 38393 4641 38427 4675
rect 41061 4641 41095 4675
rect 42165 4641 42199 4675
rect 45661 4641 45695 4675
rect 47593 4641 47627 4675
rect 50169 4641 50203 4675
rect 53389 4641 53423 4675
rect 8401 4573 8435 4607
rect 11437 4573 11471 4607
rect 12081 4573 12115 4607
rect 12725 4573 12759 4607
rect 14289 4573 14323 4607
rect 14473 4573 14507 4607
rect 16221 4573 16255 4607
rect 16865 4573 16899 4607
rect 18705 4573 18739 4607
rect 19513 4573 19547 4607
rect 21281 4573 21315 4607
rect 21741 4573 21775 4607
rect 22744 4573 22778 4607
rect 24593 4573 24627 4607
rect 27537 4573 27571 4607
rect 30021 4573 30055 4607
rect 31125 4573 31159 4607
rect 31953 4573 31987 4607
rect 35817 4573 35851 4607
rect 38853 4573 38887 4607
rect 42993 4573 43027 4607
rect 43453 4573 43487 4607
rect 44281 4573 44315 4607
rect 45201 4573 45235 4607
rect 46305 4573 46339 4607
rect 46949 4573 46983 4607
rect 48237 4573 48271 4607
rect 49525 4573 49559 4607
rect 51457 4573 51491 4607
rect 52285 4573 52319 4607
rect 15117 4505 15151 4539
rect 15301 4505 15335 4539
rect 16681 4505 16715 4539
rect 36093 4505 36127 4539
rect 40877 4505 40911 4539
rect 41981 4505 42015 4539
rect 12265 4437 12299 4471
rect 12909 4437 12943 4471
rect 21097 4437 21131 4471
rect 24777 4437 24811 4471
rect 33609 4437 33643 4471
rect 39865 4437 39899 4471
rect 40785 4437 40819 4471
rect 42073 4437 42107 4471
rect 42809 4437 42843 4471
rect 43545 4437 43579 4471
rect 44189 4437 44223 4471
rect 45017 4437 45051 4471
rect 47133 4437 47167 4471
rect 48421 4437 48455 4471
rect 51641 4437 51675 4471
rect 52101 4437 52135 4471
rect 55965 4437 55999 4471
rect 9229 4233 9263 4267
rect 12725 4233 12759 4267
rect 15853 4233 15887 4267
rect 17785 4233 17819 4267
rect 19533 4233 19567 4267
rect 26065 4233 26099 4267
rect 33057 4233 33091 4267
rect 36553 4233 36587 4267
rect 41613 4233 41647 4267
rect 46397 4233 46431 4267
rect 49525 4233 49559 4267
rect 49709 4233 49743 4267
rect 13921 4165 13955 4199
rect 14657 4165 14691 4199
rect 15669 4165 15703 4199
rect 17325 4165 17359 4199
rect 41521 4165 41555 4199
rect 44925 4165 44959 4199
rect 8677 4097 8711 4131
rect 9781 4097 9815 4131
rect 12541 4097 12575 4131
rect 14105 4097 14139 4131
rect 15485 4097 15519 4131
rect 15761 4097 15795 4131
rect 16681 4097 16715 4131
rect 17049 4097 17083 4131
rect 17969 4097 18003 4131
rect 18153 4097 18187 4131
rect 18613 4097 18647 4131
rect 19625 4097 19659 4131
rect 20821 4097 20855 4131
rect 21005 4097 21039 4131
rect 23765 4097 23799 4131
rect 24952 4097 24986 4131
rect 29469 4097 29503 4131
rect 30297 4097 30331 4131
rect 30849 4097 30883 4131
rect 31309 4097 31343 4131
rect 32229 4097 32263 4131
rect 33149 4097 33183 4131
rect 33885 4097 33919 4131
rect 36737 4097 36771 4131
rect 37473 4097 37507 4131
rect 40417 4097 40451 4131
rect 42441 4097 42475 4131
rect 46581 4097 46615 4131
rect 47777 4097 47811 4131
rect 48421 4097 48455 4131
rect 50169 4097 50203 4131
rect 51917 4097 51951 4131
rect 54677 4097 54711 4131
rect 55229 4097 55263 4131
rect 55781 4097 55815 4131
rect 56333 4097 56367 4131
rect 67373 4097 67407 4131
rect 12081 4029 12115 4063
rect 13369 4029 13403 4063
rect 17141 4029 17175 4063
rect 19809 4029 19843 4063
rect 24685 4029 24719 4063
rect 33241 4029 33275 4063
rect 38577 4029 38611 4063
rect 41797 4029 41831 4063
rect 45201 4029 45235 4063
rect 46213 4029 46247 4063
rect 50629 4029 50663 4063
rect 54033 4029 54067 4063
rect 10977 3961 11011 3995
rect 19165 3961 19199 3995
rect 39865 3961 39899 3995
rect 41153 3961 41187 3995
rect 49157 3961 49191 3995
rect 53389 3961 53423 3995
rect 8125 3893 8159 3927
rect 10333 3893 10367 3927
rect 14749 3893 14783 3927
rect 16037 3893 16071 3927
rect 20913 3893 20947 3927
rect 21833 3893 21867 3927
rect 23121 3893 23155 3927
rect 23949 3893 23983 3927
rect 27813 3893 27847 3927
rect 29009 3893 29043 3927
rect 29561 3893 29595 3927
rect 30113 3893 30147 3927
rect 31401 3893 31435 3927
rect 32689 3893 32723 3927
rect 37381 3893 37415 3927
rect 37933 3893 37967 3927
rect 39221 3893 39255 3927
rect 40509 3893 40543 3927
rect 42625 3893 42659 3927
rect 43453 3893 43487 3927
rect 46213 3893 46247 3927
rect 47593 3893 47627 3927
rect 48237 3893 48271 3927
rect 49525 3893 49559 3927
rect 50261 3893 50295 3927
rect 51089 3893 51123 3927
rect 51733 3893 51767 3927
rect 52745 3893 52779 3927
rect 67557 3893 67591 3927
rect 11621 3689 11655 3723
rect 12265 3689 12299 3723
rect 14197 3689 14231 3723
rect 14657 3689 14691 3723
rect 15577 3689 15611 3723
rect 15715 3689 15749 3723
rect 16497 3689 16531 3723
rect 16957 3689 16991 3723
rect 20269 3689 20303 3723
rect 25789 3689 25823 3723
rect 30297 3689 30331 3723
rect 32505 3689 32539 3723
rect 35541 3689 35575 3723
rect 42809 3689 42843 3723
rect 45017 3689 45051 3723
rect 46213 3689 46247 3723
rect 47317 3689 47351 3723
rect 48605 3689 48639 3723
rect 67373 3689 67407 3723
rect 10333 3621 10367 3655
rect 12725 3621 12759 3655
rect 19717 3621 19751 3655
rect 38209 3621 38243 3655
rect 44189 3621 44223 3655
rect 50721 3621 50755 3655
rect 57897 3621 57931 3655
rect 7849 3553 7883 3587
rect 10977 3553 11011 3587
rect 14381 3553 14415 3587
rect 15485 3553 15519 3587
rect 16589 3553 16623 3587
rect 18061 3553 18095 3587
rect 20545 3553 20579 3587
rect 24409 3553 24443 3587
rect 30757 3553 30791 3587
rect 33977 3553 34011 3587
rect 36001 3553 36035 3587
rect 36277 3553 36311 3587
rect 40141 3553 40175 3587
rect 42257 3553 42291 3587
rect 45661 3553 45695 3587
rect 47133 3553 47167 3587
rect 49157 3553 49191 3587
rect 51733 3553 51767 3587
rect 55321 3553 55355 3587
rect 56609 3553 56643 3587
rect 58541 3553 58575 3587
rect 10149 3485 10183 3519
rect 11437 3485 11471 3519
rect 12081 3485 12115 3519
rect 13093 3485 13127 3519
rect 14105 3485 14139 3519
rect 16037 3485 16071 3519
rect 16773 3485 16807 3519
rect 18705 3485 18739 3519
rect 20637 3485 20671 3519
rect 21925 3485 21959 3519
rect 22385 3485 22419 3519
rect 23213 3485 23247 3519
rect 23857 3485 23891 3519
rect 24665 3485 24699 3519
rect 26249 3485 26283 3519
rect 27077 3485 27111 3519
rect 27721 3485 27755 3519
rect 28365 3485 28399 3519
rect 29009 3485 29043 3519
rect 33333 3485 33367 3519
rect 38393 3485 38427 3519
rect 38945 3485 38979 3519
rect 39865 3485 39899 3519
rect 43545 3485 43579 3519
rect 44005 3485 44039 3519
rect 47041 3485 47075 3519
rect 47869 3485 47903 3519
rect 48973 3485 49007 3519
rect 51457 3485 51491 3519
rect 52193 3485 52227 3519
rect 52837 3485 52871 3519
rect 54309 3485 54343 3519
rect 55965 3485 55999 3519
rect 57253 3485 57287 3519
rect 67189 3485 67223 3519
rect 67833 3485 67867 3519
rect 8401 3417 8435 3451
rect 9045 3417 9079 3451
rect 13001 3417 13035 3451
rect 13277 3417 13311 3451
rect 16497 3417 16531 3451
rect 20177 3417 20211 3451
rect 31033 3417 31067 3451
rect 45477 3417 45511 3451
rect 49065 3417 49099 3451
rect 53481 3417 53515 3451
rect 9689 3349 9723 3383
rect 12909 3349 12943 3383
rect 15209 3349 15243 3383
rect 20821 3349 20855 3383
rect 37749 3349 37783 3383
rect 39037 3349 39071 3383
rect 41613 3349 41647 3383
rect 42349 3349 42383 3383
rect 42441 3349 42475 3383
rect 43361 3349 43395 3383
rect 45385 3349 45419 3383
rect 50169 3349 50203 3383
rect 54125 3349 54159 3383
rect 7941 3145 7975 3179
rect 10333 3145 10367 3179
rect 12725 3145 12759 3179
rect 13369 3145 13403 3179
rect 14473 3145 14507 3179
rect 19993 3145 20027 3179
rect 21097 3145 21131 3179
rect 30849 3145 30883 3179
rect 31401 3145 31435 3179
rect 32137 3145 32171 3179
rect 32597 3145 32631 3179
rect 38301 3145 38335 3179
rect 49709 3145 49743 3179
rect 50369 3145 50403 3179
rect 50537 3145 50571 3179
rect 8493 3077 8527 3111
rect 17325 3077 17359 3111
rect 29377 3077 29411 3111
rect 39773 3077 39807 3111
rect 41613 3077 41647 3111
rect 49525 3077 49559 3111
rect 50169 3077 50203 3111
rect 7389 3009 7423 3043
rect 10149 3009 10183 3043
rect 12633 3009 12667 3043
rect 13461 3009 13495 3043
rect 14013 3009 14047 3043
rect 14289 3009 14323 3043
rect 17141 3009 17175 3043
rect 19809 3009 19843 3043
rect 21281 3009 21315 3043
rect 21833 3009 21867 3043
rect 29101 3009 29135 3043
rect 31585 3009 31619 3043
rect 32505 3009 32539 3043
rect 40049 3009 40083 3043
rect 41521 3009 41555 3043
rect 42441 3009 42475 3043
rect 45293 3009 45327 3043
rect 46029 3009 46063 3043
rect 51825 3009 51859 3043
rect 52745 3009 52779 3043
rect 53757 3009 53791 3043
rect 54493 3009 54527 3043
rect 55229 3009 55263 3043
rect 9045 2941 9079 2975
rect 12081 2941 12115 2975
rect 14105 2941 14139 2975
rect 15393 2941 15427 2975
rect 15945 2941 15979 2975
rect 19349 2941 19383 2975
rect 23213 2941 23247 2975
rect 25145 2941 25179 2975
rect 27997 2941 28031 2975
rect 32781 2941 32815 2975
rect 41797 2941 41831 2975
rect 45017 2941 45051 2975
rect 49157 2941 49191 2975
rect 55689 2941 55723 2975
rect 57897 2941 57931 2975
rect 9689 2873 9723 2907
rect 15117 2873 15151 2907
rect 18061 2873 18095 2907
rect 27353 2873 27387 2907
rect 42625 2873 42659 2907
rect 46489 2873 46523 2907
rect 47593 2873 47627 2907
rect 53573 2873 53607 2907
rect 55045 2873 55079 2907
rect 56333 2873 56367 2907
rect 58541 2873 58575 2907
rect 10977 2805 11011 2839
rect 14197 2805 14231 2839
rect 15485 2805 15519 2839
rect 15577 2805 15611 2839
rect 18705 2805 18739 2839
rect 20637 2805 20671 2839
rect 22569 2805 22603 2839
rect 23857 2805 23891 2839
rect 24501 2805 24535 2839
rect 25789 2805 25823 2839
rect 26433 2805 26467 2839
rect 28641 2805 28675 2839
rect 33793 2805 33827 2839
rect 34253 2805 34287 2839
rect 34897 2805 34931 2839
rect 35541 2805 35575 2839
rect 36369 2805 36403 2839
rect 37289 2805 37323 2839
rect 40509 2805 40543 2839
rect 41153 2805 41187 2839
rect 43545 2805 43579 2839
rect 45845 2805 45879 2839
rect 48237 2805 48271 2839
rect 49525 2805 49559 2839
rect 50353 2805 50387 2839
rect 51089 2805 51123 2839
rect 51641 2805 51675 2839
rect 52929 2805 52963 2839
rect 54309 2805 54343 2839
rect 56977 2805 57011 2839
rect 14473 2601 14507 2635
rect 16037 2601 16071 2635
rect 16773 2601 16807 2635
rect 19349 2601 19383 2635
rect 19993 2601 20027 2635
rect 32229 2601 32263 2635
rect 56149 2601 56183 2635
rect 56793 2601 56827 2635
rect 8401 2533 8435 2567
rect 15117 2533 15151 2567
rect 17509 2533 17543 2567
rect 18705 2533 18739 2567
rect 22569 2533 22603 2567
rect 25789 2533 25823 2567
rect 27721 2533 27755 2567
rect 30297 2533 30331 2567
rect 32873 2533 32907 2567
rect 41521 2533 41555 2567
rect 44097 2533 44131 2567
rect 45201 2533 45235 2567
rect 45845 2533 45879 2567
rect 46489 2533 46523 2567
rect 49341 2533 49375 2567
rect 53665 2533 53699 2567
rect 58541 2533 58575 2567
rect 7757 2465 7791 2499
rect 12725 2465 12759 2499
rect 20637 2465 20671 2499
rect 23213 2465 23247 2499
rect 25145 2465 25179 2499
rect 26433 2465 26467 2499
rect 28365 2465 28399 2499
rect 30941 2465 30975 2499
rect 37933 2465 37967 2499
rect 39313 2465 39347 2499
rect 47961 2465 47995 2499
rect 59185 2465 59219 2499
rect 6653 2397 6687 2431
rect 8217 2397 8251 2431
rect 9689 2397 9723 2431
rect 10333 2397 10367 2431
rect 10977 2397 11011 2431
rect 12541 2397 12575 2431
rect 14657 2397 14691 2431
rect 17693 2397 17727 2431
rect 19809 2397 19843 2431
rect 21281 2397 21315 2431
rect 23857 2397 23891 2431
rect 29009 2397 29043 2431
rect 31585 2397 31619 2431
rect 33517 2397 33551 2431
rect 34161 2397 34195 2431
rect 34989 2397 35023 2431
rect 35633 2397 35667 2431
rect 36093 2397 36127 2431
rect 37289 2397 37323 2431
rect 38577 2397 38611 2431
rect 40233 2397 40267 2431
rect 40969 2397 41003 2431
rect 41705 2397 41739 2431
rect 42441 2397 42475 2431
rect 43177 2397 43211 2431
rect 43913 2397 43947 2431
rect 45017 2397 45051 2431
rect 46029 2397 46063 2431
rect 48697 2397 48731 2431
rect 49525 2397 49559 2431
rect 50353 2397 50387 2431
rect 51273 2397 51307 2431
rect 51733 2397 51767 2431
rect 53021 2397 53055 2431
rect 53481 2397 53515 2431
rect 54493 2397 54527 2431
rect 55597 2397 55631 2431
rect 57897 2397 57931 2431
rect 7205 2329 7239 2363
rect 11897 2329 11931 2363
rect 12081 2329 12115 2363
rect 15301 2329 15335 2363
rect 15945 2329 15979 2363
rect 16865 2329 16899 2363
rect 24409 2329 24443 2363
rect 46673 2329 46707 2363
rect 48145 2329 48179 2363
rect 56241 2329 56275 2363
rect 9045 2261 9079 2295
rect 13553 2261 13587 2295
rect 21833 2261 21867 2295
rect 40049 2261 40083 2295
rect 40785 2261 40819 2295
rect 42625 2261 42659 2295
rect 43361 2261 43395 2295
rect 50169 2261 50203 2295
rect 51089 2261 51123 2295
rect 51917 2261 51951 2295
rect 52837 2261 52871 2295
rect 54309 2261 54343 2295
rect 55413 2261 55447 2295
<< metal1 >>
rect 1104 57690 68816 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 68816 57690
rect 1104 57616 68816 57638
rect 4338 57440 4344 57452
rect 4299 57412 4344 57440
rect 4338 57400 4344 57412
rect 4396 57400 4402 57452
rect 4890 57400 4896 57452
rect 4948 57440 4954 57452
rect 4985 57443 5043 57449
rect 4985 57440 4997 57443
rect 4948 57412 4997 57440
rect 4948 57400 4954 57412
rect 4985 57409 4997 57412
rect 5031 57409 5043 57443
rect 4985 57403 5043 57409
rect 5813 57443 5871 57449
rect 5813 57409 5825 57443
rect 5859 57440 5871 57443
rect 5994 57440 6000 57452
rect 5859 57412 6000 57440
rect 5859 57409 5871 57412
rect 5813 57403 5871 57409
rect 5994 57400 6000 57412
rect 6052 57400 6058 57452
rect 6546 57400 6552 57452
rect 6604 57440 6610 57452
rect 6641 57443 6699 57449
rect 6641 57440 6653 57443
rect 6604 57412 6653 57440
rect 6604 57400 6610 57412
rect 6641 57409 6653 57412
rect 6687 57409 6699 57443
rect 6641 57403 6699 57409
rect 7561 57443 7619 57449
rect 7561 57409 7573 57443
rect 7607 57440 7619 57443
rect 7650 57440 7656 57452
rect 7607 57412 7656 57440
rect 7607 57409 7619 57412
rect 7561 57403 7619 57409
rect 7650 57400 7656 57412
rect 7708 57400 7714 57452
rect 8202 57440 8208 57452
rect 8163 57412 8208 57440
rect 8202 57400 8208 57412
rect 8260 57400 8266 57452
rect 9306 57440 9312 57452
rect 9267 57412 9312 57440
rect 9306 57400 9312 57412
rect 9364 57400 9370 57452
rect 9858 57400 9864 57452
rect 9916 57440 9922 57452
rect 9953 57443 10011 57449
rect 9953 57440 9965 57443
rect 9916 57412 9965 57440
rect 9916 57400 9922 57412
rect 9953 57409 9965 57412
rect 9999 57409 10011 57443
rect 10962 57440 10968 57452
rect 10923 57412 10968 57440
rect 9953 57403 10011 57409
rect 10962 57400 10968 57412
rect 11020 57400 11026 57452
rect 11514 57400 11520 57452
rect 11572 57440 11578 57452
rect 11609 57443 11667 57449
rect 11609 57440 11621 57443
rect 11572 57412 11621 57440
rect 11572 57400 11578 57412
rect 11609 57409 11621 57412
rect 11655 57409 11667 57443
rect 12618 57440 12624 57452
rect 12579 57412 12624 57440
rect 11609 57403 11667 57409
rect 12618 57400 12624 57412
rect 12676 57400 12682 57452
rect 13170 57400 13176 57452
rect 13228 57440 13234 57452
rect 13265 57443 13323 57449
rect 13265 57440 13277 57443
rect 13228 57412 13277 57440
rect 13228 57400 13234 57412
rect 13265 57409 13277 57412
rect 13311 57409 13323 57443
rect 14274 57440 14280 57452
rect 14235 57412 14280 57440
rect 13265 57403 13323 57409
rect 14274 57400 14280 57412
rect 14332 57400 14338 57452
rect 14826 57400 14832 57452
rect 14884 57440 14890 57452
rect 14921 57443 14979 57449
rect 14921 57440 14933 57443
rect 14884 57412 14933 57440
rect 14884 57400 14890 57412
rect 14921 57409 14933 57412
rect 14967 57409 14979 57443
rect 15930 57440 15936 57452
rect 15891 57412 15936 57440
rect 14921 57403 14979 57409
rect 15930 57400 15936 57412
rect 15988 57400 15994 57452
rect 17586 57440 17592 57452
rect 17547 57412 17592 57440
rect 17586 57400 17592 57412
rect 17644 57400 17650 57452
rect 18138 57400 18144 57452
rect 18196 57440 18202 57452
rect 18233 57443 18291 57449
rect 18233 57440 18245 57443
rect 18196 57412 18245 57440
rect 18196 57400 18202 57412
rect 18233 57409 18245 57412
rect 18279 57409 18291 57443
rect 19242 57440 19248 57452
rect 19203 57412 19248 57440
rect 18233 57403 18291 57409
rect 19242 57400 19248 57412
rect 19300 57400 19306 57452
rect 19889 57443 19947 57449
rect 19889 57409 19901 57443
rect 19935 57440 19947 57443
rect 19978 57440 19984 57452
rect 19935 57412 19984 57440
rect 19935 57409 19947 57412
rect 19889 57403 19947 57409
rect 19978 57400 19984 57412
rect 20036 57400 20042 57452
rect 20898 57400 20904 57452
rect 20956 57440 20962 57452
rect 20993 57443 21051 57449
rect 20993 57440 21005 57443
rect 20956 57412 21005 57440
rect 20956 57400 20962 57412
rect 20993 57409 21005 57412
rect 21039 57409 21051 57443
rect 20993 57403 21051 57409
rect 21450 57400 21456 57452
rect 21508 57440 21514 57452
rect 21821 57443 21879 57449
rect 21821 57440 21833 57443
rect 21508 57412 21833 57440
rect 21508 57400 21514 57412
rect 21821 57409 21833 57412
rect 21867 57409 21879 57443
rect 22554 57440 22560 57452
rect 22515 57412 22560 57440
rect 21821 57403 21879 57409
rect 22554 57400 22560 57412
rect 22612 57400 22618 57452
rect 23106 57400 23112 57452
rect 23164 57440 23170 57452
rect 23201 57443 23259 57449
rect 23201 57440 23213 57443
rect 23164 57412 23213 57440
rect 23164 57400 23170 57412
rect 23201 57409 23213 57412
rect 23247 57409 23259 57443
rect 24854 57440 24860 57452
rect 24815 57412 24860 57440
rect 23201 57403 23259 57409
rect 24854 57400 24860 57412
rect 24912 57400 24918 57452
rect 25777 57443 25835 57449
rect 25777 57409 25789 57443
rect 25823 57440 25835 57443
rect 25866 57440 25872 57452
rect 25823 57412 25872 57440
rect 25823 57409 25835 57412
rect 25777 57403 25835 57409
rect 25866 57400 25872 57412
rect 25924 57400 25930 57452
rect 26418 57440 26424 57452
rect 26379 57412 26424 57440
rect 26418 57400 26424 57412
rect 26476 57400 26482 57452
rect 27522 57440 27528 57452
rect 27483 57412 27528 57440
rect 27522 57400 27528 57412
rect 27580 57400 27586 57452
rect 28074 57400 28080 57452
rect 28132 57440 28138 57452
rect 28169 57443 28227 57449
rect 28169 57440 28181 57443
rect 28132 57412 28181 57440
rect 28132 57400 28138 57412
rect 28169 57409 28181 57412
rect 28215 57409 28227 57443
rect 28169 57403 28227 57409
rect 28997 57443 29055 57449
rect 28997 57409 29009 57443
rect 29043 57440 29055 57443
rect 29178 57440 29184 57452
rect 29043 57412 29184 57440
rect 29043 57409 29055 57412
rect 28997 57403 29055 57409
rect 29178 57400 29184 57412
rect 29236 57400 29242 57452
rect 29730 57400 29736 57452
rect 29788 57440 29794 57452
rect 29825 57443 29883 57449
rect 29825 57440 29837 57443
rect 29788 57412 29837 57440
rect 29788 57400 29794 57412
rect 29825 57409 29837 57412
rect 29871 57409 29883 57443
rect 29825 57403 29883 57409
rect 30745 57443 30803 57449
rect 30745 57409 30757 57443
rect 30791 57440 30803 57443
rect 30834 57440 30840 57452
rect 30791 57412 30840 57440
rect 30791 57409 30803 57412
rect 30745 57403 30803 57409
rect 30834 57400 30840 57412
rect 30892 57400 30898 57452
rect 31386 57440 31392 57452
rect 31347 57412 31392 57440
rect 31386 57400 31392 57412
rect 31444 57400 31450 57452
rect 32490 57440 32496 57452
rect 32451 57412 32496 57440
rect 32490 57400 32496 57412
rect 32548 57400 32554 57452
rect 33134 57440 33140 57452
rect 33095 57412 33140 57440
rect 33134 57400 33140 57412
rect 33192 57400 33198 57452
rect 34146 57440 34152 57452
rect 34107 57412 34152 57440
rect 34146 57400 34152 57412
rect 34204 57400 34210 57452
rect 34698 57400 34704 57452
rect 34756 57440 34762 57452
rect 34793 57443 34851 57449
rect 34793 57440 34805 57443
rect 34756 57412 34805 57440
rect 34756 57400 34762 57412
rect 34793 57409 34805 57412
rect 34839 57409 34851 57443
rect 34793 57403 34851 57409
rect 36354 57400 36360 57452
rect 36412 57440 36418 57452
rect 36541 57443 36599 57449
rect 36541 57440 36553 57443
rect 36412 57412 36553 57440
rect 36412 57400 36418 57412
rect 36541 57409 36553 57412
rect 36587 57409 36599 57443
rect 36541 57403 36599 57409
rect 37458 57400 37464 57452
rect 37516 57440 37522 57452
rect 37553 57443 37611 57449
rect 37553 57440 37565 57443
rect 37516 57412 37565 57440
rect 37516 57400 37522 57412
rect 37553 57409 37565 57412
rect 37599 57409 37611 57443
rect 37553 57403 37611 57409
rect 38010 57400 38016 57452
rect 38068 57440 38074 57452
rect 38197 57443 38255 57449
rect 38197 57440 38209 57443
rect 38068 57412 38209 57440
rect 38068 57400 38074 57412
rect 38197 57409 38209 57412
rect 38243 57409 38255 57443
rect 38197 57403 38255 57409
rect 39114 57400 39120 57452
rect 39172 57440 39178 57452
rect 39853 57443 39911 57449
rect 39853 57440 39865 57443
rect 39172 57412 39865 57440
rect 39172 57400 39178 57412
rect 39853 57409 39865 57412
rect 39899 57409 39911 57443
rect 39853 57403 39911 57409
rect 40034 57400 40040 57452
rect 40092 57440 40098 57452
rect 40497 57443 40555 57449
rect 40497 57440 40509 57443
rect 40092 57412 40509 57440
rect 40092 57400 40098 57412
rect 40497 57409 40509 57412
rect 40543 57409 40555 57443
rect 40497 57403 40555 57409
rect 40770 57400 40776 57452
rect 40828 57440 40834 57452
rect 41141 57443 41199 57449
rect 41141 57440 41153 57443
rect 40828 57412 41153 57440
rect 40828 57400 40834 57412
rect 41141 57409 41153 57412
rect 41187 57409 41199 57443
rect 41141 57403 41199 57409
rect 42426 57400 42432 57452
rect 42484 57440 42490 57452
rect 42521 57443 42579 57449
rect 42521 57440 42533 57443
rect 42484 57412 42533 57440
rect 42484 57400 42490 57412
rect 42521 57409 42533 57412
rect 42567 57409 42579 57443
rect 42521 57403 42579 57409
rect 42978 57400 42984 57452
rect 43036 57440 43042 57452
rect 43165 57443 43223 57449
rect 43165 57440 43177 57443
rect 43036 57412 43177 57440
rect 43036 57400 43042 57412
rect 43165 57409 43177 57412
rect 43211 57409 43223 57443
rect 44174 57440 44180 57452
rect 44135 57412 44180 57440
rect 43165 57403 43223 57409
rect 44174 57400 44180 57412
rect 44232 57400 44238 57452
rect 44634 57400 44640 57452
rect 44692 57440 44698 57452
rect 45005 57443 45063 57449
rect 45005 57440 45017 57443
rect 44692 57412 45017 57440
rect 44692 57400 44698 57412
rect 45005 57409 45017 57412
rect 45051 57409 45063 57443
rect 45005 57403 45063 57409
rect 45738 57400 45744 57452
rect 45796 57440 45802 57452
rect 45833 57443 45891 57449
rect 45833 57440 45845 57443
rect 45796 57412 45845 57440
rect 45796 57400 45802 57412
rect 45833 57409 45845 57412
rect 45879 57409 45891 57443
rect 45833 57403 45891 57409
rect 46290 57400 46296 57452
rect 46348 57440 46354 57452
rect 46477 57443 46535 57449
rect 46477 57440 46489 57443
rect 46348 57412 46489 57440
rect 46348 57400 46354 57412
rect 46477 57409 46489 57412
rect 46523 57409 46535 57443
rect 46477 57403 46535 57409
rect 47394 57400 47400 57452
rect 47452 57440 47458 57452
rect 47581 57443 47639 57449
rect 47581 57440 47593 57443
rect 47452 57412 47593 57440
rect 47452 57400 47458 57412
rect 47581 57409 47593 57412
rect 47627 57409 47639 57443
rect 47581 57403 47639 57409
rect 47946 57400 47952 57452
rect 48004 57440 48010 57452
rect 48225 57443 48283 57449
rect 48225 57440 48237 57443
rect 48004 57412 48237 57440
rect 48004 57400 48010 57412
rect 48225 57409 48237 57412
rect 48271 57409 48283 57443
rect 48225 57403 48283 57409
rect 49050 57400 49056 57452
rect 49108 57440 49114 57452
rect 49145 57443 49203 57449
rect 49145 57440 49157 57443
rect 49108 57412 49157 57440
rect 49108 57400 49114 57412
rect 49145 57409 49157 57412
rect 49191 57409 49203 57443
rect 49145 57403 49203 57409
rect 49694 57400 49700 57452
rect 49752 57440 49758 57452
rect 50157 57443 50215 57449
rect 50157 57440 50169 57443
rect 49752 57412 50169 57440
rect 49752 57400 49758 57412
rect 50157 57409 50169 57412
rect 50203 57409 50215 57443
rect 50157 57403 50215 57409
rect 50706 57400 50712 57452
rect 50764 57440 50770 57452
rect 50801 57443 50859 57449
rect 50801 57440 50813 57443
rect 50764 57412 50813 57440
rect 50764 57400 50770 57412
rect 50801 57409 50813 57412
rect 50847 57409 50859 57443
rect 50801 57403 50859 57409
rect 51258 57400 51264 57452
rect 51316 57440 51322 57452
rect 51445 57443 51503 57449
rect 51445 57440 51457 57443
rect 51316 57412 51457 57440
rect 51316 57400 51322 57412
rect 51445 57409 51457 57412
rect 51491 57409 51503 57443
rect 51445 57403 51503 57409
rect 52454 57400 52460 57452
rect 52512 57440 52518 57452
rect 52733 57443 52791 57449
rect 52733 57440 52745 57443
rect 52512 57412 52745 57440
rect 52512 57400 52518 57412
rect 52733 57409 52745 57412
rect 52779 57409 52791 57443
rect 52733 57403 52791 57409
rect 52914 57400 52920 57452
rect 52972 57440 52978 57452
rect 53377 57443 53435 57449
rect 53377 57440 53389 57443
rect 52972 57412 53389 57440
rect 52972 57400 52978 57412
rect 53377 57409 53389 57412
rect 53423 57409 53435 57443
rect 53377 57403 53435 57409
rect 54018 57400 54024 57452
rect 54076 57440 54082 57452
rect 54113 57443 54171 57449
rect 54113 57440 54125 57443
rect 54076 57412 54125 57440
rect 54076 57400 54082 57412
rect 54113 57409 54125 57412
rect 54159 57409 54171 57443
rect 54113 57403 54171 57409
rect 55674 57400 55680 57452
rect 55732 57440 55738 57452
rect 55953 57443 56011 57449
rect 55953 57440 55965 57443
rect 55732 57412 55965 57440
rect 55732 57400 55738 57412
rect 55953 57409 55965 57412
rect 55999 57409 56011 57443
rect 56594 57440 56600 57452
rect 56555 57412 56600 57440
rect 55953 57403 56011 57409
rect 56594 57400 56600 57412
rect 56652 57400 56658 57452
rect 57330 57400 57336 57452
rect 57388 57440 57394 57452
rect 57885 57443 57943 57449
rect 57885 57440 57897 57443
rect 57388 57412 57897 57440
rect 57388 57400 57394 57412
rect 57885 57409 57897 57412
rect 57931 57409 57943 57443
rect 57885 57403 57943 57409
rect 57974 57400 57980 57452
rect 58032 57440 58038 57452
rect 58529 57443 58587 57449
rect 58529 57440 58541 57443
rect 58032 57412 58541 57440
rect 58032 57400 58038 57412
rect 58529 57409 58541 57412
rect 58575 57409 58587 57443
rect 58529 57403 58587 57409
rect 58986 57400 58992 57452
rect 59044 57440 59050 57452
rect 59173 57443 59231 57449
rect 59173 57440 59185 57443
rect 59044 57412 59185 57440
rect 59044 57400 59050 57412
rect 59173 57409 59185 57412
rect 59219 57409 59231 57443
rect 59173 57403 59231 57409
rect 59538 57400 59544 57452
rect 59596 57440 59602 57452
rect 60461 57443 60519 57449
rect 60461 57440 60473 57443
rect 59596 57412 60473 57440
rect 59596 57400 59602 57412
rect 60461 57409 60473 57412
rect 60507 57409 60519 57443
rect 60461 57403 60519 57409
rect 60734 57400 60740 57452
rect 60792 57440 60798 57452
rect 61105 57443 61163 57449
rect 61105 57440 61117 57443
rect 60792 57412 61117 57440
rect 60792 57400 60798 57412
rect 61105 57409 61117 57412
rect 61151 57409 61163 57443
rect 61105 57403 61163 57409
rect 61194 57400 61200 57452
rect 61252 57440 61258 57452
rect 61749 57443 61807 57449
rect 61749 57440 61761 57443
rect 61252 57412 61761 57440
rect 61252 57400 61258 57412
rect 61749 57409 61761 57412
rect 61795 57409 61807 57443
rect 61749 57403 61807 57409
rect 62298 57400 62304 57452
rect 62356 57440 62362 57452
rect 63037 57443 63095 57449
rect 63037 57440 63049 57443
rect 62356 57412 63049 57440
rect 62356 57400 62362 57412
rect 63037 57409 63049 57412
rect 63083 57409 63095 57443
rect 63037 57403 63095 57409
rect 63954 57400 63960 57452
rect 64012 57440 64018 57452
rect 64325 57443 64383 57449
rect 64325 57440 64337 57443
rect 64012 57412 64337 57440
rect 64012 57400 64018 57412
rect 64325 57409 64337 57412
rect 64371 57409 64383 57443
rect 64325 57403 64383 57409
rect 65610 57400 65616 57452
rect 65668 57440 65674 57452
rect 65705 57443 65763 57449
rect 65705 57440 65717 57443
rect 65668 57412 65717 57440
rect 65668 57400 65674 57412
rect 65705 57409 65717 57412
rect 65751 57409 65763 57443
rect 65705 57403 65763 57409
rect 66254 57400 66260 57452
rect 66312 57440 66318 57452
rect 66349 57443 66407 57449
rect 66349 57440 66361 57443
rect 66312 57412 66361 57440
rect 66312 57400 66318 57412
rect 66349 57409 66361 57412
rect 66395 57409 66407 57443
rect 66349 57403 66407 57409
rect 16482 57332 16488 57384
rect 16540 57372 16546 57384
rect 16669 57375 16727 57381
rect 16669 57372 16681 57375
rect 16540 57344 16681 57372
rect 16540 57332 16546 57344
rect 16669 57341 16681 57344
rect 16715 57341 16727 57375
rect 16669 57335 16727 57341
rect 35802 57332 35808 57384
rect 35860 57372 35866 57384
rect 35897 57375 35955 57381
rect 35897 57372 35909 57375
rect 35860 57344 35909 57372
rect 35860 57332 35866 57344
rect 35897 57341 35909 57344
rect 35943 57341 35955 57375
rect 35897 57335 35955 57341
rect 62850 57332 62856 57384
rect 62908 57372 62914 57384
rect 63681 57375 63739 57381
rect 63681 57372 63693 57375
rect 62908 57344 63693 57372
rect 62908 57332 62914 57344
rect 63681 57341 63693 57344
rect 63727 57341 63739 57375
rect 63681 57335 63739 57341
rect 54570 57264 54576 57316
rect 54628 57304 54634 57316
rect 55309 57307 55367 57313
rect 55309 57304 55321 57307
rect 54628 57276 55321 57304
rect 54628 57264 54634 57276
rect 55309 57273 55321 57276
rect 55355 57273 55367 57307
rect 55309 57267 55367 57273
rect 1104 57146 68816 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 65654 57146
rect 65706 57094 65718 57146
rect 65770 57094 65782 57146
rect 65834 57094 65846 57146
rect 65898 57094 65910 57146
rect 65962 57094 68816 57146
rect 1104 57072 68816 57094
rect 24210 56992 24216 57044
rect 24268 57032 24274 57044
rect 24397 57035 24455 57041
rect 24397 57032 24409 57035
rect 24268 57004 24409 57032
rect 24268 56992 24274 57004
rect 24397 57001 24409 57004
rect 24443 57001 24455 57035
rect 41414 57032 41420 57044
rect 41375 57004 41420 57032
rect 24397 56995 24455 57001
rect 41414 56992 41420 57004
rect 41472 56992 41478 57044
rect 64506 56992 64512 57044
rect 64564 57032 64570 57044
rect 64601 57035 64659 57041
rect 64601 57032 64613 57035
rect 64564 57004 64613 57032
rect 64564 56992 64570 57004
rect 64601 57001 64613 57004
rect 64647 57001 64659 57035
rect 64601 56995 64659 57001
rect 1104 56602 68816 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 68816 56602
rect 1104 56528 68816 56550
rect 67358 56352 67364 56364
rect 67319 56324 67364 56352
rect 67358 56312 67364 56324
rect 67416 56312 67422 56364
rect 67542 56148 67548 56160
rect 67503 56120 67548 56148
rect 67542 56108 67548 56120
rect 67600 56108 67606 56160
rect 1104 56058 68816 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 65654 56058
rect 65706 56006 65718 56058
rect 65770 56006 65782 56058
rect 65834 56006 65846 56058
rect 65898 56006 65910 56058
rect 65962 56006 68816 56058
rect 1104 55984 68816 56006
rect 1104 55514 68816 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 68816 55514
rect 1104 55440 68816 55462
rect 1104 54970 68816 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 65654 54970
rect 65706 54918 65718 54970
rect 65770 54918 65782 54970
rect 65834 54918 65846 54970
rect 65898 54918 65910 54970
rect 65962 54918 68816 54970
rect 1104 54896 68816 54918
rect 1104 54426 68816 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 68816 54426
rect 1104 54352 68816 54374
rect 1104 53882 68816 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 65654 53882
rect 65706 53830 65718 53882
rect 65770 53830 65782 53882
rect 65834 53830 65846 53882
rect 65898 53830 65910 53882
rect 65962 53830 68816 53882
rect 1104 53808 68816 53830
rect 1104 53338 68816 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 68816 53338
rect 1104 53264 68816 53286
rect 1104 52794 68816 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 65654 52794
rect 65706 52742 65718 52794
rect 65770 52742 65782 52794
rect 65834 52742 65846 52794
rect 65898 52742 65910 52794
rect 65962 52742 68816 52794
rect 1104 52720 68816 52742
rect 1104 52250 68816 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 68816 52250
rect 1104 52176 68816 52198
rect 1104 51706 68816 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 65654 51706
rect 65706 51654 65718 51706
rect 65770 51654 65782 51706
rect 65834 51654 65846 51706
rect 65898 51654 65910 51706
rect 65962 51654 68816 51706
rect 1104 51632 68816 51654
rect 1104 51162 68816 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 68816 51162
rect 1104 51088 68816 51110
rect 1104 50618 68816 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 65654 50618
rect 65706 50566 65718 50618
rect 65770 50566 65782 50618
rect 65834 50566 65846 50618
rect 65898 50566 65910 50618
rect 65962 50566 68816 50618
rect 1104 50544 68816 50566
rect 1104 50074 68816 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 68816 50074
rect 1104 50000 68816 50022
rect 1104 49530 68816 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 65654 49530
rect 65706 49478 65718 49530
rect 65770 49478 65782 49530
rect 65834 49478 65846 49530
rect 65898 49478 65910 49530
rect 65962 49478 68816 49530
rect 1104 49456 68816 49478
rect 1104 48986 68816 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 68816 48986
rect 1104 48912 68816 48934
rect 67361 48739 67419 48745
rect 67361 48705 67373 48739
rect 67407 48736 67419 48739
rect 67450 48736 67456 48748
rect 67407 48708 67456 48736
rect 67407 48705 67419 48708
rect 67361 48699 67419 48705
rect 67450 48696 67456 48708
rect 67508 48696 67514 48748
rect 67542 48600 67548 48612
rect 67503 48572 67548 48600
rect 67542 48560 67548 48572
rect 67600 48560 67606 48612
rect 1104 48442 68816 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 65654 48442
rect 65706 48390 65718 48442
rect 65770 48390 65782 48442
rect 65834 48390 65846 48442
rect 65898 48390 65910 48442
rect 65962 48390 68816 48442
rect 1104 48368 68816 48390
rect 1104 47898 68816 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 68816 47898
rect 1104 47824 68816 47846
rect 1104 47354 68816 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 65654 47354
rect 65706 47302 65718 47354
rect 65770 47302 65782 47354
rect 65834 47302 65846 47354
rect 65898 47302 65910 47354
rect 65962 47302 68816 47354
rect 1104 47280 68816 47302
rect 1104 46810 68816 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 68816 46810
rect 1104 46736 68816 46758
rect 1104 46266 68816 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 65654 46266
rect 65706 46214 65718 46266
rect 65770 46214 65782 46266
rect 65834 46214 65846 46266
rect 65898 46214 65910 46266
rect 65962 46214 68816 46266
rect 1104 46192 68816 46214
rect 1104 45722 68816 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 68816 45722
rect 1104 45648 68816 45670
rect 43990 45432 43996 45484
rect 44048 45472 44054 45484
rect 66625 45475 66683 45481
rect 66625 45472 66637 45475
rect 44048 45444 66637 45472
rect 44048 45432 44054 45444
rect 66625 45441 66637 45444
rect 66671 45472 66683 45475
rect 67177 45475 67235 45481
rect 67177 45472 67189 45475
rect 66671 45444 67189 45472
rect 66671 45441 66683 45444
rect 66625 45435 66683 45441
rect 67177 45441 67189 45444
rect 67223 45441 67235 45475
rect 67177 45435 67235 45441
rect 67358 45336 67364 45348
rect 67319 45308 67364 45336
rect 67358 45296 67364 45308
rect 67416 45296 67422 45348
rect 1104 45178 68816 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 65654 45178
rect 65706 45126 65718 45178
rect 65770 45126 65782 45178
rect 65834 45126 65846 45178
rect 65898 45126 65910 45178
rect 65962 45126 68816 45178
rect 1104 45104 68816 45126
rect 1104 44634 68816 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 68816 44634
rect 1104 44560 68816 44582
rect 1104 44090 68816 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 65654 44090
rect 65706 44038 65718 44090
rect 65770 44038 65782 44090
rect 65834 44038 65846 44090
rect 65898 44038 65910 44090
rect 65962 44038 68816 44090
rect 1104 44016 68816 44038
rect 1104 43546 68816 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 68816 43546
rect 1104 43472 68816 43494
rect 1104 43002 68816 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 65654 43002
rect 65706 42950 65718 43002
rect 65770 42950 65782 43002
rect 65834 42950 65846 43002
rect 65898 42950 65910 43002
rect 65962 42950 68816 43002
rect 1104 42928 68816 42950
rect 1104 42458 68816 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 68816 42458
rect 1104 42384 68816 42406
rect 1104 41914 68816 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 65654 41914
rect 65706 41862 65718 41914
rect 65770 41862 65782 41914
rect 65834 41862 65846 41914
rect 65898 41862 65910 41914
rect 65962 41862 68816 41914
rect 1104 41840 68816 41862
rect 67821 41599 67879 41605
rect 67821 41596 67833 41599
rect 67284 41568 67833 41596
rect 67284 41472 67312 41568
rect 67821 41565 67833 41568
rect 67867 41565 67879 41599
rect 67821 41559 67879 41565
rect 67266 41460 67272 41472
rect 67227 41432 67272 41460
rect 67266 41420 67272 41432
rect 67324 41420 67330 41472
rect 68002 41460 68008 41472
rect 67963 41432 68008 41460
rect 68002 41420 68008 41432
rect 68060 41420 68066 41472
rect 1104 41370 68816 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 68816 41370
rect 1104 41296 68816 41318
rect 1104 40826 68816 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 65654 40826
rect 65706 40774 65718 40826
rect 65770 40774 65782 40826
rect 65834 40774 65846 40826
rect 65898 40774 65910 40826
rect 65962 40774 68816 40826
rect 1104 40752 68816 40774
rect 1104 40282 68816 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 68816 40282
rect 1104 40208 68816 40230
rect 1104 39738 68816 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 65654 39738
rect 65706 39686 65718 39738
rect 65770 39686 65782 39738
rect 65834 39686 65846 39738
rect 65898 39686 65910 39738
rect 65962 39686 68816 39738
rect 1104 39664 68816 39686
rect 67361 39627 67419 39633
rect 67361 39593 67373 39627
rect 67407 39624 67419 39627
rect 67450 39624 67456 39636
rect 67407 39596 67456 39624
rect 67407 39593 67419 39596
rect 67361 39587 67419 39593
rect 67450 39584 67456 39596
rect 67508 39584 67514 39636
rect 67174 39420 67180 39432
rect 67135 39392 67180 39420
rect 67174 39380 67180 39392
rect 67232 39420 67238 39432
rect 67821 39423 67879 39429
rect 67821 39420 67833 39423
rect 67232 39392 67833 39420
rect 67232 39380 67238 39392
rect 67821 39389 67833 39392
rect 67867 39389 67879 39423
rect 67821 39383 67879 39389
rect 1104 39194 68816 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 68816 39194
rect 1104 39120 68816 39142
rect 1104 38650 68816 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 65654 38650
rect 65706 38598 65718 38650
rect 65770 38598 65782 38650
rect 65834 38598 65846 38650
rect 65898 38598 65910 38650
rect 65962 38598 68816 38650
rect 1104 38576 68816 38598
rect 1104 38106 68816 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 68816 38106
rect 1104 38032 68816 38054
rect 1104 37562 68816 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 65654 37562
rect 65706 37510 65718 37562
rect 65770 37510 65782 37562
rect 65834 37510 65846 37562
rect 65898 37510 65910 37562
rect 65962 37510 68816 37562
rect 1104 37488 68816 37510
rect 1104 37018 68816 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 68816 37018
rect 1104 36944 68816 36966
rect 1104 36474 68816 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 65654 36474
rect 65706 36422 65718 36474
rect 65770 36422 65782 36474
rect 65834 36422 65846 36474
rect 65898 36422 65910 36474
rect 65962 36422 68816 36474
rect 1104 36400 68816 36422
rect 1104 35930 68816 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 68816 35930
rect 1104 35856 68816 35878
rect 1104 35386 68816 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 65654 35386
rect 65706 35334 65718 35386
rect 65770 35334 65782 35386
rect 65834 35334 65846 35386
rect 65898 35334 65910 35386
rect 65962 35334 68816 35386
rect 1104 35312 68816 35334
rect 1104 34842 68816 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 68816 34842
rect 1104 34768 68816 34790
rect 27614 34388 27620 34400
rect 27575 34360 27620 34388
rect 27614 34348 27620 34360
rect 27672 34348 27678 34400
rect 1104 34298 68816 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 65654 34298
rect 65706 34246 65718 34298
rect 65770 34246 65782 34298
rect 65834 34246 65846 34298
rect 65898 34246 65910 34298
rect 65962 34246 68816 34298
rect 1104 34224 68816 34246
rect 26878 34076 26884 34128
rect 26936 34116 26942 34128
rect 29086 34116 29092 34128
rect 26936 34088 29092 34116
rect 26936 34076 26942 34088
rect 29086 34076 29092 34088
rect 29144 34076 29150 34128
rect 27246 34048 27252 34060
rect 26712 34020 27252 34048
rect 26712 33989 26740 34020
rect 27246 34008 27252 34020
rect 27304 34048 27310 34060
rect 27709 34051 27767 34057
rect 27709 34048 27721 34051
rect 27304 34020 27721 34048
rect 27304 34008 27310 34020
rect 27709 34017 27721 34020
rect 27755 34048 27767 34051
rect 27890 34048 27896 34060
rect 27755 34020 27896 34048
rect 27755 34017 27767 34020
rect 27709 34011 27767 34017
rect 27890 34008 27896 34020
rect 27948 34008 27954 34060
rect 28169 34051 28227 34057
rect 28169 34017 28181 34051
rect 28215 34048 28227 34051
rect 28994 34048 29000 34060
rect 28215 34020 29000 34048
rect 28215 34017 28227 34020
rect 28169 34011 28227 34017
rect 28994 34008 29000 34020
rect 29052 34008 29058 34060
rect 26697 33983 26755 33989
rect 26697 33949 26709 33983
rect 26743 33949 26755 33983
rect 26697 33943 26755 33949
rect 26878 33940 26884 33992
rect 26936 33980 26942 33992
rect 26973 33983 27031 33989
rect 26973 33980 26985 33983
rect 26936 33952 26985 33980
rect 26936 33940 26942 33952
rect 26973 33949 26985 33952
rect 27019 33949 27031 33983
rect 26973 33943 27031 33949
rect 27801 33983 27859 33989
rect 27801 33949 27813 33983
rect 27847 33949 27859 33983
rect 27801 33943 27859 33949
rect 26789 33915 26847 33921
rect 26789 33881 26801 33915
rect 26835 33912 26847 33915
rect 27062 33912 27068 33924
rect 26835 33884 27068 33912
rect 26835 33881 26847 33884
rect 26789 33875 26847 33881
rect 27062 33872 27068 33884
rect 27120 33912 27126 33924
rect 27816 33912 27844 33943
rect 67358 33940 67364 33992
rect 67416 33980 67422 33992
rect 67821 33983 67879 33989
rect 67821 33980 67833 33983
rect 67416 33952 67833 33980
rect 67416 33940 67422 33952
rect 67821 33949 67833 33952
rect 67867 33949 67879 33983
rect 67821 33943 67879 33949
rect 27120 33884 27844 33912
rect 27120 33872 27126 33884
rect 12894 33804 12900 33856
rect 12952 33844 12958 33856
rect 13173 33847 13231 33853
rect 13173 33844 13185 33847
rect 12952 33816 13185 33844
rect 12952 33804 12958 33816
rect 13173 33813 13185 33816
rect 13219 33813 13231 33847
rect 13173 33807 13231 33813
rect 27157 33847 27215 33853
rect 27157 33813 27169 33847
rect 27203 33844 27215 33847
rect 27430 33844 27436 33856
rect 27203 33816 27436 33844
rect 27203 33813 27215 33816
rect 27157 33807 27215 33813
rect 27430 33804 27436 33816
rect 27488 33804 27494 33856
rect 27614 33804 27620 33856
rect 27672 33844 27678 33856
rect 28166 33844 28172 33856
rect 27672 33816 28172 33844
rect 27672 33804 27678 33816
rect 28166 33804 28172 33816
rect 28224 33804 28230 33856
rect 28810 33844 28816 33856
rect 28771 33816 28816 33844
rect 28810 33804 28816 33816
rect 28868 33804 28874 33856
rect 68002 33844 68008 33856
rect 67963 33816 68008 33844
rect 68002 33804 68008 33816
rect 68060 33804 68066 33856
rect 1104 33754 68816 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 68816 33754
rect 1104 33680 68816 33702
rect 13170 33640 13176 33652
rect 13131 33612 13176 33640
rect 13170 33600 13176 33612
rect 13228 33600 13234 33652
rect 31202 33640 31208 33652
rect 24688 33612 31208 33640
rect 14274 33572 14280 33584
rect 13004 33544 14280 33572
rect 7466 33464 7472 33516
rect 7524 33504 7530 33516
rect 13004 33513 13032 33544
rect 14274 33532 14280 33544
rect 14332 33572 14338 33584
rect 14332 33544 14596 33572
rect 14332 33532 14338 33544
rect 8757 33507 8815 33513
rect 8757 33504 8769 33507
rect 7524 33476 8769 33504
rect 7524 33464 7530 33476
rect 8757 33473 8769 33476
rect 8803 33473 8815 33507
rect 8757 33467 8815 33473
rect 12989 33507 13047 33513
rect 12989 33473 13001 33507
rect 13035 33473 13047 33507
rect 13262 33504 13268 33516
rect 13223 33476 13268 33504
rect 12989 33467 13047 33473
rect 13262 33464 13268 33476
rect 13320 33464 13326 33516
rect 14568 33513 14596 33544
rect 13909 33507 13967 33513
rect 13909 33504 13921 33507
rect 13372 33476 13921 33504
rect 8849 33439 8907 33445
rect 8849 33405 8861 33439
rect 8895 33436 8907 33439
rect 12526 33436 12532 33448
rect 8895 33408 12532 33436
rect 8895 33405 8907 33408
rect 8849 33399 8907 33405
rect 12526 33396 12532 33408
rect 12584 33436 12590 33448
rect 13372 33436 13400 33476
rect 13909 33473 13921 33476
rect 13955 33473 13967 33507
rect 13909 33467 13967 33473
rect 14553 33507 14611 33513
rect 14553 33473 14565 33507
rect 14599 33473 14611 33507
rect 14553 33467 14611 33473
rect 14737 33507 14795 33513
rect 14737 33473 14749 33507
rect 14783 33504 14795 33507
rect 16206 33504 16212 33516
rect 14783 33476 16212 33504
rect 14783 33473 14795 33476
rect 14737 33467 14795 33473
rect 16206 33464 16212 33476
rect 16264 33464 16270 33516
rect 22186 33464 22192 33516
rect 22244 33504 22250 33516
rect 24688 33513 24716 33612
rect 31202 33600 31208 33612
rect 31260 33600 31266 33652
rect 32398 33640 32404 33652
rect 31726 33612 32404 33640
rect 28166 33532 28172 33584
rect 28224 33572 28230 33584
rect 28902 33572 28908 33584
rect 28224 33544 28269 33572
rect 28863 33544 28908 33572
rect 28224 33532 28230 33544
rect 28902 33532 28908 33544
rect 28960 33532 28966 33584
rect 29012 33544 29316 33572
rect 24029 33507 24087 33513
rect 24029 33504 24041 33507
rect 22244 33476 24041 33504
rect 22244 33464 22250 33476
rect 24029 33473 24041 33476
rect 24075 33504 24087 33507
rect 24673 33507 24731 33513
rect 24673 33504 24685 33507
rect 24075 33476 24685 33504
rect 24075 33473 24087 33476
rect 24029 33467 24087 33473
rect 24673 33473 24685 33476
rect 24719 33473 24731 33507
rect 25958 33504 25964 33516
rect 25919 33476 25964 33504
rect 24673 33467 24731 33473
rect 25958 33464 25964 33476
rect 26016 33464 26022 33516
rect 27157 33507 27215 33513
rect 27157 33504 27169 33507
rect 26068 33476 27169 33504
rect 12584 33408 13400 33436
rect 13725 33439 13783 33445
rect 12584 33396 12590 33408
rect 13725 33405 13737 33439
rect 13771 33405 13783 33439
rect 13725 33399 13783 33405
rect 9125 33371 9183 33377
rect 9125 33337 9137 33371
rect 9171 33368 9183 33371
rect 9766 33368 9772 33380
rect 9171 33340 9772 33368
rect 9171 33337 9183 33340
rect 9125 33331 9183 33337
rect 9766 33328 9772 33340
rect 9824 33328 9830 33380
rect 13170 33328 13176 33380
rect 13228 33368 13234 33380
rect 13740 33368 13768 33399
rect 23658 33396 23664 33448
rect 23716 33436 23722 33448
rect 26068 33445 26096 33476
rect 27157 33473 27169 33476
rect 27203 33473 27215 33507
rect 27157 33467 27215 33473
rect 27706 33464 27712 33516
rect 27764 33504 27770 33516
rect 27801 33507 27859 33513
rect 27801 33504 27813 33507
rect 27764 33476 27813 33504
rect 27764 33464 27770 33476
rect 27801 33473 27813 33476
rect 27847 33473 27859 33507
rect 27801 33467 27859 33473
rect 27891 33464 27897 33516
rect 27949 33513 27955 33516
rect 27949 33507 27997 33513
rect 27949 33473 27951 33507
rect 27985 33473 27997 33507
rect 28074 33504 28080 33516
rect 28035 33476 28080 33504
rect 27949 33467 27997 33473
rect 27949 33464 27955 33467
rect 28074 33464 28080 33476
rect 28132 33464 28138 33516
rect 28285 33507 28343 33513
rect 28285 33504 28297 33507
rect 28281 33473 28297 33504
rect 28331 33473 28343 33507
rect 28281 33467 28343 33473
rect 24581 33439 24639 33445
rect 24581 33436 24593 33439
rect 23716 33408 24593 33436
rect 23716 33396 23722 33408
rect 24581 33405 24593 33408
rect 24627 33405 24639 33439
rect 26053 33439 26111 33445
rect 26053 33436 26065 33439
rect 24581 33399 24639 33405
rect 25056 33408 26065 33436
rect 25056 33377 25084 33408
rect 26053 33405 26065 33408
rect 26099 33405 26111 33439
rect 26053 33399 26111 33405
rect 26973 33439 27031 33445
rect 26973 33405 26985 33439
rect 27019 33436 27031 33439
rect 27062 33436 27068 33448
rect 27019 33408 27068 33436
rect 27019 33405 27031 33408
rect 26973 33399 27031 33405
rect 27062 33396 27068 33408
rect 27120 33396 27126 33448
rect 28281 33436 28309 33467
rect 28442 33464 28448 33516
rect 28500 33504 28506 33516
rect 29012 33504 29040 33544
rect 28500 33476 29040 33504
rect 28500 33464 28506 33476
rect 29086 33464 29092 33516
rect 29144 33504 29150 33516
rect 29288 33504 29316 33544
rect 31726 33504 31754 33612
rect 32398 33600 32404 33612
rect 32456 33600 32462 33652
rect 29144 33476 29189 33504
rect 29288 33476 31754 33504
rect 29144 33464 29150 33476
rect 34514 33464 34520 33516
rect 34572 33504 34578 33516
rect 35161 33507 35219 33513
rect 35161 33504 35173 33507
rect 34572 33476 35173 33504
rect 34572 33464 34578 33476
rect 35161 33473 35173 33476
rect 35207 33473 35219 33507
rect 35342 33504 35348 33516
rect 35303 33476 35348 33504
rect 35161 33467 35219 33473
rect 35342 33464 35348 33476
rect 35400 33464 35406 33516
rect 28281 33408 28396 33436
rect 14553 33371 14611 33377
rect 14553 33368 14565 33371
rect 13228 33340 14565 33368
rect 13228 33328 13234 33340
rect 14553 33337 14565 33340
rect 14599 33337 14611 33371
rect 14553 33331 14611 33337
rect 25041 33371 25099 33377
rect 25041 33337 25053 33371
rect 25087 33337 25099 33371
rect 26326 33368 26332 33380
rect 26287 33340 26332 33368
rect 25041 33331 25099 33337
rect 26326 33328 26332 33340
rect 26384 33328 26390 33380
rect 27341 33371 27399 33377
rect 27341 33337 27353 33371
rect 27387 33368 27399 33371
rect 28074 33368 28080 33380
rect 27387 33340 28080 33368
rect 27387 33337 27399 33340
rect 27341 33331 27399 33337
rect 28074 33328 28080 33340
rect 28132 33368 28138 33380
rect 28258 33368 28264 33380
rect 28132 33340 28264 33368
rect 28132 33328 28138 33340
rect 28258 33328 28264 33340
rect 28316 33328 28322 33380
rect 11146 33260 11152 33312
rect 11204 33300 11210 33312
rect 12805 33303 12863 33309
rect 12805 33300 12817 33303
rect 11204 33272 12817 33300
rect 11204 33260 11210 33272
rect 12805 33269 12817 33272
rect 12851 33269 12863 33303
rect 14090 33300 14096 33312
rect 14051 33272 14096 33300
rect 12805 33263 12863 33269
rect 14090 33260 14096 33272
rect 14148 33260 14154 33312
rect 15289 33303 15347 33309
rect 15289 33269 15301 33303
rect 15335 33300 15347 33303
rect 16022 33300 16028 33312
rect 15335 33272 16028 33300
rect 15335 33269 15347 33272
rect 15289 33263 15347 33269
rect 16022 33260 16028 33272
rect 16080 33260 16086 33312
rect 26050 33260 26056 33312
rect 26108 33300 26114 33312
rect 28368 33300 28396 33408
rect 28810 33396 28816 33448
rect 28868 33436 28874 33448
rect 29365 33439 29423 33445
rect 29365 33436 29377 33439
rect 28868 33408 29377 33436
rect 28868 33396 28874 33408
rect 29365 33405 29377 33408
rect 29411 33436 29423 33439
rect 37277 33439 37335 33445
rect 37277 33436 37289 33439
rect 29411 33408 37289 33436
rect 29411 33405 29423 33408
rect 29365 33399 29423 33405
rect 37277 33405 37289 33408
rect 37323 33436 37335 33439
rect 37734 33436 37740 33448
rect 37323 33408 37740 33436
rect 37323 33405 37335 33408
rect 37277 33399 37335 33405
rect 37734 33396 37740 33408
rect 37792 33396 37798 33448
rect 28445 33371 28503 33377
rect 28445 33337 28457 33371
rect 28491 33368 28503 33371
rect 31110 33368 31116 33380
rect 28491 33340 31116 33368
rect 28491 33337 28503 33340
rect 28445 33331 28503 33337
rect 31110 33328 31116 33340
rect 31168 33328 31174 33380
rect 31202 33328 31208 33380
rect 31260 33368 31266 33380
rect 35894 33368 35900 33380
rect 31260 33340 35900 33368
rect 31260 33328 31266 33340
rect 35894 33328 35900 33340
rect 35952 33368 35958 33380
rect 35952 33340 35997 33368
rect 35952 33328 35958 33340
rect 29273 33303 29331 33309
rect 29273 33300 29285 33303
rect 26108 33272 29285 33300
rect 26108 33260 26114 33272
rect 29273 33269 29285 33272
rect 29319 33269 29331 33303
rect 29273 33263 29331 33269
rect 34514 33260 34520 33312
rect 34572 33300 34578 33312
rect 34609 33303 34667 33309
rect 34609 33300 34621 33303
rect 34572 33272 34621 33300
rect 34572 33260 34578 33272
rect 34609 33269 34621 33272
rect 34655 33269 34667 33303
rect 34609 33263 34667 33269
rect 35345 33303 35403 33309
rect 35345 33269 35357 33303
rect 35391 33300 35403 33303
rect 37182 33300 37188 33312
rect 35391 33272 37188 33300
rect 35391 33269 35403 33272
rect 35345 33263 35403 33269
rect 37182 33260 37188 33272
rect 37240 33260 37246 33312
rect 1104 33210 68816 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 65654 33210
rect 65706 33158 65718 33210
rect 65770 33158 65782 33210
rect 65834 33158 65846 33210
rect 65898 33158 65910 33210
rect 65962 33158 68816 33210
rect 1104 33136 68816 33158
rect 16206 33096 16212 33108
rect 16167 33068 16212 33096
rect 16206 33056 16212 33068
rect 16264 33056 16270 33108
rect 26050 33096 26056 33108
rect 26011 33068 26056 33096
rect 26050 33056 26056 33068
rect 26108 33056 26114 33108
rect 26789 33099 26847 33105
rect 26789 33065 26801 33099
rect 26835 33096 26847 33099
rect 27062 33096 27068 33108
rect 26835 33068 27068 33096
rect 26835 33065 26847 33068
rect 26789 33059 26847 33065
rect 27062 33056 27068 33068
rect 27120 33056 27126 33108
rect 34057 33099 34115 33105
rect 34057 33096 34069 33099
rect 27172 33068 34069 33096
rect 12526 33028 12532 33040
rect 12487 33000 12532 33028
rect 12526 32988 12532 33000
rect 12584 32988 12590 33040
rect 12894 32988 12900 33040
rect 12952 33028 12958 33040
rect 19334 33028 19340 33040
rect 12952 33000 16528 33028
rect 19247 33000 19340 33028
rect 12952 32988 12958 33000
rect 9766 32960 9772 32972
rect 9727 32932 9772 32960
rect 9766 32920 9772 32932
rect 9824 32920 9830 32972
rect 12986 32960 12992 32972
rect 12947 32932 12992 32960
rect 12986 32920 12992 32932
rect 13044 32920 13050 32972
rect 15105 32963 15163 32969
rect 15105 32960 15117 32963
rect 14292 32932 15117 32960
rect 14292 32904 14320 32932
rect 15105 32929 15117 32932
rect 15151 32929 15163 32963
rect 15105 32923 15163 32929
rect 9677 32895 9735 32901
rect 9677 32861 9689 32895
rect 9723 32892 9735 32895
rect 11146 32892 11152 32904
rect 9723 32864 11152 32892
rect 9723 32861 9735 32864
rect 9677 32855 9735 32861
rect 11146 32852 11152 32864
rect 11204 32852 11210 32904
rect 12894 32892 12900 32904
rect 12855 32864 12900 32892
rect 12894 32852 12900 32864
rect 12952 32852 12958 32904
rect 14274 32892 14280 32904
rect 14235 32864 14280 32892
rect 14274 32852 14280 32864
rect 14332 32852 14338 32904
rect 14458 32892 14464 32904
rect 14419 32864 14464 32892
rect 14458 32852 14464 32864
rect 14516 32852 14522 32904
rect 14553 32895 14611 32901
rect 14553 32861 14565 32895
rect 14599 32861 14611 32895
rect 15010 32892 15016 32904
rect 14971 32864 15016 32892
rect 14553 32855 14611 32861
rect 14568 32824 14596 32855
rect 15010 32852 15016 32864
rect 15068 32852 15074 32904
rect 15197 32895 15255 32901
rect 15197 32861 15209 32895
rect 15243 32892 15255 32895
rect 16390 32892 16396 32904
rect 15243 32864 16396 32892
rect 15243 32861 15255 32864
rect 15197 32855 15255 32861
rect 16390 32852 16396 32864
rect 16448 32852 16454 32904
rect 16022 32824 16028 32836
rect 14568 32796 16028 32824
rect 16022 32784 16028 32796
rect 16080 32784 16086 32836
rect 16500 32824 16528 33000
rect 19334 32988 19340 33000
rect 19392 33028 19398 33040
rect 27172 33028 27200 33068
rect 34057 33065 34069 33068
rect 34103 33065 34115 33099
rect 34057 33059 34115 33065
rect 19392 33000 24532 33028
rect 19392 32988 19398 33000
rect 16577 32963 16635 32969
rect 16577 32929 16589 32963
rect 16623 32929 16635 32963
rect 16577 32923 16635 32929
rect 21468 32932 22508 32960
rect 16592 32892 16620 32923
rect 17129 32895 17187 32901
rect 17129 32892 17141 32895
rect 16592 32864 17141 32892
rect 17129 32861 17141 32864
rect 17175 32892 17187 32895
rect 18049 32895 18107 32901
rect 18049 32892 18061 32895
rect 17175 32864 18061 32892
rect 17175 32861 17187 32864
rect 17129 32855 17187 32861
rect 18049 32861 18061 32864
rect 18095 32892 18107 32895
rect 19334 32892 19340 32904
rect 18095 32864 19340 32892
rect 18095 32861 18107 32864
rect 18049 32855 18107 32861
rect 19334 32852 19340 32864
rect 19392 32852 19398 32904
rect 21468 32824 21496 32932
rect 22186 32892 22192 32904
rect 22066 32864 22192 32892
rect 22066 32824 22094 32864
rect 22186 32852 22192 32864
rect 22244 32852 22250 32904
rect 16500 32796 21496 32824
rect 21560 32796 22094 32824
rect 10045 32759 10103 32765
rect 10045 32725 10057 32759
rect 10091 32756 10103 32759
rect 10226 32756 10232 32768
rect 10091 32728 10232 32756
rect 10091 32725 10103 32728
rect 10045 32719 10103 32725
rect 10226 32716 10232 32728
rect 10284 32716 10290 32768
rect 13814 32716 13820 32768
rect 13872 32756 13878 32768
rect 14093 32759 14151 32765
rect 14093 32756 14105 32759
rect 13872 32728 14105 32756
rect 13872 32716 13878 32728
rect 14093 32725 14105 32728
rect 14139 32725 14151 32759
rect 14093 32719 14151 32725
rect 15010 32716 15016 32768
rect 15068 32756 15074 32768
rect 15657 32759 15715 32765
rect 15657 32756 15669 32759
rect 15068 32728 15669 32756
rect 15068 32716 15074 32728
rect 15657 32725 15669 32728
rect 15703 32756 15715 32759
rect 18230 32756 18236 32768
rect 15703 32728 18236 32756
rect 15703 32725 15715 32728
rect 15657 32719 15715 32725
rect 18230 32716 18236 32728
rect 18288 32716 18294 32768
rect 20162 32716 20168 32768
rect 20220 32756 20226 32768
rect 21560 32765 21588 32796
rect 22480 32765 22508 32932
rect 24504 32892 24532 33000
rect 25148 33000 27200 33028
rect 27801 33031 27859 33037
rect 25148 32901 25176 33000
rect 27801 32997 27813 33031
rect 27847 32997 27859 33031
rect 27801 32991 27859 32997
rect 26326 32920 26332 32972
rect 26384 32960 26390 32972
rect 27341 32963 27399 32969
rect 27341 32960 27353 32963
rect 26384 32932 27353 32960
rect 26384 32920 26390 32932
rect 27341 32929 27353 32932
rect 27387 32929 27399 32963
rect 27341 32923 27399 32929
rect 24673 32895 24731 32901
rect 24673 32892 24685 32895
rect 24504 32864 24685 32892
rect 24673 32861 24685 32864
rect 24719 32892 24731 32895
rect 25133 32895 25191 32901
rect 25133 32892 25145 32895
rect 24719 32864 25145 32892
rect 24719 32861 24731 32864
rect 24673 32855 24731 32861
rect 25133 32861 25145 32864
rect 25179 32861 25191 32895
rect 25314 32892 25320 32904
rect 25275 32864 25320 32892
rect 25133 32855 25191 32861
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 25961 32895 26019 32901
rect 25961 32892 25973 32895
rect 25424 32864 25973 32892
rect 23658 32784 23664 32836
rect 23716 32824 23722 32836
rect 25424 32824 25452 32864
rect 25961 32861 25973 32864
rect 26007 32861 26019 32895
rect 25961 32855 26019 32861
rect 26605 32895 26663 32901
rect 26605 32861 26617 32895
rect 26651 32861 26663 32895
rect 26786 32892 26792 32904
rect 26747 32864 26792 32892
rect 26605 32855 26663 32861
rect 23716 32796 25452 32824
rect 25501 32827 25559 32833
rect 23716 32784 23722 32796
rect 25501 32793 25513 32827
rect 25547 32824 25559 32827
rect 26620 32824 26648 32855
rect 26786 32852 26792 32864
rect 26844 32852 26850 32904
rect 27430 32892 27436 32904
rect 27391 32864 27436 32892
rect 27430 32852 27436 32864
rect 27488 32852 27494 32904
rect 27816 32892 27844 32991
rect 28813 32963 28871 32969
rect 28813 32929 28825 32963
rect 28859 32960 28871 32963
rect 33134 32960 33140 32972
rect 28859 32932 33140 32960
rect 28859 32929 28871 32932
rect 28813 32923 28871 32929
rect 33134 32920 33140 32932
rect 33192 32920 33198 32972
rect 34072 32960 34100 33059
rect 35069 32963 35127 32969
rect 35069 32960 35081 32963
rect 34072 32932 35081 32960
rect 35069 32929 35081 32932
rect 35115 32929 35127 32963
rect 35069 32923 35127 32929
rect 36265 32963 36323 32969
rect 36265 32929 36277 32963
rect 36311 32960 36323 32963
rect 36538 32960 36544 32972
rect 36311 32932 36544 32960
rect 36311 32929 36323 32932
rect 36265 32923 36323 32929
rect 36538 32920 36544 32932
rect 36596 32920 36602 32972
rect 37093 32963 37151 32969
rect 37093 32929 37105 32963
rect 37139 32960 37151 32963
rect 38473 32963 38531 32969
rect 38473 32960 38485 32963
rect 37139 32932 38485 32960
rect 37139 32929 37151 32932
rect 37093 32923 37151 32929
rect 38473 32929 38485 32932
rect 38519 32960 38531 32963
rect 38654 32960 38660 32972
rect 38519 32932 38660 32960
rect 38519 32929 38531 32932
rect 38473 32923 38531 32929
rect 38654 32920 38660 32932
rect 38712 32920 38718 32972
rect 28261 32895 28319 32901
rect 28261 32892 28273 32895
rect 27816 32864 28273 32892
rect 28261 32861 28273 32864
rect 28307 32861 28319 32895
rect 28261 32855 28319 32861
rect 28350 32852 28356 32904
rect 28408 32892 28414 32904
rect 28537 32895 28595 32901
rect 28408 32864 28453 32892
rect 28408 32852 28414 32864
rect 28537 32861 28549 32895
rect 28583 32861 28595 32895
rect 28537 32855 28595 32861
rect 25547 32796 26648 32824
rect 28552 32824 28580 32855
rect 28626 32852 28632 32904
rect 28684 32892 28690 32904
rect 28684 32864 28729 32892
rect 28684 32852 28690 32864
rect 28994 32852 29000 32904
rect 29052 32892 29058 32904
rect 29549 32895 29607 32901
rect 29549 32892 29561 32895
rect 29052 32864 29561 32892
rect 29052 32852 29058 32864
rect 29549 32861 29561 32864
rect 29595 32861 29607 32895
rect 29730 32892 29736 32904
rect 29691 32864 29736 32892
rect 29549 32855 29607 32861
rect 29730 32852 29736 32864
rect 29788 32852 29794 32904
rect 32398 32892 32404 32904
rect 32359 32864 32404 32892
rect 32398 32852 32404 32864
rect 32456 32852 32462 32904
rect 35253 32895 35311 32901
rect 35253 32861 35265 32895
rect 35299 32892 35311 32895
rect 35342 32892 35348 32904
rect 35299 32864 35348 32892
rect 35299 32861 35311 32864
rect 35253 32855 35311 32861
rect 35342 32852 35348 32864
rect 35400 32852 35406 32904
rect 35894 32852 35900 32904
rect 35952 32892 35958 32904
rect 36173 32895 36231 32901
rect 36173 32892 36185 32895
rect 35952 32864 36185 32892
rect 35952 32852 35958 32864
rect 36173 32861 36185 32864
rect 36219 32861 36231 32895
rect 36173 32855 36231 32861
rect 37001 32895 37059 32901
rect 37001 32861 37013 32895
rect 37047 32861 37059 32895
rect 37182 32892 37188 32904
rect 37143 32864 37188 32892
rect 37001 32855 37059 32861
rect 29641 32827 29699 32833
rect 29641 32824 29653 32827
rect 28552 32796 29653 32824
rect 25547 32793 25559 32796
rect 25501 32787 25559 32793
rect 29641 32793 29653 32796
rect 29687 32793 29699 32827
rect 29641 32787 29699 32793
rect 35437 32827 35495 32833
rect 35437 32793 35449 32827
rect 35483 32824 35495 32827
rect 37016 32824 37044 32855
rect 37182 32852 37188 32864
rect 37240 32852 37246 32904
rect 38286 32892 38292 32904
rect 37752 32864 38292 32892
rect 35483 32796 37044 32824
rect 35483 32793 35495 32796
rect 35437 32787 35495 32793
rect 21545 32759 21603 32765
rect 21545 32756 21557 32759
rect 20220 32728 21557 32756
rect 20220 32716 20226 32728
rect 21545 32725 21557 32728
rect 21591 32725 21603 32759
rect 21545 32719 21603 32725
rect 22465 32759 22523 32765
rect 22465 32725 22477 32759
rect 22511 32756 22523 32759
rect 26418 32756 26424 32768
rect 22511 32728 26424 32756
rect 22511 32725 22523 32728
rect 22465 32719 22523 32725
rect 26418 32716 26424 32728
rect 26476 32716 26482 32768
rect 32493 32759 32551 32765
rect 32493 32725 32505 32759
rect 32539 32756 32551 32759
rect 33318 32756 33324 32768
rect 32539 32728 33324 32756
rect 32539 32725 32551 32728
rect 32493 32719 32551 32725
rect 33318 32716 33324 32728
rect 33376 32716 33382 32768
rect 36541 32759 36599 32765
rect 36541 32725 36553 32759
rect 36587 32756 36599 32759
rect 37752 32756 37780 32864
rect 38286 32852 38292 32864
rect 38344 32852 38350 32904
rect 36587 32728 37780 32756
rect 38105 32759 38163 32765
rect 36587 32725 36599 32728
rect 36541 32719 36599 32725
rect 38105 32725 38117 32759
rect 38151 32756 38163 32759
rect 38746 32756 38752 32768
rect 38151 32728 38752 32756
rect 38151 32725 38163 32728
rect 38105 32719 38163 32725
rect 38746 32716 38752 32728
rect 38804 32716 38810 32768
rect 1104 32666 68816 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 68816 32666
rect 1104 32592 68816 32614
rect 18230 32512 18236 32564
rect 18288 32552 18294 32564
rect 25409 32555 25467 32561
rect 18288 32524 22094 32552
rect 18288 32512 18294 32524
rect 14185 32487 14243 32493
rect 14185 32453 14197 32487
rect 14231 32484 14243 32487
rect 22066 32484 22094 32524
rect 25409 32521 25421 32555
rect 25455 32552 25467 32555
rect 26786 32552 26792 32564
rect 25455 32524 26792 32552
rect 25455 32521 25467 32524
rect 25409 32515 25467 32521
rect 26786 32512 26792 32524
rect 26844 32512 26850 32564
rect 28626 32552 28632 32564
rect 28587 32524 28632 32552
rect 28626 32512 28632 32524
rect 28684 32512 28690 32564
rect 34514 32552 34520 32564
rect 31726 32524 34520 32552
rect 24857 32487 24915 32493
rect 24857 32484 24869 32487
rect 14231 32456 16068 32484
rect 22066 32456 24869 32484
rect 14231 32453 14243 32456
rect 14185 32447 14243 32453
rect 16040 32428 16068 32456
rect 24857 32453 24869 32456
rect 24903 32484 24915 32487
rect 31726 32484 31754 32524
rect 34514 32512 34520 32524
rect 34572 32512 34578 32564
rect 38654 32552 38660 32564
rect 38615 32524 38660 32552
rect 38654 32512 38660 32524
rect 38712 32552 38718 32564
rect 38712 32524 39896 32552
rect 38712 32512 38718 32524
rect 24903 32456 31754 32484
rect 34609 32487 34667 32493
rect 24903 32453 24915 32456
rect 24857 32447 24915 32453
rect 6549 32419 6607 32425
rect 6549 32385 6561 32419
rect 6595 32416 6607 32419
rect 7098 32416 7104 32428
rect 6595 32388 7104 32416
rect 6595 32385 6607 32388
rect 6549 32379 6607 32385
rect 7098 32376 7104 32388
rect 7156 32376 7162 32428
rect 9030 32416 9036 32428
rect 8991 32388 9036 32416
rect 9030 32376 9036 32388
rect 9088 32376 9094 32428
rect 12713 32419 12771 32425
rect 12713 32385 12725 32419
rect 12759 32416 12771 32419
rect 13170 32416 13176 32428
rect 12759 32388 13176 32416
rect 12759 32385 12771 32388
rect 12713 32379 12771 32385
rect 13170 32376 13176 32388
rect 13228 32376 13234 32428
rect 13814 32416 13820 32428
rect 13775 32388 13820 32416
rect 13814 32376 13820 32388
rect 13872 32376 13878 32428
rect 13910 32419 13968 32425
rect 13910 32385 13922 32419
rect 13956 32385 13968 32419
rect 13910 32379 13968 32385
rect 9125 32351 9183 32357
rect 9125 32317 9137 32351
rect 9171 32317 9183 32351
rect 12802 32348 12808 32360
rect 12763 32320 12808 32348
rect 9125 32311 9183 32317
rect 9140 32280 9168 32311
rect 12802 32308 12808 32320
rect 12860 32348 12866 32360
rect 13262 32348 13268 32360
rect 12860 32320 13268 32348
rect 12860 32308 12866 32320
rect 13262 32308 13268 32320
rect 13320 32348 13326 32360
rect 13924 32348 13952 32379
rect 14090 32376 14096 32428
rect 14148 32416 14154 32428
rect 14323 32419 14381 32425
rect 14148 32388 14241 32416
rect 14148 32376 14154 32388
rect 14323 32385 14335 32419
rect 14369 32416 14381 32419
rect 14458 32416 14464 32428
rect 14369 32388 14464 32416
rect 14369 32385 14381 32388
rect 14323 32379 14381 32385
rect 14458 32376 14464 32388
rect 14516 32376 14522 32428
rect 15470 32416 15476 32428
rect 15431 32388 15476 32416
rect 15470 32376 15476 32388
rect 15528 32376 15534 32428
rect 16022 32416 16028 32428
rect 15935 32388 16028 32416
rect 16022 32376 16028 32388
rect 16080 32416 16086 32428
rect 18601 32419 18659 32425
rect 16080 32388 18000 32416
rect 16080 32376 16086 32388
rect 13320 32320 13952 32348
rect 14108 32348 14136 32376
rect 14734 32348 14740 32360
rect 14108 32320 14740 32348
rect 13320 32308 13326 32320
rect 14734 32308 14740 32320
rect 14792 32308 14798 32360
rect 17402 32308 17408 32360
rect 17460 32348 17466 32360
rect 17972 32357 18000 32388
rect 18601 32385 18613 32419
rect 18647 32416 18659 32419
rect 18690 32416 18696 32428
rect 18647 32388 18696 32416
rect 18647 32385 18659 32388
rect 18601 32379 18659 32385
rect 18690 32376 18696 32388
rect 18748 32376 18754 32428
rect 23198 32416 23204 32428
rect 23159 32388 23204 32416
rect 23198 32376 23204 32388
rect 23256 32376 23262 32428
rect 23382 32376 23388 32428
rect 23440 32416 23446 32428
rect 25314 32416 25320 32428
rect 23440 32388 25320 32416
rect 23440 32376 23446 32388
rect 25314 32376 25320 32388
rect 25372 32376 25378 32428
rect 25516 32425 25544 32456
rect 34609 32453 34621 32487
rect 34655 32484 34667 32487
rect 35342 32484 35348 32496
rect 34655 32456 35348 32484
rect 34655 32453 34667 32456
rect 34609 32447 34667 32453
rect 35342 32444 35348 32456
rect 35400 32444 35406 32496
rect 37476 32456 38700 32484
rect 25501 32419 25559 32425
rect 25501 32385 25513 32419
rect 25547 32385 25559 32419
rect 26418 32416 26424 32428
rect 26331 32388 26424 32416
rect 25501 32379 25559 32385
rect 26418 32376 26424 32388
rect 26476 32416 26482 32428
rect 27433 32419 27491 32425
rect 27433 32416 27445 32419
rect 26476 32388 27445 32416
rect 26476 32376 26482 32388
rect 27433 32385 27445 32388
rect 27479 32385 27491 32419
rect 27433 32379 27491 32385
rect 17681 32351 17739 32357
rect 17681 32348 17693 32351
rect 17460 32320 17693 32348
rect 17460 32308 17466 32320
rect 17681 32317 17693 32320
rect 17727 32317 17739 32351
rect 17681 32311 17739 32317
rect 17957 32351 18015 32357
rect 17957 32317 17969 32351
rect 18003 32317 18015 32351
rect 27448 32348 27476 32379
rect 27890 32376 27896 32428
rect 27948 32416 27954 32428
rect 28813 32419 28871 32425
rect 28813 32416 28825 32419
rect 27948 32388 28825 32416
rect 27948 32376 27954 32388
rect 28813 32385 28825 32388
rect 28859 32385 28871 32419
rect 28994 32416 29000 32428
rect 28955 32388 29000 32416
rect 28813 32379 28871 32385
rect 28718 32348 28724 32360
rect 27448 32320 28724 32348
rect 17957 32311 18015 32317
rect 12345 32283 12403 32289
rect 12345 32280 12357 32283
rect 9140 32252 12357 32280
rect 12345 32249 12357 32252
rect 12391 32249 12403 32283
rect 17972 32280 18000 32311
rect 28718 32308 28724 32320
rect 28776 32308 28782 32360
rect 28828 32348 28856 32379
rect 28994 32376 29000 32388
rect 29052 32376 29058 32428
rect 33505 32419 33563 32425
rect 33505 32385 33517 32419
rect 33551 32416 33563 32419
rect 34514 32416 34520 32428
rect 33551 32388 34192 32416
rect 34475 32388 34520 32416
rect 33551 32385 33563 32388
rect 33505 32379 33563 32385
rect 29730 32348 29736 32360
rect 28828 32320 29736 32348
rect 29730 32308 29736 32320
rect 29788 32308 29794 32360
rect 19153 32283 19211 32289
rect 19153 32280 19165 32283
rect 17972 32252 19165 32280
rect 12345 32243 12403 32249
rect 19153 32249 19165 32252
rect 19199 32280 19211 32283
rect 27614 32280 27620 32292
rect 19199 32252 27620 32280
rect 19199 32249 19211 32252
rect 19153 32243 19211 32249
rect 27614 32240 27620 32252
rect 27672 32240 27678 32292
rect 34164 32289 34192 32388
rect 34514 32376 34520 32388
rect 34572 32376 34578 32428
rect 35713 32419 35771 32425
rect 35713 32385 35725 32419
rect 35759 32416 35771 32419
rect 35802 32416 35808 32428
rect 35759 32388 35808 32416
rect 35759 32385 35771 32388
rect 35713 32379 35771 32385
rect 35802 32376 35808 32388
rect 35860 32376 35866 32428
rect 36538 32416 36544 32428
rect 36499 32388 36544 32416
rect 36538 32376 36544 32388
rect 36596 32376 36602 32428
rect 37182 32376 37188 32428
rect 37240 32416 37246 32428
rect 37476 32425 37504 32456
rect 37461 32419 37519 32425
rect 37461 32416 37473 32419
rect 37240 32388 37473 32416
rect 37240 32376 37246 32388
rect 37461 32385 37473 32388
rect 37507 32385 37519 32419
rect 37734 32416 37740 32428
rect 37695 32388 37740 32416
rect 37461 32379 37519 32385
rect 37734 32376 37740 32388
rect 37792 32376 37798 32428
rect 38565 32419 38623 32425
rect 38565 32385 38577 32419
rect 38611 32385 38623 32419
rect 38672 32416 38700 32456
rect 39868 32425 39896 32524
rect 38841 32419 38899 32425
rect 38841 32416 38853 32419
rect 38672 32388 38853 32416
rect 38565 32379 38623 32385
rect 38841 32385 38853 32388
rect 38887 32385 38899 32419
rect 38841 32379 38899 32385
rect 39853 32419 39911 32425
rect 39853 32385 39865 32419
rect 39899 32385 39911 32419
rect 39853 32379 39911 32385
rect 34793 32351 34851 32357
rect 34793 32317 34805 32351
rect 34839 32348 34851 32351
rect 35526 32348 35532 32360
rect 34839 32320 35532 32348
rect 34839 32317 34851 32320
rect 34793 32311 34851 32317
rect 35526 32308 35532 32320
rect 35584 32308 35590 32360
rect 35621 32351 35679 32357
rect 35621 32317 35633 32351
rect 35667 32348 35679 32351
rect 36556 32348 36584 32376
rect 35667 32320 36584 32348
rect 35667 32317 35679 32320
rect 35621 32311 35679 32317
rect 34149 32283 34207 32289
rect 34149 32249 34161 32283
rect 34195 32249 34207 32283
rect 34149 32243 34207 32249
rect 36633 32283 36691 32289
rect 36633 32249 36645 32283
rect 36679 32280 36691 32283
rect 37642 32280 37648 32292
rect 36679 32252 37648 32280
rect 36679 32249 36691 32252
rect 36633 32243 36691 32249
rect 37642 32240 37648 32252
rect 37700 32240 37706 32292
rect 38580 32280 38608 32379
rect 39945 32351 40003 32357
rect 39945 32317 39957 32351
rect 39991 32348 40003 32351
rect 40494 32348 40500 32360
rect 39991 32320 40500 32348
rect 39991 32317 40003 32320
rect 39945 32311 40003 32317
rect 39960 32280 39988 32311
rect 40494 32308 40500 32320
rect 40552 32308 40558 32360
rect 38580 32252 39988 32280
rect 6362 32212 6368 32224
rect 6323 32184 6368 32212
rect 6362 32172 6368 32184
rect 6420 32172 6426 32224
rect 9309 32215 9367 32221
rect 9309 32181 9321 32215
rect 9355 32212 9367 32215
rect 9674 32212 9680 32224
rect 9355 32184 9680 32212
rect 9355 32181 9367 32184
rect 9309 32175 9367 32181
rect 9674 32172 9680 32184
rect 9732 32172 9738 32224
rect 14274 32172 14280 32224
rect 14332 32212 14338 32224
rect 14461 32215 14519 32221
rect 14461 32212 14473 32215
rect 14332 32184 14473 32212
rect 14332 32172 14338 32184
rect 14461 32181 14473 32184
rect 14507 32181 14519 32215
rect 15286 32212 15292 32224
rect 15247 32184 15292 32212
rect 14461 32175 14519 32181
rect 15286 32172 15292 32184
rect 15344 32172 15350 32224
rect 17586 32172 17592 32224
rect 17644 32212 17650 32224
rect 18417 32215 18475 32221
rect 18417 32212 18429 32215
rect 17644 32184 18429 32212
rect 17644 32172 17650 32184
rect 18417 32181 18429 32184
rect 18463 32181 18475 32215
rect 18417 32175 18475 32181
rect 22738 32172 22744 32224
rect 22796 32212 22802 32224
rect 23017 32215 23075 32221
rect 23017 32212 23029 32215
rect 22796 32184 23029 32212
rect 22796 32172 22802 32184
rect 23017 32181 23029 32184
rect 23063 32181 23075 32215
rect 23017 32175 23075 32181
rect 33689 32215 33747 32221
rect 33689 32181 33701 32215
rect 33735 32212 33747 32215
rect 33962 32212 33968 32224
rect 33735 32184 33968 32212
rect 33735 32181 33747 32184
rect 33689 32175 33747 32181
rect 33962 32172 33968 32184
rect 34020 32172 34026 32224
rect 35894 32172 35900 32224
rect 35952 32212 35958 32224
rect 36081 32215 36139 32221
rect 36081 32212 36093 32215
rect 35952 32184 36093 32212
rect 35952 32172 35958 32184
rect 36081 32181 36093 32184
rect 36127 32181 36139 32215
rect 37274 32212 37280 32224
rect 37235 32184 37280 32212
rect 36081 32175 36139 32181
rect 37274 32172 37280 32184
rect 37332 32172 37338 32224
rect 37458 32172 37464 32224
rect 37516 32212 37522 32224
rect 38580 32212 38608 32252
rect 37516 32184 38608 32212
rect 39025 32215 39083 32221
rect 37516 32172 37522 32184
rect 39025 32181 39037 32215
rect 39071 32212 39083 32215
rect 40034 32212 40040 32224
rect 39071 32184 40040 32212
rect 39071 32181 39083 32184
rect 39025 32175 39083 32181
rect 40034 32172 40040 32184
rect 40092 32172 40098 32224
rect 40129 32215 40187 32221
rect 40129 32181 40141 32215
rect 40175 32212 40187 32215
rect 41138 32212 41144 32224
rect 40175 32184 41144 32212
rect 40175 32181 40187 32184
rect 40129 32175 40187 32181
rect 41138 32172 41144 32184
rect 41196 32172 41202 32224
rect 1104 32122 68816 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 65654 32122
rect 65706 32070 65718 32122
rect 65770 32070 65782 32122
rect 65834 32070 65846 32122
rect 65898 32070 65910 32122
rect 65962 32070 68816 32122
rect 1104 32048 68816 32070
rect 7098 32008 7104 32020
rect 7059 31980 7104 32008
rect 7098 31968 7104 31980
rect 7156 31968 7162 32020
rect 8389 32011 8447 32017
rect 8389 31977 8401 32011
rect 8435 32008 8447 32011
rect 8435 31980 12940 32008
rect 8435 31977 8447 31980
rect 8389 31971 8447 31977
rect 7006 31832 7012 31884
rect 7064 31872 7070 31884
rect 7653 31875 7711 31881
rect 7653 31872 7665 31875
rect 7064 31844 7665 31872
rect 7064 31832 7070 31844
rect 7653 31841 7665 31844
rect 7699 31841 7711 31875
rect 7653 31835 7711 31841
rect 5258 31804 5264 31816
rect 5219 31776 5264 31804
rect 5258 31764 5264 31776
rect 5316 31764 5322 31816
rect 7282 31764 7288 31816
rect 7340 31804 7346 31816
rect 7561 31807 7619 31813
rect 7561 31804 7573 31807
rect 7340 31776 7573 31804
rect 7340 31764 7346 31776
rect 7561 31773 7573 31776
rect 7607 31804 7619 31807
rect 8404 31804 8432 31971
rect 12912 31940 12940 31980
rect 12986 31968 12992 32020
rect 13044 32008 13050 32020
rect 13357 32011 13415 32017
rect 13357 32008 13369 32011
rect 13044 31980 13369 32008
rect 13044 31968 13050 31980
rect 13357 31977 13369 31980
rect 13403 32008 13415 32011
rect 13630 32008 13636 32020
rect 13403 31980 13636 32008
rect 13403 31977 13415 31980
rect 13357 31971 13415 31977
rect 13630 31968 13636 31980
rect 13688 31968 13694 32020
rect 14185 32011 14243 32017
rect 14185 31977 14197 32011
rect 14231 32008 14243 32011
rect 14458 32008 14464 32020
rect 14231 31980 14464 32008
rect 14231 31977 14243 31980
rect 14185 31971 14243 31977
rect 14458 31968 14464 31980
rect 14516 31968 14522 32020
rect 16390 32008 16396 32020
rect 14568 31980 15976 32008
rect 16351 31980 16396 32008
rect 14568 31940 14596 31980
rect 12912 31912 14596 31940
rect 15948 31940 15976 31980
rect 16390 31968 16396 31980
rect 16448 31968 16454 32020
rect 19334 32008 19340 32020
rect 19295 31980 19340 32008
rect 19334 31968 19340 31980
rect 19392 31968 19398 32020
rect 22005 32011 22063 32017
rect 22005 31977 22017 32011
rect 22051 32008 22063 32011
rect 22278 32008 22284 32020
rect 22051 31980 22284 32008
rect 22051 31977 22063 31980
rect 22005 31971 22063 31977
rect 22278 31968 22284 31980
rect 22336 32008 22342 32020
rect 23382 32008 23388 32020
rect 22336 31980 23388 32008
rect 22336 31968 22342 31980
rect 23382 31968 23388 31980
rect 23440 31968 23446 32020
rect 25777 32011 25835 32017
rect 25777 31977 25789 32011
rect 25823 32008 25835 32011
rect 25958 32008 25964 32020
rect 25823 31980 25964 32008
rect 25823 31977 25835 31980
rect 25777 31971 25835 31977
rect 25958 31968 25964 31980
rect 26016 31968 26022 32020
rect 27614 31968 27620 32020
rect 27672 32008 27678 32020
rect 36081 32011 36139 32017
rect 27672 31980 35894 32008
rect 27672 31968 27678 31980
rect 16574 31940 16580 31952
rect 15948 31912 16580 31940
rect 16574 31900 16580 31912
rect 16632 31900 16638 31952
rect 18693 31943 18751 31949
rect 18693 31909 18705 31943
rect 18739 31909 18751 31943
rect 18693 31903 18751 31909
rect 13004 31844 15056 31872
rect 7607 31776 8432 31804
rect 11977 31807 12035 31813
rect 7607 31773 7619 31776
rect 7561 31767 7619 31773
rect 11977 31773 11989 31807
rect 12023 31804 12035 31807
rect 12066 31804 12072 31816
rect 12023 31776 12072 31804
rect 12023 31773 12035 31776
rect 11977 31767 12035 31773
rect 12066 31764 12072 31776
rect 12124 31804 12130 31816
rect 13004 31804 13032 31844
rect 12124 31776 13032 31804
rect 12124 31764 12130 31776
rect 13630 31764 13636 31816
rect 13688 31804 13694 31816
rect 15028 31813 15056 31844
rect 14093 31807 14151 31813
rect 14093 31804 14105 31807
rect 13688 31776 14105 31804
rect 13688 31764 13694 31776
rect 14093 31773 14105 31776
rect 14139 31773 14151 31807
rect 14093 31767 14151 31773
rect 15013 31807 15071 31813
rect 15013 31773 15025 31807
rect 15059 31804 15071 31807
rect 17313 31807 17371 31813
rect 15059 31776 15424 31804
rect 15059 31773 15071 31776
rect 15013 31767 15071 31773
rect 15396 31748 15424 31776
rect 17313 31773 17325 31807
rect 17359 31804 17371 31807
rect 18138 31804 18144 31816
rect 17359 31776 18144 31804
rect 17359 31773 17371 31776
rect 17313 31767 17371 31773
rect 18138 31764 18144 31776
rect 18196 31764 18202 31816
rect 18708 31804 18736 31903
rect 23658 31900 23664 31952
rect 23716 31940 23722 31952
rect 23845 31943 23903 31949
rect 23845 31940 23857 31943
rect 23716 31912 23857 31940
rect 23716 31900 23722 31912
rect 23845 31909 23857 31912
rect 23891 31909 23903 31943
rect 23845 31903 23903 31909
rect 28353 31943 28411 31949
rect 28353 31909 28365 31943
rect 28399 31909 28411 31943
rect 35866 31940 35894 31980
rect 36081 31977 36093 32011
rect 36127 32008 36139 32011
rect 36538 32008 36544 32020
rect 36127 31980 36544 32008
rect 36127 31977 36139 31980
rect 36081 31971 36139 31977
rect 36538 31968 36544 31980
rect 36596 31968 36602 32020
rect 38654 32008 38660 32020
rect 37568 31980 38660 32008
rect 36446 31940 36452 31952
rect 35866 31912 36452 31940
rect 28353 31903 28411 31909
rect 27709 31875 27767 31881
rect 27709 31841 27721 31875
rect 27755 31841 27767 31875
rect 27890 31872 27896 31884
rect 27851 31844 27896 31872
rect 27709 31835 27767 31841
rect 19150 31804 19156 31816
rect 18708 31776 19156 31804
rect 19150 31764 19156 31776
rect 19208 31804 19214 31816
rect 19429 31807 19487 31813
rect 19429 31804 19441 31807
rect 19208 31776 19441 31804
rect 19208 31764 19214 31776
rect 19429 31773 19441 31776
rect 19475 31773 19487 31807
rect 20622 31804 20628 31816
rect 20583 31776 20628 31804
rect 19429 31767 19487 31773
rect 20622 31764 20628 31776
rect 20680 31804 20686 31816
rect 22465 31807 22523 31813
rect 22465 31804 22477 31807
rect 20680 31776 22477 31804
rect 20680 31764 20686 31776
rect 22465 31773 22477 31776
rect 22511 31804 22523 31807
rect 24397 31807 24455 31813
rect 24397 31804 24409 31807
rect 22511 31776 24409 31804
rect 22511 31773 22523 31776
rect 22465 31767 22523 31773
rect 5534 31745 5540 31748
rect 5528 31699 5540 31745
rect 5592 31736 5598 31748
rect 12244 31739 12302 31745
rect 5592 31708 5628 31736
rect 5534 31696 5540 31699
rect 5592 31696 5598 31708
rect 12244 31705 12256 31739
rect 12290 31736 12302 31739
rect 12618 31736 12624 31748
rect 12290 31708 12624 31736
rect 12290 31705 12302 31708
rect 12244 31699 12302 31705
rect 12618 31696 12624 31708
rect 12676 31696 12682 31748
rect 15286 31745 15292 31748
rect 15280 31736 15292 31745
rect 15247 31708 15292 31736
rect 15280 31699 15292 31708
rect 15286 31696 15292 31699
rect 15344 31696 15350 31748
rect 15378 31696 15384 31748
rect 15436 31696 15442 31748
rect 17586 31745 17592 31748
rect 17580 31699 17592 31745
rect 17644 31736 17650 31748
rect 20892 31739 20950 31745
rect 17644 31708 17680 31736
rect 17586 31696 17592 31699
rect 17644 31696 17650 31708
rect 20892 31705 20904 31739
rect 20938 31736 20950 31739
rect 20990 31736 20996 31748
rect 20938 31708 20996 31736
rect 20938 31705 20950 31708
rect 20892 31699 20950 31705
rect 20990 31696 20996 31708
rect 21048 31696 21054 31748
rect 22738 31745 22744 31748
rect 22732 31699 22744 31745
rect 22796 31736 22802 31748
rect 24044 31736 24072 31776
rect 24397 31773 24409 31776
rect 24443 31773 24455 31807
rect 24397 31767 24455 31773
rect 24302 31736 24308 31748
rect 22796 31708 22832 31736
rect 24044 31708 24308 31736
rect 22738 31696 22744 31699
rect 22796 31696 22802 31708
rect 24302 31696 24308 31708
rect 24360 31696 24366 31748
rect 24486 31696 24492 31748
rect 24544 31736 24550 31748
rect 24642 31739 24700 31745
rect 24642 31736 24654 31739
rect 24544 31708 24654 31736
rect 24544 31696 24550 31708
rect 24642 31705 24654 31708
rect 24688 31705 24700 31739
rect 24642 31699 24700 31705
rect 27430 31696 27436 31748
rect 27488 31736 27494 31748
rect 27724 31736 27752 31835
rect 27890 31832 27896 31844
rect 27948 31832 27954 31884
rect 28368 31804 28396 31903
rect 36446 31900 36452 31912
rect 36504 31900 36510 31952
rect 28997 31807 29055 31813
rect 28997 31804 29009 31807
rect 28368 31776 29009 31804
rect 28997 31773 29009 31776
rect 29043 31773 29055 31807
rect 28997 31767 29055 31773
rect 31205 31807 31263 31813
rect 31205 31773 31217 31807
rect 31251 31804 31263 31807
rect 34698 31804 34704 31816
rect 31251 31776 34704 31804
rect 31251 31773 31263 31776
rect 31205 31767 31263 31773
rect 34698 31764 34704 31776
rect 34756 31764 34762 31816
rect 37274 31804 37280 31816
rect 37235 31776 37280 31804
rect 37274 31764 37280 31776
rect 37332 31764 37338 31816
rect 37458 31813 37464 31816
rect 37425 31807 37464 31813
rect 37425 31773 37437 31807
rect 37425 31767 37464 31773
rect 37458 31764 37464 31767
rect 37516 31764 37522 31816
rect 37568 31813 37596 31980
rect 38654 31968 38660 31980
rect 38712 31968 38718 32020
rect 37921 31943 37979 31949
rect 37921 31909 37933 31943
rect 37967 31940 37979 31943
rect 38194 31940 38200 31952
rect 37967 31912 38200 31940
rect 37967 31909 37979 31912
rect 37921 31903 37979 31909
rect 38194 31900 38200 31912
rect 38252 31900 38258 31952
rect 38933 31943 38991 31949
rect 38933 31909 38945 31943
rect 38979 31940 38991 31943
rect 57885 31943 57943 31949
rect 38979 31912 39988 31940
rect 38979 31909 38991 31912
rect 38933 31903 38991 31909
rect 37642 31832 37648 31884
rect 37700 31832 37706 31884
rect 38286 31832 38292 31884
rect 38344 31872 38350 31884
rect 39960 31881 39988 31912
rect 57885 31909 57897 31943
rect 57931 31940 57943 31943
rect 67266 31940 67272 31952
rect 57931 31912 67272 31940
rect 57931 31909 57943 31912
rect 57885 31903 57943 31909
rect 67266 31900 67272 31912
rect 67324 31900 67330 31952
rect 38473 31875 38531 31881
rect 38473 31872 38485 31875
rect 38344 31844 38485 31872
rect 38344 31832 38350 31844
rect 38473 31841 38485 31844
rect 38519 31841 38531 31875
rect 38473 31835 38531 31841
rect 39945 31875 40003 31881
rect 39945 31841 39957 31875
rect 39991 31841 40003 31875
rect 41138 31872 41144 31884
rect 41099 31844 41144 31872
rect 39945 31835 40003 31841
rect 41138 31832 41144 31844
rect 41196 31832 41202 31884
rect 37553 31807 37611 31813
rect 37553 31773 37565 31807
rect 37599 31773 37611 31807
rect 37660 31804 37688 31832
rect 37742 31807 37800 31813
rect 37742 31804 37754 31807
rect 37660 31776 37754 31804
rect 37553 31767 37611 31773
rect 37742 31773 37754 31776
rect 37788 31773 37800 31807
rect 38562 31804 38568 31816
rect 38523 31776 38568 31804
rect 37742 31767 37800 31773
rect 38562 31764 38568 31776
rect 38620 31764 38626 31816
rect 40034 31804 40040 31816
rect 39995 31776 40040 31804
rect 40034 31764 40040 31776
rect 40092 31764 40098 31816
rect 41230 31804 41236 31816
rect 41191 31776 41236 31804
rect 41230 31764 41236 31776
rect 41288 31764 41294 31816
rect 41874 31804 41880 31816
rect 41835 31776 41880 31804
rect 41874 31764 41880 31776
rect 41932 31764 41938 31816
rect 57698 31804 57704 31816
rect 57659 31776 57704 31804
rect 57698 31764 57704 31776
rect 57756 31804 57762 31816
rect 58345 31807 58403 31813
rect 58345 31804 58357 31807
rect 57756 31776 58357 31804
rect 57756 31764 57762 31776
rect 58345 31773 58357 31776
rect 58391 31773 58403 31807
rect 58345 31767 58403 31773
rect 31478 31745 31484 31748
rect 27488 31708 27752 31736
rect 27488 31696 27494 31708
rect 31472 31699 31484 31745
rect 31536 31736 31542 31748
rect 34968 31739 35026 31745
rect 31536 31708 31572 31736
rect 31478 31696 31484 31699
rect 31536 31696 31542 31708
rect 34968 31705 34980 31739
rect 35014 31736 35026 31739
rect 35710 31736 35716 31748
rect 35014 31708 35716 31736
rect 35014 31705 35026 31708
rect 34968 31699 35026 31705
rect 35710 31696 35716 31708
rect 35768 31696 35774 31748
rect 36446 31696 36452 31748
rect 36504 31736 36510 31748
rect 37645 31739 37703 31745
rect 37645 31736 37657 31739
rect 36504 31708 37657 31736
rect 36504 31696 36510 31708
rect 37645 31705 37657 31708
rect 37691 31705 37703 31739
rect 37645 31699 37703 31705
rect 5626 31628 5632 31680
rect 5684 31668 5690 31680
rect 6454 31668 6460 31680
rect 5684 31640 6460 31668
rect 5684 31628 5690 31640
rect 6454 31628 6460 31640
rect 6512 31668 6518 31680
rect 6641 31671 6699 31677
rect 6641 31668 6653 31671
rect 6512 31640 6653 31668
rect 6512 31628 6518 31640
rect 6641 31637 6653 31640
rect 6687 31637 6699 31671
rect 7466 31668 7472 31680
rect 7427 31640 7472 31668
rect 6641 31631 6699 31637
rect 7466 31628 7472 31640
rect 7524 31628 7530 31680
rect 19978 31668 19984 31680
rect 19939 31640 19984 31668
rect 19978 31628 19984 31640
rect 20036 31628 20042 31680
rect 22186 31628 22192 31680
rect 22244 31668 22250 31680
rect 27157 31671 27215 31677
rect 27157 31668 27169 31671
rect 22244 31640 27169 31668
rect 22244 31628 22250 31640
rect 27157 31637 27169 31640
rect 27203 31668 27215 31671
rect 27985 31671 28043 31677
rect 27985 31668 27997 31671
rect 27203 31640 27997 31668
rect 27203 31637 27215 31640
rect 27157 31631 27215 31637
rect 27985 31637 27997 31640
rect 28031 31668 28043 31671
rect 28442 31668 28448 31680
rect 28031 31640 28448 31668
rect 28031 31637 28043 31640
rect 27985 31631 28043 31637
rect 28442 31628 28448 31640
rect 28500 31628 28506 31680
rect 28810 31668 28816 31680
rect 28771 31640 28816 31668
rect 28810 31628 28816 31640
rect 28868 31628 28874 31680
rect 32306 31628 32312 31680
rect 32364 31668 32370 31680
rect 32585 31671 32643 31677
rect 32585 31668 32597 31671
rect 32364 31640 32597 31668
rect 32364 31628 32370 31640
rect 32585 31637 32597 31640
rect 32631 31637 32643 31671
rect 32585 31631 32643 31637
rect 34057 31671 34115 31677
rect 34057 31637 34069 31671
rect 34103 31668 34115 31671
rect 34514 31668 34520 31680
rect 34103 31640 34520 31668
rect 34103 31637 34115 31640
rect 34057 31631 34115 31637
rect 34514 31628 34520 31640
rect 34572 31628 34578 31680
rect 35802 31628 35808 31680
rect 35860 31668 35866 31680
rect 36541 31671 36599 31677
rect 36541 31668 36553 31671
rect 35860 31640 36553 31668
rect 35860 31628 35866 31640
rect 36541 31637 36553 31640
rect 36587 31637 36599 31671
rect 40402 31668 40408 31680
rect 40363 31640 40408 31668
rect 36541 31631 36599 31637
rect 40402 31628 40408 31640
rect 40460 31628 40466 31680
rect 40862 31668 40868 31680
rect 40823 31640 40868 31668
rect 40862 31628 40868 31640
rect 40920 31628 40926 31680
rect 42058 31668 42064 31680
rect 42019 31640 42064 31668
rect 42058 31628 42064 31640
rect 42116 31628 42122 31680
rect 1104 31578 68816 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 68816 31578
rect 1104 31504 68816 31526
rect 5445 31467 5503 31473
rect 5445 31433 5457 31467
rect 5491 31464 5503 31467
rect 5626 31464 5632 31476
rect 5491 31436 5632 31464
rect 5491 31433 5503 31436
rect 5445 31427 5503 31433
rect 5626 31424 5632 31436
rect 5684 31424 5690 31476
rect 7098 31464 7104 31476
rect 5736 31436 7104 31464
rect 5736 31269 5764 31436
rect 7098 31424 7104 31436
rect 7156 31424 7162 31476
rect 8205 31467 8263 31473
rect 8205 31433 8217 31467
rect 8251 31433 8263 31467
rect 12618 31464 12624 31476
rect 12579 31436 12624 31464
rect 8205 31427 8263 31433
rect 6632 31399 6690 31405
rect 6632 31365 6644 31399
rect 6678 31396 6690 31399
rect 8220 31396 8248 31427
rect 12618 31424 12624 31436
rect 12676 31424 12682 31476
rect 13265 31467 13323 31473
rect 13265 31433 13277 31467
rect 13311 31433 13323 31467
rect 13630 31464 13636 31476
rect 13591 31436 13636 31464
rect 13265 31427 13323 31433
rect 6678 31368 8248 31396
rect 6678 31365 6690 31368
rect 6632 31359 6690 31365
rect 6454 31288 6460 31340
rect 6512 31328 6518 31340
rect 8386 31328 8392 31340
rect 6512 31300 7420 31328
rect 8347 31300 8392 31328
rect 6512 31288 6518 31300
rect 5537 31263 5595 31269
rect 5537 31260 5549 31263
rect 5368 31232 5549 31260
rect 4617 31195 4675 31201
rect 4617 31161 4629 31195
rect 4663 31192 4675 31195
rect 5368 31192 5396 31232
rect 5537 31229 5549 31232
rect 5583 31229 5595 31263
rect 5537 31223 5595 31229
rect 5721 31263 5779 31269
rect 5721 31229 5733 31263
rect 5767 31229 5779 31263
rect 5721 31223 5779 31229
rect 6365 31263 6423 31269
rect 6365 31229 6377 31263
rect 6411 31229 6423 31263
rect 7392 31260 7420 31300
rect 8386 31288 8392 31300
rect 8444 31288 8450 31340
rect 9125 31331 9183 31337
rect 9125 31297 9137 31331
rect 9171 31297 9183 31331
rect 9766 31328 9772 31340
rect 9125 31291 9183 31297
rect 9232 31300 9772 31328
rect 9140 31260 9168 31291
rect 9232 31269 9260 31300
rect 9766 31288 9772 31300
rect 9824 31288 9830 31340
rect 9950 31328 9956 31340
rect 9911 31300 9956 31328
rect 9950 31288 9956 31300
rect 10008 31288 10014 31340
rect 10226 31328 10232 31340
rect 10187 31300 10232 31328
rect 10226 31288 10232 31300
rect 10284 31288 10290 31340
rect 12805 31331 12863 31337
rect 12805 31297 12817 31331
rect 12851 31328 12863 31331
rect 13280 31328 13308 31427
rect 13630 31424 13636 31436
rect 13688 31424 13694 31476
rect 15381 31467 15439 31473
rect 15381 31433 15393 31467
rect 15427 31464 15439 31467
rect 15470 31464 15476 31476
rect 15427 31436 15476 31464
rect 15427 31433 15439 31436
rect 15381 31427 15439 31433
rect 15470 31424 15476 31436
rect 15528 31424 15534 31476
rect 15749 31467 15807 31473
rect 15749 31433 15761 31467
rect 15795 31464 15807 31467
rect 16390 31464 16396 31476
rect 15795 31436 16396 31464
rect 15795 31433 15807 31436
rect 15749 31427 15807 31433
rect 16390 31424 16396 31436
rect 16448 31424 16454 31476
rect 17218 31424 17224 31476
rect 17276 31464 17282 31476
rect 17313 31467 17371 31473
rect 17313 31464 17325 31467
rect 17276 31436 17325 31464
rect 17276 31424 17282 31436
rect 17313 31433 17325 31436
rect 17359 31464 17371 31467
rect 17402 31464 17408 31476
rect 17359 31436 17408 31464
rect 17359 31433 17371 31436
rect 17313 31427 17371 31433
rect 17402 31424 17408 31436
rect 17460 31424 17466 31476
rect 19521 31467 19579 31473
rect 19521 31433 19533 31467
rect 19567 31464 19579 31467
rect 20162 31464 20168 31476
rect 19567 31436 20168 31464
rect 19567 31433 19579 31436
rect 19521 31427 19579 31433
rect 20162 31424 20168 31436
rect 20220 31424 20226 31476
rect 20990 31464 20996 31476
rect 20951 31436 20996 31464
rect 20990 31424 20996 31436
rect 21048 31424 21054 31476
rect 21821 31467 21879 31473
rect 21821 31433 21833 31467
rect 21867 31433 21879 31467
rect 22278 31464 22284 31476
rect 22239 31436 22284 31464
rect 21821 31427 21879 31433
rect 17034 31328 17040 31340
rect 12851 31300 13308 31328
rect 15856 31300 17040 31328
rect 12851 31297 12863 31300
rect 12805 31291 12863 31297
rect 7392 31232 9168 31260
rect 9217 31263 9275 31269
rect 6365 31223 6423 31229
rect 9217 31229 9229 31263
rect 9263 31229 9275 31263
rect 10045 31263 10103 31269
rect 10045 31260 10057 31263
rect 9217 31223 9275 31229
rect 9508 31232 10057 31260
rect 4663 31164 5396 31192
rect 4663 31161 4675 31164
rect 4617 31155 4675 31161
rect 5077 31127 5135 31133
rect 5077 31093 5089 31127
rect 5123 31124 5135 31127
rect 5166 31124 5172 31136
rect 5123 31096 5172 31124
rect 5123 31093 5135 31096
rect 5077 31087 5135 31093
rect 5166 31084 5172 31096
rect 5224 31084 5230 31136
rect 5368 31124 5396 31164
rect 5442 31152 5448 31204
rect 5500 31192 5506 31204
rect 6380 31192 6408 31223
rect 5500 31164 6408 31192
rect 7745 31195 7803 31201
rect 5500 31152 5506 31164
rect 7745 31161 7757 31195
rect 7791 31192 7803 31195
rect 8294 31192 8300 31204
rect 7791 31164 8300 31192
rect 7791 31161 7803 31164
rect 7745 31155 7803 31161
rect 8294 31152 8300 31164
rect 8352 31192 8358 31204
rect 9030 31192 9036 31204
rect 8352 31164 9036 31192
rect 8352 31152 8358 31164
rect 9030 31152 9036 31164
rect 9088 31152 9094 31204
rect 9508 31201 9536 31232
rect 10045 31229 10057 31232
rect 10091 31229 10103 31263
rect 13722 31260 13728 31272
rect 13683 31232 13728 31260
rect 10045 31223 10103 31229
rect 13722 31220 13728 31232
rect 13780 31220 13786 31272
rect 13814 31220 13820 31272
rect 13872 31260 13878 31272
rect 13872 31232 13917 31260
rect 13872 31220 13878 31232
rect 14918 31220 14924 31272
rect 14976 31260 14982 31272
rect 15856 31269 15884 31300
rect 17034 31288 17040 31300
rect 17092 31288 17098 31340
rect 18141 31331 18199 31337
rect 18141 31297 18153 31331
rect 18187 31328 18199 31331
rect 18230 31328 18236 31340
rect 18187 31300 18236 31328
rect 18187 31297 18199 31300
rect 18141 31291 18199 31297
rect 18230 31288 18236 31300
rect 18288 31288 18294 31340
rect 18414 31337 18420 31340
rect 18408 31291 18420 31337
rect 18472 31328 18478 31340
rect 18472 31300 18508 31328
rect 18414 31288 18420 31291
rect 18472 31288 18478 31300
rect 18966 31288 18972 31340
rect 19024 31328 19030 31340
rect 19978 31328 19984 31340
rect 19024 31300 19984 31328
rect 19024 31288 19030 31300
rect 19978 31288 19984 31300
rect 20036 31328 20042 31340
rect 20165 31331 20223 31337
rect 20165 31328 20177 31331
rect 20036 31300 20177 31328
rect 20036 31288 20042 31300
rect 20165 31297 20177 31300
rect 20211 31297 20223 31331
rect 20165 31291 20223 31297
rect 21177 31331 21235 31337
rect 21177 31297 21189 31331
rect 21223 31328 21235 31331
rect 21836 31328 21864 31427
rect 22278 31424 22284 31436
rect 22336 31424 22342 31476
rect 23198 31464 23204 31476
rect 23159 31436 23204 31464
rect 23198 31424 23204 31436
rect 23256 31424 23262 31476
rect 23658 31464 23664 31476
rect 23619 31436 23664 31464
rect 23658 31424 23664 31436
rect 23716 31424 23722 31476
rect 24486 31464 24492 31476
rect 24447 31436 24492 31464
rect 24486 31424 24492 31436
rect 24544 31424 24550 31476
rect 25133 31467 25191 31473
rect 25133 31433 25145 31467
rect 25179 31433 25191 31467
rect 25133 31427 25191 31433
rect 25593 31467 25651 31473
rect 25593 31433 25605 31467
rect 25639 31464 25651 31467
rect 25958 31464 25964 31476
rect 25639 31436 25964 31464
rect 25639 31433 25651 31436
rect 25593 31427 25651 31433
rect 22186 31396 22192 31408
rect 21223 31300 21864 31328
rect 22066 31368 22192 31396
rect 21223 31297 21235 31300
rect 21177 31291 21235 31297
rect 15841 31263 15899 31269
rect 15841 31260 15853 31263
rect 14976 31232 15853 31260
rect 14976 31220 14982 31232
rect 15841 31229 15853 31232
rect 15887 31229 15899 31263
rect 15841 31223 15899 31229
rect 15933 31263 15991 31269
rect 15933 31229 15945 31263
rect 15979 31229 15991 31263
rect 17126 31260 17132 31272
rect 17087 31232 17132 31260
rect 15933 31223 15991 31229
rect 9493 31195 9551 31201
rect 9493 31161 9505 31195
rect 9539 31161 9551 31195
rect 13832 31192 13860 31220
rect 15948 31192 15976 31223
rect 17126 31220 17132 31232
rect 17184 31220 17190 31272
rect 17221 31263 17279 31269
rect 17221 31229 17233 31263
rect 17267 31229 17279 31263
rect 17221 31223 17279 31229
rect 13832 31164 15976 31192
rect 9493 31155 9551 31161
rect 16942 31152 16948 31204
rect 17000 31192 17006 31204
rect 17236 31192 17264 31223
rect 17000 31164 17264 31192
rect 20349 31195 20407 31201
rect 17000 31152 17006 31164
rect 20349 31161 20361 31195
rect 20395 31192 20407 31195
rect 22066 31192 22094 31368
rect 22186 31356 22192 31368
rect 22244 31356 22250 31408
rect 23569 31331 23627 31337
rect 23569 31297 23581 31331
rect 23615 31328 23627 31331
rect 24673 31331 24731 31337
rect 23615 31300 24624 31328
rect 23615 31297 23627 31300
rect 23569 31291 23627 31297
rect 22465 31263 22523 31269
rect 22465 31229 22477 31263
rect 22511 31260 22523 31263
rect 22738 31260 22744 31272
rect 22511 31232 22744 31260
rect 22511 31229 22523 31232
rect 22465 31223 22523 31229
rect 22738 31220 22744 31232
rect 22796 31260 22802 31272
rect 23753 31263 23811 31269
rect 23753 31260 23765 31263
rect 22796 31232 23765 31260
rect 22796 31220 22802 31232
rect 23753 31229 23765 31232
rect 23799 31229 23811 31263
rect 24596 31260 24624 31300
rect 24673 31297 24685 31331
rect 24719 31328 24731 31331
rect 25148 31328 25176 31427
rect 25958 31424 25964 31436
rect 26016 31424 26022 31476
rect 27525 31467 27583 31473
rect 27525 31433 27537 31467
rect 27571 31464 27583 31467
rect 28350 31464 28356 31476
rect 27571 31436 28356 31464
rect 27571 31433 27583 31436
rect 27525 31427 27583 31433
rect 28350 31424 28356 31436
rect 28408 31424 28414 31476
rect 28442 31424 28448 31476
rect 28500 31464 28506 31476
rect 29730 31464 29736 31476
rect 28500 31436 28948 31464
rect 29691 31436 29736 31464
rect 28500 31424 28506 31436
rect 28620 31399 28678 31405
rect 28620 31365 28632 31399
rect 28666 31396 28678 31399
rect 28810 31396 28816 31408
rect 28666 31368 28816 31396
rect 28666 31365 28678 31368
rect 28620 31359 28678 31365
rect 28810 31356 28816 31368
rect 28868 31356 28874 31408
rect 28920 31396 28948 31436
rect 29730 31424 29736 31436
rect 29788 31424 29794 31476
rect 31389 31467 31447 31473
rect 31389 31433 31401 31467
rect 31435 31464 31447 31467
rect 31478 31464 31484 31476
rect 31435 31436 31484 31464
rect 31435 31433 31447 31436
rect 31389 31427 31447 31433
rect 31478 31424 31484 31436
rect 31536 31424 31542 31476
rect 32493 31467 32551 31473
rect 32493 31433 32505 31467
rect 32539 31464 32551 31467
rect 33413 31467 33471 31473
rect 33413 31464 33425 31467
rect 32539 31436 33425 31464
rect 32539 31433 32551 31436
rect 32493 31427 32551 31433
rect 33413 31433 33425 31436
rect 33459 31464 33471 31467
rect 34514 31464 34520 31476
rect 33459 31436 34520 31464
rect 33459 31433 33471 31436
rect 33413 31427 33471 31433
rect 32508 31396 32536 31427
rect 34514 31424 34520 31436
rect 34572 31464 34578 31476
rect 35253 31467 35311 31473
rect 34572 31436 34836 31464
rect 34572 31424 34578 31436
rect 34698 31396 34704 31408
rect 28920 31368 32536 31396
rect 33888 31368 34704 31396
rect 25498 31328 25504 31340
rect 24719 31300 25176 31328
rect 25459 31300 25504 31328
rect 24719 31297 24731 31300
rect 24673 31291 24731 31297
rect 25498 31288 25504 31300
rect 25556 31288 25562 31340
rect 27154 31328 27160 31340
rect 27115 31300 27160 31328
rect 27154 31288 27160 31300
rect 27212 31288 27218 31340
rect 31573 31331 31631 31337
rect 31573 31297 31585 31331
rect 31619 31328 31631 31331
rect 31619 31300 31754 31328
rect 31619 31297 31631 31300
rect 31573 31291 31631 31297
rect 25516 31260 25544 31288
rect 24596 31232 25544 31260
rect 25685 31263 25743 31269
rect 23753 31223 23811 31229
rect 25685 31229 25697 31263
rect 25731 31229 25743 31263
rect 25685 31223 25743 31229
rect 20395 31164 22094 31192
rect 25700 31192 25728 31223
rect 25774 31220 25780 31272
rect 25832 31260 25838 31272
rect 27065 31263 27123 31269
rect 27065 31260 27077 31263
rect 25832 31232 27077 31260
rect 25832 31220 25838 31232
rect 27065 31229 27077 31232
rect 27111 31229 27123 31263
rect 28350 31260 28356 31272
rect 28311 31232 28356 31260
rect 27065 31223 27123 31229
rect 28350 31220 28356 31232
rect 28408 31220 28414 31272
rect 27430 31192 27436 31204
rect 25700 31164 27436 31192
rect 20395 31161 20407 31164
rect 20349 31155 20407 31161
rect 27430 31152 27436 31164
rect 27488 31152 27494 31204
rect 8478 31124 8484 31136
rect 5368 31096 8484 31124
rect 8478 31084 8484 31096
rect 8536 31084 8542 31136
rect 9674 31084 9680 31136
rect 9732 31124 9738 31136
rect 9953 31127 10011 31133
rect 9953 31124 9965 31127
rect 9732 31096 9965 31124
rect 9732 31084 9738 31096
rect 9953 31093 9965 31096
rect 9999 31093 10011 31127
rect 9953 31087 10011 31093
rect 10413 31127 10471 31133
rect 10413 31093 10425 31127
rect 10459 31124 10471 31127
rect 14182 31124 14188 31136
rect 10459 31096 14188 31124
rect 10459 31093 10471 31096
rect 10413 31087 10471 31093
rect 14182 31084 14188 31096
rect 14240 31084 14246 31136
rect 14918 31124 14924 31136
rect 14879 31096 14924 31124
rect 14918 31084 14924 31096
rect 14976 31084 14982 31136
rect 17310 31084 17316 31136
rect 17368 31124 17374 31136
rect 17681 31127 17739 31133
rect 17681 31124 17693 31127
rect 17368 31096 17693 31124
rect 17368 31084 17374 31096
rect 17681 31093 17693 31096
rect 17727 31093 17739 31127
rect 31726 31124 31754 31300
rect 32306 31220 32312 31272
rect 32364 31260 32370 31272
rect 32585 31263 32643 31269
rect 32585 31260 32597 31263
rect 32364 31232 32597 31260
rect 32364 31220 32370 31232
rect 32585 31229 32597 31232
rect 32631 31229 32643 31263
rect 32585 31223 32643 31229
rect 32674 31220 32680 31272
rect 32732 31260 32738 31272
rect 33888 31269 33916 31368
rect 34698 31356 34704 31368
rect 34756 31356 34762 31408
rect 34808 31396 34836 31436
rect 35253 31433 35265 31467
rect 35299 31464 35311 31467
rect 35342 31464 35348 31476
rect 35299 31436 35348 31464
rect 35299 31433 35311 31436
rect 35253 31427 35311 31433
rect 35342 31424 35348 31436
rect 35400 31424 35406 31476
rect 35710 31464 35716 31476
rect 35671 31436 35716 31464
rect 35710 31424 35716 31436
rect 35768 31424 35774 31476
rect 41049 31467 41107 31473
rect 35820 31436 40356 31464
rect 35820 31396 35848 31436
rect 40328 31405 40356 31436
rect 41049 31433 41061 31467
rect 41095 31464 41107 31467
rect 41230 31464 41236 31476
rect 41095 31436 41236 31464
rect 41095 31433 41107 31436
rect 41049 31427 41107 31433
rect 41230 31424 41236 31436
rect 41288 31424 41294 31476
rect 41509 31467 41567 31473
rect 41509 31433 41521 31467
rect 41555 31464 41567 31467
rect 41874 31464 41880 31476
rect 41555 31436 41880 31464
rect 41555 31433 41567 31436
rect 41509 31427 41567 31433
rect 41874 31424 41880 31436
rect 41932 31424 41938 31476
rect 37522 31399 37580 31405
rect 37522 31396 37534 31399
rect 34808 31368 35848 31396
rect 37384 31368 37534 31396
rect 33962 31288 33968 31340
rect 34020 31328 34026 31340
rect 34129 31331 34187 31337
rect 34129 31328 34141 31331
rect 34020 31300 34141 31328
rect 34020 31288 34026 31300
rect 34129 31297 34141 31300
rect 34175 31297 34187 31331
rect 35894 31328 35900 31340
rect 35855 31300 35900 31328
rect 34129 31291 34187 31297
rect 35894 31288 35900 31300
rect 35952 31288 35958 31340
rect 36541 31331 36599 31337
rect 36541 31297 36553 31331
rect 36587 31328 36599 31331
rect 36998 31328 37004 31340
rect 36587 31300 37004 31328
rect 36587 31297 36599 31300
rect 36541 31291 36599 31297
rect 36998 31288 37004 31300
rect 37056 31288 37062 31340
rect 37277 31331 37335 31337
rect 37277 31328 37289 31331
rect 37108 31300 37289 31328
rect 33873 31263 33931 31269
rect 32732 31232 32777 31260
rect 32732 31220 32738 31232
rect 33873 31229 33885 31263
rect 33919 31229 33931 31263
rect 33873 31223 33931 31229
rect 31938 31152 31944 31204
rect 31996 31192 32002 31204
rect 33888 31192 33916 31223
rect 35986 31220 35992 31272
rect 36044 31260 36050 31272
rect 37108 31260 37136 31300
rect 37277 31297 37289 31300
rect 37323 31297 37335 31331
rect 37277 31291 37335 31297
rect 37384 31260 37412 31368
rect 37522 31365 37534 31368
rect 37568 31365 37580 31399
rect 37522 31359 37580 31365
rect 40313 31399 40371 31405
rect 40313 31365 40325 31399
rect 40359 31396 40371 31399
rect 41141 31399 41199 31405
rect 41141 31396 41153 31399
rect 40359 31368 41153 31396
rect 40359 31365 40371 31368
rect 40313 31359 40371 31365
rect 41141 31365 41153 31368
rect 41187 31365 41199 31399
rect 41141 31359 41199 31365
rect 42426 31328 42432 31340
rect 42387 31300 42432 31328
rect 42426 31288 42432 31300
rect 42484 31288 42490 31340
rect 36044 31232 37136 31260
rect 37292 31232 37412 31260
rect 40957 31263 41015 31269
rect 36044 31220 36050 31232
rect 31996 31164 33916 31192
rect 36725 31195 36783 31201
rect 31996 31152 32002 31164
rect 36725 31161 36737 31195
rect 36771 31192 36783 31195
rect 37292 31192 37320 31232
rect 40957 31229 40969 31263
rect 41003 31229 41015 31263
rect 40957 31223 41015 31229
rect 36771 31164 37320 31192
rect 40972 31192 41000 31223
rect 41506 31192 41512 31204
rect 40972 31164 41512 31192
rect 36771 31161 36783 31164
rect 36725 31155 36783 31161
rect 41506 31152 41512 31164
rect 41564 31152 41570 31204
rect 32125 31127 32183 31133
rect 32125 31124 32137 31127
rect 31726 31096 32137 31124
rect 17681 31087 17739 31093
rect 32125 31093 32137 31096
rect 32171 31093 32183 31127
rect 32125 31087 32183 31093
rect 37458 31084 37464 31136
rect 37516 31124 37522 31136
rect 38562 31124 38568 31136
rect 37516 31096 38568 31124
rect 37516 31084 37522 31096
rect 38562 31084 38568 31096
rect 38620 31124 38626 31136
rect 38657 31127 38715 31133
rect 38657 31124 38669 31127
rect 38620 31096 38669 31124
rect 38620 31084 38626 31096
rect 38657 31093 38669 31096
rect 38703 31093 38715 31127
rect 38657 31087 38715 31093
rect 42613 31127 42671 31133
rect 42613 31093 42625 31127
rect 42659 31124 42671 31127
rect 43530 31124 43536 31136
rect 42659 31096 43536 31124
rect 42659 31093 42671 31096
rect 42613 31087 42671 31093
rect 43530 31084 43536 31096
rect 43588 31084 43594 31136
rect 1104 31034 68816 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 65654 31034
rect 65706 30982 65718 31034
rect 65770 30982 65782 31034
rect 65834 30982 65846 31034
rect 65898 30982 65910 31034
rect 65962 30982 68816 31034
rect 1104 30960 68816 30982
rect 5353 30923 5411 30929
rect 5353 30889 5365 30923
rect 5399 30920 5411 30923
rect 5534 30920 5540 30932
rect 5399 30892 5540 30920
rect 5399 30889 5411 30892
rect 5353 30883 5411 30889
rect 5534 30880 5540 30892
rect 5592 30880 5598 30932
rect 7193 30923 7251 30929
rect 7193 30889 7205 30923
rect 7239 30920 7251 30923
rect 7466 30920 7472 30932
rect 7239 30892 7472 30920
rect 7239 30889 7251 30892
rect 7193 30883 7251 30889
rect 7466 30880 7472 30892
rect 7524 30880 7530 30932
rect 8386 30920 8392 30932
rect 8347 30892 8392 30920
rect 8386 30880 8392 30892
rect 8444 30880 8450 30932
rect 8478 30880 8484 30932
rect 8536 30920 8542 30932
rect 15930 30920 15936 30932
rect 8536 30892 15936 30920
rect 8536 30880 8542 30892
rect 15930 30880 15936 30892
rect 15988 30880 15994 30932
rect 16574 30920 16580 30932
rect 16535 30892 16580 30920
rect 16574 30880 16580 30892
rect 16632 30880 16638 30932
rect 17497 30923 17555 30929
rect 17497 30889 17509 30923
rect 17543 30920 17555 30923
rect 18414 30920 18420 30932
rect 17543 30892 18420 30920
rect 17543 30889 17555 30892
rect 17497 30883 17555 30889
rect 18414 30880 18420 30892
rect 18472 30880 18478 30932
rect 18690 30920 18696 30932
rect 18651 30892 18696 30920
rect 18690 30880 18696 30892
rect 18748 30880 18754 30932
rect 19797 30923 19855 30929
rect 19797 30889 19809 30923
rect 19843 30920 19855 30923
rect 19843 30892 22094 30920
rect 19843 30889 19855 30892
rect 19797 30883 19855 30889
rect 16592 30852 16620 30880
rect 17954 30852 17960 30864
rect 16592 30824 17960 30852
rect 17954 30812 17960 30824
rect 18012 30812 18018 30864
rect 5074 30744 5080 30796
rect 5132 30784 5138 30796
rect 5442 30784 5448 30796
rect 5132 30756 5448 30784
rect 5132 30744 5138 30756
rect 5442 30744 5448 30756
rect 5500 30784 5506 30796
rect 5813 30787 5871 30793
rect 5813 30784 5825 30787
rect 5500 30756 5825 30784
rect 5500 30744 5506 30756
rect 5813 30753 5825 30756
rect 5859 30753 5871 30787
rect 5813 30747 5871 30753
rect 7098 30744 7104 30796
rect 7156 30784 7162 30796
rect 7745 30787 7803 30793
rect 7745 30784 7757 30787
rect 7156 30756 7757 30784
rect 7156 30744 7162 30756
rect 7745 30753 7757 30756
rect 7791 30753 7803 30787
rect 7745 30747 7803 30753
rect 12406 30756 17080 30784
rect 5166 30716 5172 30728
rect 5127 30688 5172 30716
rect 5166 30676 5172 30688
rect 5224 30676 5230 30728
rect 6080 30719 6138 30725
rect 6080 30685 6092 30719
rect 6126 30716 6138 30719
rect 6362 30716 6368 30728
rect 6126 30688 6368 30716
rect 6126 30685 6138 30688
rect 6080 30679 6138 30685
rect 6362 30676 6368 30688
rect 6420 30676 6426 30728
rect 8021 30719 8079 30725
rect 8021 30685 8033 30719
rect 8067 30716 8079 30719
rect 8294 30716 8300 30728
rect 8067 30688 8300 30716
rect 8067 30685 8079 30688
rect 8021 30679 8079 30685
rect 8294 30676 8300 30688
rect 8352 30676 8358 30728
rect 9033 30719 9091 30725
rect 9033 30685 9045 30719
rect 9079 30716 9091 30719
rect 9079 30688 12020 30716
rect 9079 30685 9091 30688
rect 9033 30679 9091 30685
rect 7926 30648 7932 30660
rect 7839 30620 7932 30648
rect 7926 30608 7932 30620
rect 7984 30648 7990 30660
rect 9048 30648 9076 30679
rect 7984 30620 9076 30648
rect 7984 30608 7990 30620
rect 11698 30608 11704 30660
rect 11756 30648 11762 30660
rect 11894 30651 11952 30657
rect 11894 30648 11906 30651
rect 11756 30620 11906 30648
rect 11756 30608 11762 30620
rect 11894 30617 11906 30620
rect 11940 30617 11952 30651
rect 11992 30648 12020 30688
rect 12066 30676 12072 30728
rect 12124 30716 12130 30728
rect 12161 30719 12219 30725
rect 12161 30716 12173 30719
rect 12124 30688 12173 30716
rect 12124 30676 12130 30688
rect 12161 30685 12173 30688
rect 12207 30685 12219 30719
rect 12161 30679 12219 30685
rect 12406 30648 12434 30756
rect 15470 30716 15476 30728
rect 15431 30688 15476 30716
rect 15470 30676 15476 30688
rect 15528 30676 15534 30728
rect 11992 30620 12434 30648
rect 11894 30611 11952 30617
rect 13722 30608 13728 30660
rect 13780 30648 13786 30660
rect 14185 30651 14243 30657
rect 14185 30648 14197 30651
rect 13780 30620 14197 30648
rect 13780 30608 13786 30620
rect 14185 30617 14197 30620
rect 14231 30648 14243 30651
rect 15013 30651 15071 30657
rect 15013 30648 15025 30651
rect 14231 30620 15025 30648
rect 14231 30617 14243 30620
rect 14185 30611 14243 30617
rect 15013 30617 15025 30620
rect 15059 30648 15071 30651
rect 16485 30651 16543 30657
rect 16485 30648 16497 30651
rect 15059 30620 16497 30648
rect 15059 30617 15071 30620
rect 15013 30611 15071 30617
rect 16485 30617 16497 30620
rect 16531 30648 16543 30651
rect 16942 30648 16948 30660
rect 16531 30620 16948 30648
rect 16531 30617 16543 30620
rect 16485 30611 16543 30617
rect 16942 30608 16948 30620
rect 17000 30608 17006 30660
rect 17052 30648 17080 30756
rect 17126 30744 17132 30796
rect 17184 30784 17190 30796
rect 18141 30787 18199 30793
rect 18141 30784 18153 30787
rect 17184 30756 18153 30784
rect 17184 30744 17190 30756
rect 18141 30753 18153 30756
rect 18187 30784 18199 30787
rect 20254 30784 20260 30796
rect 18187 30756 20260 30784
rect 18187 30753 18199 30756
rect 18141 30747 18199 30753
rect 20254 30744 20260 30756
rect 20312 30744 20318 30796
rect 17310 30716 17316 30728
rect 17271 30688 17316 30716
rect 17310 30676 17316 30688
rect 17368 30676 17374 30728
rect 20622 30716 20628 30728
rect 20583 30688 20628 30716
rect 20622 30676 20628 30688
rect 20680 30676 20686 30728
rect 18046 30648 18052 30660
rect 17052 30620 18052 30648
rect 18046 30608 18052 30620
rect 18104 30608 18110 30660
rect 19426 30608 19432 30660
rect 19484 30648 19490 30660
rect 19705 30651 19763 30657
rect 19705 30648 19717 30651
rect 19484 30620 19717 30648
rect 19484 30608 19490 30620
rect 19705 30617 19717 30620
rect 19751 30617 19763 30651
rect 19705 30611 19763 30617
rect 20892 30651 20950 30657
rect 20892 30617 20904 30651
rect 20938 30648 20950 30651
rect 21082 30648 21088 30660
rect 20938 30620 21088 30648
rect 20938 30617 20950 30620
rect 20892 30611 20950 30617
rect 21082 30608 21088 30620
rect 21140 30608 21146 30660
rect 22066 30648 22094 30892
rect 22186 30880 22192 30932
rect 22244 30920 22250 30932
rect 22465 30923 22523 30929
rect 22465 30920 22477 30923
rect 22244 30892 22477 30920
rect 22244 30880 22250 30892
rect 22465 30889 22477 30892
rect 22511 30889 22523 30923
rect 31294 30920 31300 30932
rect 22465 30883 22523 30889
rect 30208 30892 31300 30920
rect 27065 30855 27123 30861
rect 27065 30821 27077 30855
rect 27111 30852 27123 30855
rect 27154 30852 27160 30864
rect 27111 30824 27160 30852
rect 27111 30821 27123 30824
rect 27065 30815 27123 30821
rect 24394 30744 24400 30796
rect 24452 30784 24458 30796
rect 25685 30787 25743 30793
rect 25685 30784 25697 30787
rect 24452 30756 25697 30784
rect 24452 30744 24458 30756
rect 25685 30753 25697 30756
rect 25731 30753 25743 30787
rect 27080 30784 27108 30815
rect 27154 30812 27160 30824
rect 27212 30812 27218 30864
rect 30208 30793 30236 30892
rect 31294 30880 31300 30892
rect 31352 30920 31358 30932
rect 32674 30920 32680 30932
rect 31352 30892 32680 30920
rect 31352 30880 31358 30892
rect 32674 30880 32680 30892
rect 32732 30880 32738 30932
rect 36446 30920 36452 30932
rect 36407 30892 36452 30920
rect 36446 30880 36452 30892
rect 36504 30880 36510 30932
rect 36998 30920 37004 30932
rect 36959 30892 37004 30920
rect 36998 30880 37004 30892
rect 37056 30880 37062 30932
rect 41230 30920 41236 30932
rect 41191 30892 41236 30920
rect 41230 30880 41236 30892
rect 41288 30880 41294 30932
rect 31481 30855 31539 30861
rect 31481 30821 31493 30855
rect 31527 30852 31539 30855
rect 31527 30824 31754 30852
rect 31527 30821 31539 30824
rect 31481 30815 31539 30821
rect 27985 30787 28043 30793
rect 27985 30784 27997 30787
rect 27080 30756 27997 30784
rect 25685 30747 25743 30753
rect 27985 30753 27997 30756
rect 28031 30753 28043 30787
rect 27985 30747 28043 30753
rect 28077 30787 28135 30793
rect 28077 30753 28089 30787
rect 28123 30753 28135 30787
rect 28077 30747 28135 30753
rect 30193 30787 30251 30793
rect 30193 30753 30205 30787
rect 30239 30753 30251 30787
rect 31726 30784 31754 30824
rect 37458 30784 37464 30796
rect 31726 30756 32076 30784
rect 37419 30756 37464 30784
rect 30193 30747 30251 30753
rect 24670 30716 24676 30728
rect 24631 30688 24676 30716
rect 24670 30676 24676 30688
rect 24728 30676 24734 30728
rect 25225 30719 25283 30725
rect 25225 30685 25237 30719
rect 25271 30716 25283 30719
rect 25498 30716 25504 30728
rect 25271 30688 25504 30716
rect 25271 30685 25283 30688
rect 25225 30679 25283 30685
rect 23109 30651 23167 30657
rect 23109 30648 23121 30651
rect 22066 30620 23121 30648
rect 23109 30617 23121 30620
rect 23155 30648 23167 30651
rect 25240 30648 25268 30679
rect 25498 30676 25504 30688
rect 25556 30716 25562 30728
rect 25556 30688 26280 30716
rect 25556 30676 25562 30688
rect 25958 30657 25964 30660
rect 23155 30620 25268 30648
rect 23155 30617 23167 30620
rect 23109 30611 23167 30617
rect 25952 30611 25964 30657
rect 26016 30648 26022 30660
rect 26252 30648 26280 30688
rect 27430 30676 27436 30728
rect 27488 30716 27494 30728
rect 28092 30716 28120 30747
rect 27488 30688 28120 30716
rect 28997 30719 29055 30725
rect 27488 30676 27494 30688
rect 28997 30685 29009 30719
rect 29043 30716 29055 30719
rect 31297 30719 31355 30725
rect 29043 30688 30144 30716
rect 29043 30685 29055 30688
rect 28997 30679 29055 30685
rect 29012 30648 29040 30679
rect 26016 30620 26052 30648
rect 26252 30620 29040 30648
rect 25958 30608 25964 30611
rect 26016 30608 26022 30620
rect 29638 30608 29644 30660
rect 29696 30648 29702 30660
rect 30009 30651 30067 30657
rect 30009 30648 30021 30651
rect 29696 30620 30021 30648
rect 29696 30608 29702 30620
rect 30009 30617 30021 30620
rect 30055 30617 30067 30651
rect 30009 30611 30067 30617
rect 10781 30583 10839 30589
rect 10781 30549 10793 30583
rect 10827 30580 10839 30583
rect 12158 30580 12164 30592
rect 10827 30552 12164 30580
rect 10827 30549 10839 30552
rect 10781 30543 10839 30549
rect 12158 30540 12164 30552
rect 12216 30540 12222 30592
rect 15562 30540 15568 30592
rect 15620 30580 15626 30592
rect 15657 30583 15715 30589
rect 15657 30580 15669 30583
rect 15620 30552 15669 30580
rect 15620 30540 15626 30552
rect 15657 30549 15669 30552
rect 15703 30549 15715 30583
rect 15657 30543 15715 30549
rect 18138 30540 18144 30592
rect 18196 30580 18202 30592
rect 18233 30583 18291 30589
rect 18233 30580 18245 30583
rect 18196 30552 18245 30580
rect 18196 30540 18202 30552
rect 18233 30549 18245 30552
rect 18279 30549 18291 30583
rect 18233 30543 18291 30549
rect 18325 30583 18383 30589
rect 18325 30549 18337 30583
rect 18371 30580 18383 30583
rect 19334 30580 19340 30592
rect 18371 30552 19340 30580
rect 18371 30549 18383 30552
rect 18325 30543 18383 30549
rect 19334 30540 19340 30552
rect 19392 30540 19398 30592
rect 21910 30540 21916 30592
rect 21968 30580 21974 30592
rect 22005 30583 22063 30589
rect 22005 30580 22017 30583
rect 21968 30552 22017 30580
rect 21968 30540 21974 30552
rect 22005 30549 22017 30552
rect 22051 30549 22063 30583
rect 24486 30580 24492 30592
rect 24447 30552 24492 30580
rect 22005 30543 22063 30549
rect 24486 30540 24492 30552
rect 24544 30540 24550 30592
rect 27522 30580 27528 30592
rect 27483 30552 27528 30580
rect 27522 30540 27528 30552
rect 27580 30540 27586 30592
rect 27890 30580 27896 30592
rect 27851 30552 27896 30580
rect 27890 30540 27896 30552
rect 27948 30540 27954 30592
rect 28994 30540 29000 30592
rect 29052 30580 29058 30592
rect 29549 30583 29607 30589
rect 29549 30580 29561 30583
rect 29052 30552 29561 30580
rect 29052 30540 29058 30552
rect 29549 30549 29561 30552
rect 29595 30549 29607 30583
rect 29549 30543 29607 30549
rect 29917 30583 29975 30589
rect 29917 30549 29929 30583
rect 29963 30580 29975 30583
rect 30116 30580 30144 30688
rect 31297 30685 31309 30719
rect 31343 30716 31355 30719
rect 31938 30716 31944 30728
rect 31343 30688 31754 30716
rect 31899 30688 31944 30716
rect 31343 30685 31355 30688
rect 31297 30679 31355 30685
rect 31726 30648 31754 30688
rect 31938 30676 31944 30688
rect 31996 30676 32002 30728
rect 32048 30716 32076 30756
rect 37458 30744 37464 30756
rect 37516 30744 37522 30796
rect 37553 30787 37611 30793
rect 37553 30753 37565 30787
rect 37599 30753 37611 30787
rect 37553 30747 37611 30753
rect 32197 30719 32255 30725
rect 32197 30716 32209 30719
rect 32048 30688 32209 30716
rect 32197 30685 32209 30688
rect 32243 30685 32255 30719
rect 32197 30679 32255 30685
rect 37274 30676 37280 30728
rect 37332 30716 37338 30728
rect 37568 30716 37596 30747
rect 37332 30688 37596 30716
rect 37332 30676 37338 30688
rect 42058 30676 42064 30728
rect 42116 30716 42122 30728
rect 42346 30719 42404 30725
rect 42346 30716 42358 30719
rect 42116 30688 42358 30716
rect 42116 30676 42122 30688
rect 42346 30685 42358 30688
rect 42392 30685 42404 30719
rect 42346 30679 42404 30685
rect 42613 30719 42671 30725
rect 42613 30685 42625 30719
rect 42659 30716 42671 30719
rect 43806 30716 43812 30728
rect 42659 30688 43812 30716
rect 42659 30685 42671 30688
rect 42613 30679 42671 30685
rect 43806 30676 43812 30688
rect 43864 30676 43870 30728
rect 32030 30648 32036 30660
rect 31726 30620 32036 30648
rect 32030 30608 32036 30620
rect 32088 30608 32094 30660
rect 35802 30648 35808 30660
rect 32508 30620 35808 30648
rect 32508 30580 32536 30620
rect 35802 30608 35808 30620
rect 35860 30648 35866 30660
rect 35897 30651 35955 30657
rect 35897 30648 35909 30651
rect 35860 30620 35909 30648
rect 35860 30608 35866 30620
rect 35897 30617 35909 30620
rect 35943 30648 35955 30651
rect 37369 30651 37427 30657
rect 37369 30648 37381 30651
rect 35943 30620 37381 30648
rect 35943 30617 35955 30620
rect 35897 30611 35955 30617
rect 37369 30617 37381 30620
rect 37415 30617 37427 30651
rect 37369 30611 37427 30617
rect 29963 30552 32536 30580
rect 29963 30549 29975 30552
rect 29917 30543 29975 30549
rect 32582 30540 32588 30592
rect 32640 30580 32646 30592
rect 33321 30583 33379 30589
rect 33321 30580 33333 30583
rect 32640 30552 33333 30580
rect 32640 30540 32646 30552
rect 33321 30549 33333 30552
rect 33367 30549 33379 30583
rect 33321 30543 33379 30549
rect 1104 30490 68816 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 68816 30490
rect 1104 30416 68816 30438
rect 9766 30336 9772 30388
rect 9824 30376 9830 30388
rect 10321 30379 10379 30385
rect 10321 30376 10333 30379
rect 9824 30348 10333 30376
rect 9824 30336 9830 30348
rect 10321 30345 10333 30348
rect 10367 30345 10379 30379
rect 11698 30376 11704 30388
rect 11659 30348 11704 30376
rect 10321 30339 10379 30345
rect 11698 30336 11704 30348
rect 11756 30336 11762 30388
rect 15381 30379 15439 30385
rect 15381 30345 15393 30379
rect 15427 30376 15439 30379
rect 15470 30376 15476 30388
rect 15427 30348 15476 30376
rect 15427 30345 15439 30348
rect 15381 30339 15439 30345
rect 15470 30336 15476 30348
rect 15528 30336 15534 30388
rect 18046 30376 18052 30388
rect 18007 30348 18052 30376
rect 18046 30336 18052 30348
rect 18104 30376 18110 30388
rect 21082 30376 21088 30388
rect 18104 30348 19288 30376
rect 21043 30348 21088 30376
rect 18104 30336 18110 30348
rect 17034 30268 17040 30320
rect 17092 30308 17098 30320
rect 17313 30311 17371 30317
rect 17313 30308 17325 30311
rect 17092 30280 17325 30308
rect 17092 30268 17098 30280
rect 17313 30277 17325 30280
rect 17359 30308 17371 30311
rect 17957 30311 18015 30317
rect 17957 30308 17969 30311
rect 17359 30280 17969 30308
rect 17359 30277 17371 30280
rect 17313 30271 17371 30277
rect 17957 30277 17969 30280
rect 18003 30308 18015 30311
rect 18138 30308 18144 30320
rect 18003 30280 18144 30308
rect 18003 30277 18015 30280
rect 17957 30271 18015 30277
rect 18138 30268 18144 30280
rect 18196 30308 18202 30320
rect 18601 30311 18659 30317
rect 18601 30308 18613 30311
rect 18196 30280 18613 30308
rect 18196 30268 18202 30280
rect 18601 30277 18613 30280
rect 18647 30308 18659 30311
rect 18966 30308 18972 30320
rect 18647 30280 18972 30308
rect 18647 30277 18659 30280
rect 18601 30271 18659 30277
rect 18966 30268 18972 30280
rect 19024 30268 19030 30320
rect 19260 30308 19288 30348
rect 21082 30336 21088 30348
rect 21140 30336 21146 30388
rect 25958 30376 25964 30388
rect 25919 30348 25964 30376
rect 25958 30336 25964 30348
rect 26016 30336 26022 30388
rect 32030 30336 32036 30388
rect 32088 30376 32094 30388
rect 32125 30379 32183 30385
rect 32125 30376 32137 30379
rect 32088 30348 32137 30376
rect 32088 30336 32094 30348
rect 32125 30345 32137 30348
rect 32171 30345 32183 30379
rect 32125 30339 32183 30345
rect 41877 30379 41935 30385
rect 41877 30345 41889 30379
rect 41923 30376 41935 30379
rect 42426 30376 42432 30388
rect 41923 30348 42432 30376
rect 41923 30345 41935 30348
rect 41877 30339 41935 30345
rect 42426 30336 42432 30348
rect 42484 30336 42490 30388
rect 20530 30308 20536 30320
rect 19260 30280 20536 30308
rect 20530 30268 20536 30280
rect 20588 30268 20594 30320
rect 24296 30311 24354 30317
rect 24296 30277 24308 30311
rect 24342 30308 24354 30311
rect 24486 30308 24492 30320
rect 24342 30280 24492 30308
rect 24342 30277 24354 30280
rect 24296 30271 24354 30277
rect 24486 30268 24492 30280
rect 24544 30268 24550 30320
rect 27890 30268 27896 30320
rect 27948 30308 27954 30320
rect 31481 30311 31539 30317
rect 31481 30308 31493 30311
rect 27948 30280 31493 30308
rect 27948 30268 27954 30280
rect 31481 30277 31493 30280
rect 31527 30308 31539 30311
rect 32582 30308 32588 30320
rect 31527 30280 31754 30308
rect 32543 30280 32588 30308
rect 31527 30277 31539 30280
rect 31481 30271 31539 30277
rect 10689 30243 10747 30249
rect 10689 30209 10701 30243
rect 10735 30240 10747 30243
rect 11146 30240 11152 30252
rect 10735 30212 11152 30240
rect 10735 30209 10747 30212
rect 10689 30203 10747 30209
rect 11146 30200 11152 30212
rect 11204 30200 11210 30252
rect 11517 30243 11575 30249
rect 11517 30209 11529 30243
rect 11563 30240 11575 30243
rect 11790 30240 11796 30252
rect 11563 30212 11796 30240
rect 11563 30209 11575 30212
rect 11517 30203 11575 30209
rect 11790 30200 11796 30212
rect 11848 30200 11854 30252
rect 15749 30243 15807 30249
rect 15749 30209 15761 30243
rect 15795 30240 15807 30243
rect 16666 30240 16672 30252
rect 15795 30212 16672 30240
rect 15795 30209 15807 30212
rect 15749 30203 15807 30209
rect 16666 30200 16672 30212
rect 16724 30200 16730 30252
rect 21269 30243 21327 30249
rect 21269 30209 21281 30243
rect 21315 30240 21327 30243
rect 22186 30240 22192 30252
rect 21315 30212 21864 30240
rect 22147 30212 22192 30240
rect 21315 30209 21327 30212
rect 21269 30203 21327 30209
rect 10781 30175 10839 30181
rect 10781 30141 10793 30175
rect 10827 30172 10839 30175
rect 11054 30172 11060 30184
rect 10827 30144 11060 30172
rect 10827 30141 10839 30144
rect 10781 30135 10839 30141
rect 11054 30132 11060 30144
rect 11112 30132 11118 30184
rect 14921 30175 14979 30181
rect 14921 30141 14933 30175
rect 14967 30172 14979 30175
rect 15838 30172 15844 30184
rect 14967 30144 15844 30172
rect 14967 30141 14979 30144
rect 14921 30135 14979 30141
rect 15838 30132 15844 30144
rect 15896 30132 15902 30184
rect 15933 30175 15991 30181
rect 15933 30141 15945 30175
rect 15979 30141 15991 30175
rect 15933 30135 15991 30141
rect 13814 30064 13820 30116
rect 13872 30104 13878 30116
rect 15948 30104 15976 30135
rect 19426 30104 19432 30116
rect 13872 30076 15976 30104
rect 16960 30076 19432 30104
rect 13872 30064 13878 30076
rect 16960 30048 16988 30076
rect 19426 30064 19432 30076
rect 19484 30064 19490 30116
rect 21836 30113 21864 30212
rect 22186 30200 22192 30212
rect 22244 30240 22250 30252
rect 26145 30243 26203 30249
rect 22244 30212 26096 30240
rect 22244 30200 22250 30212
rect 21910 30132 21916 30184
rect 21968 30172 21974 30184
rect 22281 30175 22339 30181
rect 22281 30172 22293 30175
rect 21968 30144 22293 30172
rect 21968 30132 21974 30144
rect 22281 30141 22293 30144
rect 22327 30141 22339 30175
rect 22281 30135 22339 30141
rect 22465 30175 22523 30181
rect 22465 30141 22477 30175
rect 22511 30172 22523 30175
rect 22738 30172 22744 30184
rect 22511 30144 22744 30172
rect 22511 30141 22523 30144
rect 22465 30135 22523 30141
rect 22738 30132 22744 30144
rect 22796 30132 22802 30184
rect 24029 30175 24087 30181
rect 24029 30141 24041 30175
rect 24075 30141 24087 30175
rect 26068 30172 26096 30212
rect 26145 30209 26157 30243
rect 26191 30240 26203 30243
rect 27522 30240 27528 30252
rect 26191 30212 27528 30240
rect 26191 30209 26203 30212
rect 26145 30203 26203 30209
rect 27522 30200 27528 30212
rect 27580 30200 27586 30252
rect 28261 30243 28319 30249
rect 28261 30209 28273 30243
rect 28307 30240 28319 30243
rect 28350 30240 28356 30252
rect 28307 30212 28356 30240
rect 28307 30209 28319 30212
rect 28261 30203 28319 30209
rect 28350 30200 28356 30212
rect 28408 30200 28414 30252
rect 28528 30243 28586 30249
rect 28528 30209 28540 30243
rect 28574 30240 28586 30243
rect 28810 30240 28816 30252
rect 28574 30212 28816 30240
rect 28574 30209 28586 30212
rect 28528 30203 28586 30209
rect 28810 30200 28816 30212
rect 28868 30200 28874 30252
rect 30834 30240 30840 30252
rect 30795 30212 30840 30240
rect 30834 30200 30840 30212
rect 30892 30200 30898 30252
rect 31726 30240 31754 30280
rect 32582 30268 32588 30280
rect 32640 30268 32646 30320
rect 43530 30268 43536 30320
rect 43588 30317 43594 30320
rect 43588 30308 43600 30317
rect 43588 30280 43633 30308
rect 43588 30271 43600 30280
rect 43588 30268 43594 30271
rect 32490 30240 32496 30252
rect 31726 30212 32496 30240
rect 32490 30200 32496 30212
rect 32548 30200 32554 30252
rect 36449 30243 36507 30249
rect 36449 30209 36461 30243
rect 36495 30240 36507 30243
rect 37274 30240 37280 30252
rect 36495 30212 37280 30240
rect 36495 30209 36507 30212
rect 36449 30203 36507 30209
rect 37274 30200 37280 30212
rect 37332 30200 37338 30252
rect 40402 30240 40408 30252
rect 40363 30212 40408 30240
rect 40402 30200 40408 30212
rect 40460 30200 40466 30252
rect 40678 30240 40684 30252
rect 40639 30212 40684 30240
rect 40678 30200 40684 30212
rect 40736 30200 40742 30252
rect 40770 30200 40776 30252
rect 40828 30240 40834 30252
rect 41509 30243 41567 30249
rect 41509 30240 41521 30243
rect 40828 30212 41521 30240
rect 40828 30200 40834 30212
rect 41509 30209 41521 30212
rect 41555 30209 41567 30243
rect 43806 30240 43812 30252
rect 43767 30212 43812 30240
rect 41509 30203 41567 30209
rect 43806 30200 43812 30212
rect 43864 30200 43870 30252
rect 27341 30175 27399 30181
rect 27341 30172 27353 30175
rect 26068 30144 27353 30172
rect 24029 30135 24087 30141
rect 27341 30141 27353 30144
rect 27387 30172 27399 30175
rect 27890 30172 27896 30184
rect 27387 30144 27896 30172
rect 27387 30141 27399 30144
rect 27341 30135 27399 30141
rect 21821 30107 21879 30113
rect 21821 30073 21833 30107
rect 21867 30073 21879 30107
rect 21821 30067 21879 30073
rect 16853 30039 16911 30045
rect 16853 30005 16865 30039
rect 16899 30036 16911 30039
rect 16942 30036 16948 30048
rect 16899 30008 16948 30036
rect 16899 30005 16911 30008
rect 16853 29999 16911 30005
rect 16942 29996 16948 30008
rect 17000 29996 17006 30048
rect 20070 30036 20076 30048
rect 20031 30008 20076 30036
rect 20070 29996 20076 30008
rect 20128 29996 20134 30048
rect 24044 30036 24072 30135
rect 27890 30132 27896 30144
rect 27948 30132 27954 30184
rect 32674 30172 32680 30184
rect 32635 30144 32680 30172
rect 32674 30132 32680 30144
rect 32732 30132 32738 30184
rect 40586 30172 40592 30184
rect 40547 30144 40592 30172
rect 40586 30132 40592 30144
rect 40644 30132 40650 30184
rect 41325 30175 41383 30181
rect 41325 30141 41337 30175
rect 41371 30141 41383 30175
rect 41325 30135 41383 30141
rect 41417 30175 41475 30181
rect 41417 30141 41429 30175
rect 41463 30141 41475 30175
rect 41417 30135 41475 30141
rect 24394 30036 24400 30048
rect 24044 30008 24400 30036
rect 24394 29996 24400 30008
rect 24452 29996 24458 30048
rect 24762 29996 24768 30048
rect 24820 30036 24826 30048
rect 25409 30039 25467 30045
rect 25409 30036 25421 30039
rect 24820 30008 25421 30036
rect 24820 29996 24826 30008
rect 25409 30005 25421 30008
rect 25455 30005 25467 30039
rect 29638 30036 29644 30048
rect 29599 30008 29644 30036
rect 25409 29999 25467 30005
rect 29638 29996 29644 30008
rect 29696 29996 29702 30048
rect 30650 30036 30656 30048
rect 30611 30008 30656 30036
rect 30650 29996 30656 30008
rect 30708 29996 30714 30048
rect 36265 30039 36323 30045
rect 36265 30005 36277 30039
rect 36311 30036 36323 30039
rect 36354 30036 36360 30048
rect 36311 30008 36360 30036
rect 36311 30005 36323 30008
rect 36265 29999 36323 30005
rect 36354 29996 36360 30008
rect 36412 29996 36418 30048
rect 40126 29996 40132 30048
rect 40184 30036 40190 30048
rect 40221 30039 40279 30045
rect 40221 30036 40233 30039
rect 40184 30008 40233 30036
rect 40184 29996 40190 30008
rect 40221 30005 40233 30008
rect 40267 30005 40279 30039
rect 40221 29999 40279 30005
rect 40681 30039 40739 30045
rect 40681 30005 40693 30039
rect 40727 30036 40739 30039
rect 40862 30036 40868 30048
rect 40727 30008 40868 30036
rect 40727 30005 40739 30008
rect 40681 29999 40739 30005
rect 40862 29996 40868 30008
rect 40920 29996 40926 30048
rect 41340 30036 41368 30135
rect 41432 30104 41460 30135
rect 41598 30104 41604 30116
rect 41432 30076 41604 30104
rect 41598 30064 41604 30076
rect 41656 30104 41662 30116
rect 42429 30107 42487 30113
rect 42429 30104 42441 30107
rect 41656 30076 42441 30104
rect 41656 30064 41662 30076
rect 42429 30073 42441 30076
rect 42475 30073 42487 30107
rect 42429 30067 42487 30073
rect 41506 30036 41512 30048
rect 41340 30008 41512 30036
rect 41506 29996 41512 30008
rect 41564 29996 41570 30048
rect 1104 29946 68816 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 65654 29946
rect 65706 29894 65718 29946
rect 65770 29894 65782 29946
rect 65834 29894 65846 29946
rect 65898 29894 65910 29946
rect 65962 29894 68816 29946
rect 1104 29872 68816 29894
rect 11790 29832 11796 29844
rect 11751 29804 11796 29832
rect 11790 29792 11796 29804
rect 11848 29792 11854 29844
rect 16666 29832 16672 29844
rect 16627 29804 16672 29832
rect 16666 29792 16672 29804
rect 16724 29792 16730 29844
rect 24670 29792 24676 29844
rect 24728 29832 24734 29844
rect 24765 29835 24823 29841
rect 24765 29832 24777 29835
rect 24728 29804 24777 29832
rect 24728 29792 24734 29804
rect 24765 29801 24777 29804
rect 24811 29801 24823 29835
rect 28810 29832 28816 29844
rect 28771 29804 28816 29832
rect 24765 29795 24823 29801
rect 28810 29792 28816 29804
rect 28868 29792 28874 29844
rect 32490 29792 32496 29844
rect 32548 29832 32554 29844
rect 37642 29832 37648 29844
rect 32548 29804 37648 29832
rect 32548 29792 32554 29804
rect 37642 29792 37648 29804
rect 37700 29832 37706 29844
rect 37829 29835 37887 29841
rect 37829 29832 37841 29835
rect 37700 29804 37841 29832
rect 37700 29792 37706 29804
rect 37829 29801 37841 29804
rect 37875 29801 37887 29835
rect 37829 29795 37887 29801
rect 6273 29767 6331 29773
rect 6273 29733 6285 29767
rect 6319 29733 6331 29767
rect 6273 29727 6331 29733
rect 7285 29767 7343 29773
rect 7285 29733 7297 29767
rect 7331 29764 7343 29767
rect 9493 29767 9551 29773
rect 7331 29736 9076 29764
rect 7331 29733 7343 29736
rect 7285 29727 7343 29733
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29628 4951 29631
rect 4982 29628 4988 29640
rect 4939 29600 4988 29628
rect 4939 29597 4951 29600
rect 4893 29591 4951 29597
rect 4982 29588 4988 29600
rect 5040 29588 5046 29640
rect 6288 29628 6316 29727
rect 7006 29696 7012 29708
rect 6967 29668 7012 29696
rect 7006 29656 7012 29668
rect 7064 29656 7070 29708
rect 9048 29705 9076 29736
rect 9493 29733 9505 29767
rect 9539 29764 9551 29767
rect 9950 29764 9956 29776
rect 9539 29736 9956 29764
rect 9539 29733 9551 29736
rect 9493 29727 9551 29733
rect 9950 29724 9956 29736
rect 10008 29724 10014 29776
rect 37844 29764 37872 29795
rect 40586 29792 40592 29844
rect 40644 29832 40650 29844
rect 41325 29835 41383 29841
rect 41325 29832 41337 29835
rect 40644 29804 41337 29832
rect 40644 29792 40650 29804
rect 41325 29801 41337 29804
rect 41371 29801 41383 29835
rect 67358 29832 67364 29844
rect 67319 29804 67364 29832
rect 41325 29795 41383 29801
rect 67358 29792 67364 29804
rect 67416 29792 67422 29844
rect 40681 29767 40739 29773
rect 40681 29764 40693 29767
rect 37844 29736 40693 29764
rect 40681 29733 40693 29736
rect 40727 29764 40739 29767
rect 40770 29764 40776 29776
rect 40727 29736 40776 29764
rect 40727 29733 40739 29736
rect 40681 29727 40739 29733
rect 40770 29724 40776 29736
rect 40828 29724 40834 29776
rect 9033 29699 9091 29705
rect 9033 29665 9045 29699
rect 9079 29665 9091 29699
rect 9033 29659 9091 29665
rect 12345 29699 12403 29705
rect 12345 29665 12357 29699
rect 12391 29696 12403 29699
rect 13814 29696 13820 29708
rect 12391 29668 13820 29696
rect 12391 29665 12403 29668
rect 12345 29659 12403 29665
rect 13814 29656 13820 29668
rect 13872 29656 13878 29708
rect 25409 29699 25467 29705
rect 25409 29665 25421 29699
rect 25455 29696 25467 29699
rect 27522 29696 27528 29708
rect 25455 29668 27528 29696
rect 25455 29665 25467 29668
rect 25409 29659 25467 29665
rect 27522 29656 27528 29668
rect 27580 29656 27586 29708
rect 28350 29656 28356 29708
rect 28408 29696 28414 29708
rect 30466 29696 30472 29708
rect 28408 29668 30472 29696
rect 28408 29656 28414 29668
rect 30466 29656 30472 29668
rect 30524 29656 30530 29708
rect 35986 29696 35992 29708
rect 35947 29668 35992 29696
rect 35986 29656 35992 29668
rect 36044 29656 36050 29708
rect 41046 29656 41052 29708
rect 41104 29696 41110 29708
rect 41509 29699 41567 29705
rect 41509 29696 41521 29699
rect 41104 29668 41521 29696
rect 41104 29656 41110 29668
rect 41509 29665 41521 29668
rect 41555 29665 41567 29699
rect 41509 29659 41567 29665
rect 6730 29628 6736 29640
rect 6288 29600 6736 29628
rect 6730 29588 6736 29600
rect 6788 29628 6794 29640
rect 6917 29631 6975 29637
rect 6917 29628 6929 29631
rect 6788 29600 6929 29628
rect 6788 29588 6794 29600
rect 6917 29597 6929 29600
rect 6963 29597 6975 29631
rect 9122 29628 9128 29640
rect 9083 29600 9128 29628
rect 6917 29591 6975 29597
rect 9122 29588 9128 29600
rect 9180 29588 9186 29640
rect 10962 29628 10968 29640
rect 10923 29600 10968 29628
rect 10962 29588 10968 29600
rect 11020 29588 11026 29640
rect 11146 29628 11152 29640
rect 11107 29600 11152 29628
rect 11146 29588 11152 29600
rect 11204 29628 11210 29640
rect 11790 29628 11796 29640
rect 11204 29600 11796 29628
rect 11204 29588 11210 29600
rect 11790 29588 11796 29600
rect 11848 29628 11854 29640
rect 15289 29631 15347 29637
rect 11848 29600 12434 29628
rect 11848 29588 11854 29600
rect 5160 29563 5218 29569
rect 5160 29529 5172 29563
rect 5206 29560 5218 29563
rect 5258 29560 5264 29572
rect 5206 29532 5264 29560
rect 5206 29529 5218 29532
rect 5160 29523 5218 29529
rect 5258 29520 5264 29532
rect 5316 29520 5322 29572
rect 12158 29560 12164 29572
rect 12119 29532 12164 29560
rect 12158 29520 12164 29532
rect 12216 29520 12222 29572
rect 12406 29560 12434 29600
rect 15289 29597 15301 29631
rect 15335 29628 15347 29631
rect 15378 29628 15384 29640
rect 15335 29600 15384 29628
rect 15335 29597 15347 29600
rect 15289 29591 15347 29597
rect 15378 29588 15384 29600
rect 15436 29588 15442 29640
rect 15562 29637 15568 29640
rect 15556 29628 15568 29637
rect 15523 29600 15568 29628
rect 15556 29591 15568 29600
rect 15562 29588 15568 29591
rect 15620 29588 15626 29640
rect 16666 29588 16672 29640
rect 16724 29628 16730 29640
rect 17497 29631 17555 29637
rect 17497 29628 17509 29631
rect 16724 29600 17509 29628
rect 16724 29588 16730 29600
rect 17497 29597 17509 29600
rect 17543 29597 17555 29631
rect 17497 29591 17555 29597
rect 17957 29631 18015 29637
rect 17957 29597 17969 29631
rect 18003 29628 18015 29631
rect 18322 29628 18328 29640
rect 18003 29600 18328 29628
rect 18003 29597 18015 29600
rect 17957 29591 18015 29597
rect 18322 29588 18328 29600
rect 18380 29588 18386 29640
rect 19242 29588 19248 29640
rect 19300 29628 19306 29640
rect 19429 29631 19487 29637
rect 19429 29628 19441 29631
rect 19300 29600 19441 29628
rect 19300 29588 19306 29600
rect 19429 29597 19441 29600
rect 19475 29597 19487 29631
rect 19429 29591 19487 29597
rect 20441 29631 20499 29637
rect 20441 29597 20453 29631
rect 20487 29628 20499 29631
rect 21637 29631 21695 29637
rect 21637 29628 21649 29631
rect 20487 29600 21649 29628
rect 20487 29597 20499 29600
rect 20441 29591 20499 29597
rect 21637 29597 21649 29600
rect 21683 29628 21695 29631
rect 22186 29628 22192 29640
rect 21683 29600 22192 29628
rect 21683 29597 21695 29600
rect 21637 29591 21695 29597
rect 22186 29588 22192 29600
rect 22244 29588 22250 29640
rect 28994 29628 29000 29640
rect 28955 29600 29000 29628
rect 28994 29588 29000 29600
rect 29052 29588 29058 29640
rect 30736 29631 30794 29637
rect 30736 29597 30748 29631
rect 30782 29597 30794 29631
rect 30736 29591 30794 29597
rect 35345 29631 35403 29637
rect 35345 29597 35357 29631
rect 35391 29628 35403 29631
rect 35894 29628 35900 29640
rect 35391 29600 35900 29628
rect 35391 29597 35403 29600
rect 35345 29591 35403 29597
rect 17129 29563 17187 29569
rect 17129 29560 17141 29563
rect 12406 29532 17141 29560
rect 17129 29529 17141 29532
rect 17175 29529 17187 29563
rect 17129 29523 17187 29529
rect 20070 29520 20076 29572
rect 20128 29560 20134 29572
rect 20257 29563 20315 29569
rect 20257 29560 20269 29563
rect 20128 29532 20269 29560
rect 20128 29520 20134 29532
rect 20257 29529 20269 29532
rect 20303 29529 20315 29563
rect 20257 29523 20315 29529
rect 24762 29520 24768 29572
rect 24820 29560 24826 29572
rect 25225 29563 25283 29569
rect 25225 29560 25237 29563
rect 24820 29532 25237 29560
rect 24820 29520 24826 29532
rect 25225 29529 25237 29532
rect 25271 29529 25283 29563
rect 25225 29523 25283 29529
rect 30650 29520 30656 29572
rect 30708 29560 30714 29572
rect 30760 29560 30788 29591
rect 35894 29588 35900 29600
rect 35952 29588 35958 29640
rect 41598 29628 41604 29640
rect 41559 29600 41604 29628
rect 41598 29588 41604 29600
rect 41656 29588 41662 29640
rect 61378 29588 61384 29640
rect 61436 29628 61442 29640
rect 67177 29631 67235 29637
rect 67177 29628 67189 29631
rect 61436 29600 67189 29628
rect 61436 29588 61442 29600
rect 67177 29597 67189 29600
rect 67223 29628 67235 29631
rect 67821 29631 67879 29637
rect 67821 29628 67833 29631
rect 67223 29600 67833 29628
rect 67223 29597 67235 29600
rect 67177 29591 67235 29597
rect 67821 29597 67833 29600
rect 67867 29597 67879 29631
rect 67821 29591 67879 29597
rect 36234 29563 36292 29569
rect 36234 29560 36246 29563
rect 30708 29532 30788 29560
rect 35544 29532 36246 29560
rect 30708 29520 30714 29532
rect 11333 29495 11391 29501
rect 11333 29461 11345 29495
rect 11379 29492 11391 29495
rect 11698 29492 11704 29504
rect 11379 29464 11704 29492
rect 11379 29461 11391 29464
rect 11333 29455 11391 29461
rect 11698 29452 11704 29464
rect 11756 29452 11762 29504
rect 12253 29495 12311 29501
rect 12253 29461 12265 29495
rect 12299 29492 12311 29495
rect 13081 29495 13139 29501
rect 13081 29492 13093 29495
rect 12299 29464 13093 29492
rect 12299 29461 12311 29464
rect 12253 29455 12311 29461
rect 13081 29461 13093 29464
rect 13127 29492 13139 29495
rect 13906 29492 13912 29504
rect 13127 29464 13912 29492
rect 13127 29461 13139 29464
rect 13081 29455 13139 29461
rect 13906 29452 13912 29464
rect 13964 29452 13970 29504
rect 14737 29495 14795 29501
rect 14737 29461 14749 29495
rect 14783 29492 14795 29495
rect 15102 29492 15108 29504
rect 14783 29464 15108 29492
rect 14783 29461 14795 29464
rect 14737 29455 14795 29461
rect 15102 29452 15108 29464
rect 15160 29452 15166 29504
rect 19245 29495 19303 29501
rect 19245 29461 19257 29495
rect 19291 29492 19303 29495
rect 19426 29492 19432 29504
rect 19291 29464 19432 29492
rect 19291 29461 19303 29464
rect 19245 29455 19303 29461
rect 19426 29452 19432 29464
rect 19484 29452 19490 29504
rect 23842 29492 23848 29504
rect 23755 29464 23848 29492
rect 23842 29452 23848 29464
rect 23900 29492 23906 29504
rect 25133 29495 25191 29501
rect 25133 29492 25145 29495
rect 23900 29464 25145 29492
rect 23900 29452 23906 29464
rect 25133 29461 25145 29464
rect 25179 29492 25191 29495
rect 25406 29492 25412 29504
rect 25179 29464 25412 29492
rect 25179 29461 25191 29464
rect 25133 29455 25191 29461
rect 25406 29452 25412 29464
rect 25464 29452 25470 29504
rect 31386 29452 31392 29504
rect 31444 29492 31450 29504
rect 35544 29501 35572 29532
rect 36234 29529 36246 29532
rect 36280 29529 36292 29563
rect 36234 29523 36292 29529
rect 31849 29495 31907 29501
rect 31849 29492 31861 29495
rect 31444 29464 31861 29492
rect 31444 29452 31450 29464
rect 31849 29461 31861 29464
rect 31895 29461 31907 29495
rect 31849 29455 31907 29461
rect 35529 29495 35587 29501
rect 35529 29461 35541 29495
rect 35575 29461 35587 29495
rect 37366 29492 37372 29504
rect 37327 29464 37372 29492
rect 35529 29455 35587 29461
rect 37366 29452 37372 29464
rect 37424 29452 37430 29504
rect 38654 29452 38660 29504
rect 38712 29492 38718 29504
rect 40954 29492 40960 29504
rect 38712 29464 40960 29492
rect 38712 29452 38718 29464
rect 40954 29452 40960 29464
rect 41012 29452 41018 29504
rect 42794 29452 42800 29504
rect 42852 29492 42858 29504
rect 43073 29495 43131 29501
rect 43073 29492 43085 29495
rect 42852 29464 43085 29492
rect 42852 29452 42858 29464
rect 43073 29461 43085 29464
rect 43119 29461 43131 29495
rect 43073 29455 43131 29461
rect 1104 29402 68816 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 68816 29402
rect 1104 29328 68816 29350
rect 5258 29288 5264 29300
rect 5219 29260 5264 29288
rect 5258 29248 5264 29260
rect 5316 29248 5322 29300
rect 6730 29288 6736 29300
rect 6691 29260 6736 29288
rect 6730 29248 6736 29260
rect 6788 29248 6794 29300
rect 12897 29291 12955 29297
rect 12897 29257 12909 29291
rect 12943 29288 12955 29291
rect 13998 29288 14004 29300
rect 12943 29260 14004 29288
rect 12943 29257 12955 29260
rect 12897 29251 12955 29257
rect 13998 29248 14004 29260
rect 14056 29248 14062 29300
rect 14550 29248 14556 29300
rect 14608 29288 14614 29300
rect 37274 29288 37280 29300
rect 14608 29260 36584 29288
rect 37235 29260 37280 29288
rect 14608 29248 14614 29260
rect 6178 29180 6184 29232
rect 6236 29220 6242 29232
rect 6825 29223 6883 29229
rect 6825 29220 6837 29223
rect 6236 29192 6837 29220
rect 6236 29180 6242 29192
rect 6825 29189 6837 29192
rect 6871 29220 6883 29223
rect 7561 29223 7619 29229
rect 7561 29220 7573 29223
rect 6871 29192 7573 29220
rect 6871 29189 6883 29192
rect 6825 29183 6883 29189
rect 7561 29189 7573 29192
rect 7607 29189 7619 29223
rect 7561 29183 7619 29189
rect 9309 29223 9367 29229
rect 9309 29189 9321 29223
rect 9355 29220 9367 29223
rect 10413 29223 10471 29229
rect 10413 29220 10425 29223
rect 9355 29192 10425 29220
rect 9355 29189 9367 29192
rect 9309 29183 9367 29189
rect 10413 29189 10425 29192
rect 10459 29220 10471 29223
rect 15930 29220 15936 29232
rect 10459 29192 11560 29220
rect 15891 29192 15936 29220
rect 10459 29189 10471 29192
rect 10413 29183 10471 29189
rect 5445 29155 5503 29161
rect 5445 29121 5457 29155
rect 5491 29152 5503 29155
rect 5491 29124 6408 29152
rect 5491 29121 5503 29124
rect 5445 29115 5503 29121
rect 6380 29025 6408 29124
rect 7006 29112 7012 29164
rect 7064 29152 7070 29164
rect 9125 29155 9183 29161
rect 9125 29152 9137 29155
rect 7064 29124 9137 29152
rect 7064 29112 7070 29124
rect 9125 29121 9137 29124
rect 9171 29121 9183 29155
rect 10318 29152 10324 29164
rect 10279 29124 10324 29152
rect 9125 29115 9183 29121
rect 10318 29112 10324 29124
rect 10376 29112 10382 29164
rect 10597 29155 10655 29161
rect 10597 29121 10609 29155
rect 10643 29152 10655 29155
rect 11146 29152 11152 29164
rect 10643 29124 11152 29152
rect 10643 29121 10655 29124
rect 10597 29115 10655 29121
rect 11146 29112 11152 29124
rect 11204 29112 11210 29164
rect 11532 29161 11560 29192
rect 15930 29180 15936 29192
rect 15988 29180 15994 29232
rect 16500 29192 17724 29220
rect 11517 29155 11575 29161
rect 11517 29121 11529 29155
rect 11563 29121 11575 29155
rect 11698 29152 11704 29164
rect 11659 29124 11704 29152
rect 11517 29115 11575 29121
rect 11698 29112 11704 29124
rect 11756 29112 11762 29164
rect 12526 29152 12532 29164
rect 12487 29124 12532 29152
rect 12526 29112 12532 29124
rect 12584 29112 12590 29164
rect 14369 29155 14427 29161
rect 14369 29121 14381 29155
rect 14415 29152 14427 29155
rect 15102 29152 15108 29164
rect 14415 29124 15108 29152
rect 14415 29121 14427 29124
rect 14369 29115 14427 29121
rect 15102 29112 15108 29124
rect 15160 29112 15166 29164
rect 15197 29155 15255 29161
rect 15197 29121 15209 29155
rect 15243 29152 15255 29155
rect 15749 29155 15807 29161
rect 15749 29152 15761 29155
rect 15243 29124 15761 29152
rect 15243 29121 15255 29124
rect 15197 29115 15255 29121
rect 15749 29121 15761 29124
rect 15795 29152 15807 29155
rect 15838 29152 15844 29164
rect 15795 29124 15844 29152
rect 15795 29121 15807 29124
rect 15749 29115 15807 29121
rect 15838 29112 15844 29124
rect 15896 29152 15902 29164
rect 16500 29152 16528 29192
rect 16666 29152 16672 29164
rect 15896 29124 16528 29152
rect 16627 29124 16672 29152
rect 15896 29112 15902 29124
rect 16666 29112 16672 29124
rect 16724 29112 16730 29164
rect 16850 29112 16856 29164
rect 16908 29152 16914 29164
rect 17696 29152 17724 29192
rect 18230 29180 18236 29232
rect 18288 29220 18294 29232
rect 18288 29192 19748 29220
rect 18288 29180 18294 29192
rect 19058 29152 19064 29164
rect 16908 29124 17448 29152
rect 17696 29124 19064 29152
rect 16908 29112 16914 29124
rect 6917 29087 6975 29093
rect 6917 29053 6929 29087
rect 6963 29084 6975 29087
rect 7098 29084 7104 29096
rect 6963 29056 7104 29084
rect 6963 29053 6975 29056
rect 6917 29047 6975 29053
rect 7098 29044 7104 29056
rect 7156 29044 7162 29096
rect 8941 29087 8999 29093
rect 8941 29053 8953 29087
rect 8987 29084 8999 29087
rect 9582 29084 9588 29096
rect 8987 29056 9588 29084
rect 8987 29053 8999 29056
rect 8941 29047 8999 29053
rect 9582 29044 9588 29056
rect 9640 29044 9646 29096
rect 12621 29087 12679 29093
rect 12621 29053 12633 29087
rect 12667 29053 12679 29087
rect 14274 29084 14280 29096
rect 14235 29056 14280 29084
rect 12621 29047 12679 29053
rect 6365 29019 6423 29025
rect 6365 28985 6377 29019
rect 6411 28985 6423 29019
rect 6365 28979 6423 28985
rect 10781 29019 10839 29025
rect 10781 28985 10793 29019
rect 10827 29016 10839 29019
rect 11054 29016 11060 29028
rect 10827 28988 11060 29016
rect 10827 28985 10839 28988
rect 10781 28979 10839 28985
rect 11054 28976 11060 28988
rect 11112 28976 11118 29028
rect 11885 29019 11943 29025
rect 11885 28985 11897 29019
rect 11931 29016 11943 29019
rect 12434 29016 12440 29028
rect 11931 28988 12440 29016
rect 11931 28985 11943 28988
rect 11885 28979 11943 28985
rect 12434 28976 12440 28988
rect 12492 28976 12498 29028
rect 12636 29016 12664 29047
rect 14274 29044 14280 29056
rect 14332 29044 14338 29096
rect 17420 29025 17448 29124
rect 19058 29112 19064 29124
rect 19116 29112 19122 29164
rect 19426 29112 19432 29164
rect 19484 29161 19490 29164
rect 19720 29161 19748 29192
rect 30466 29180 30472 29232
rect 30524 29220 30530 29232
rect 31938 29220 31944 29232
rect 30524 29192 31944 29220
rect 30524 29180 30530 29192
rect 19484 29152 19496 29161
rect 19705 29155 19763 29161
rect 19484 29124 19529 29152
rect 19484 29115 19496 29124
rect 19705 29121 19717 29155
rect 19751 29152 19763 29155
rect 20714 29152 20720 29164
rect 19751 29124 20720 29152
rect 19751 29121 19763 29124
rect 19705 29115 19763 29121
rect 19484 29112 19490 29115
rect 20714 29112 20720 29124
rect 20772 29152 20778 29164
rect 21726 29152 21732 29164
rect 20772 29124 21732 29152
rect 20772 29112 20778 29124
rect 21726 29112 21732 29124
rect 21784 29112 21790 29164
rect 22094 29112 22100 29164
rect 22152 29152 22158 29164
rect 24578 29152 24584 29164
rect 22152 29124 22197 29152
rect 24539 29124 24584 29152
rect 22152 29112 22158 29124
rect 24578 29112 24584 29124
rect 24636 29112 24642 29164
rect 31588 29161 31616 29192
rect 31938 29180 31944 29192
rect 31996 29220 32002 29232
rect 35152 29223 35210 29229
rect 31996 29192 34744 29220
rect 31996 29180 32002 29192
rect 31317 29155 31375 29161
rect 31317 29121 31329 29155
rect 31363 29152 31375 29155
rect 31573 29155 31631 29161
rect 31363 29124 31524 29152
rect 31363 29121 31375 29124
rect 31317 29115 31375 29121
rect 31496 29084 31524 29124
rect 31573 29121 31585 29155
rect 31619 29152 31631 29155
rect 32309 29155 32367 29161
rect 32309 29152 32321 29155
rect 31619 29124 31653 29152
rect 31726 29124 32321 29152
rect 31619 29121 31631 29124
rect 31573 29115 31631 29121
rect 31726 29096 31754 29124
rect 32309 29121 32321 29124
rect 32355 29121 32367 29155
rect 32309 29115 32367 29121
rect 34716 29096 34744 29192
rect 35152 29189 35164 29223
rect 35198 29220 35210 29223
rect 35342 29220 35348 29232
rect 35198 29192 35348 29220
rect 35198 29189 35210 29192
rect 35152 29183 35210 29189
rect 35342 29180 35348 29192
rect 35400 29180 35406 29232
rect 36556 29220 36584 29260
rect 37274 29248 37280 29260
rect 37332 29248 37338 29300
rect 37642 29288 37648 29300
rect 37603 29260 37648 29288
rect 37642 29248 37648 29260
rect 37700 29248 37706 29300
rect 40037 29291 40095 29297
rect 40037 29257 40049 29291
rect 40083 29288 40095 29291
rect 40678 29288 40684 29300
rect 40083 29260 40684 29288
rect 40083 29257 40095 29260
rect 40037 29251 40095 29257
rect 40678 29248 40684 29260
rect 40736 29248 40742 29300
rect 41046 29288 41052 29300
rect 41007 29260 41052 29288
rect 41046 29248 41052 29260
rect 41104 29248 41110 29300
rect 45097 29291 45155 29297
rect 45097 29288 45109 29291
rect 43364 29260 45109 29288
rect 42797 29223 42855 29229
rect 42797 29220 42809 29223
rect 36556 29192 42809 29220
rect 42797 29189 42809 29192
rect 42843 29189 42855 29223
rect 42797 29183 42855 29189
rect 35526 29112 35532 29164
rect 35584 29152 35590 29164
rect 38657 29155 38715 29161
rect 35584 29124 37872 29152
rect 35584 29112 35590 29124
rect 31496 29056 31616 29084
rect 14001 29019 14059 29025
rect 14001 29016 14013 29019
rect 12636 28988 14013 29016
rect 14001 28985 14013 28988
rect 14047 28985 14059 29019
rect 14001 28979 14059 28985
rect 17405 29019 17463 29025
rect 17405 28985 17417 29019
rect 17451 29016 17463 29019
rect 31588 29016 31616 29056
rect 31662 29044 31668 29096
rect 31720 29056 31754 29096
rect 31720 29044 31726 29056
rect 34698 29044 34704 29096
rect 34756 29084 34762 29096
rect 34885 29087 34943 29093
rect 34885 29084 34897 29087
rect 34756 29056 34897 29084
rect 34756 29044 34762 29056
rect 34885 29053 34897 29056
rect 34931 29053 34943 29087
rect 34885 29047 34943 29053
rect 37458 29044 37464 29096
rect 37516 29084 37522 29096
rect 37844 29093 37872 29124
rect 38657 29121 38669 29155
rect 38703 29121 38715 29155
rect 39666 29152 39672 29164
rect 39627 29124 39672 29152
rect 38657 29115 38715 29121
rect 37737 29087 37795 29093
rect 37737 29084 37749 29087
rect 37516 29056 37749 29084
rect 37516 29044 37522 29056
rect 37737 29053 37749 29056
rect 37783 29053 37795 29087
rect 37737 29047 37795 29053
rect 37829 29087 37887 29093
rect 37829 29053 37841 29087
rect 37875 29053 37887 29087
rect 37829 29047 37887 29053
rect 32125 29019 32183 29025
rect 32125 29016 32137 29019
rect 17451 28988 18828 29016
rect 31588 28988 32137 29016
rect 17451 28985 17463 28988
rect 17405 28979 17463 28985
rect 16666 28948 16672 28960
rect 16627 28920 16672 28948
rect 16666 28908 16672 28920
rect 16724 28908 16730 28960
rect 18322 28948 18328 28960
rect 18283 28920 18328 28948
rect 18322 28908 18328 28920
rect 18380 28908 18386 28960
rect 18800 28948 18828 28988
rect 32125 28985 32137 28988
rect 32171 28985 32183 29019
rect 32125 28979 32183 28985
rect 36170 28976 36176 29028
rect 36228 29016 36234 29028
rect 36265 29019 36323 29025
rect 36265 29016 36277 29019
rect 36228 28988 36277 29016
rect 36228 28976 36234 28988
rect 36265 28985 36277 28988
rect 36311 29016 36323 29019
rect 38672 29016 38700 29115
rect 39666 29112 39672 29124
rect 39724 29112 39730 29164
rect 40678 29152 40684 29164
rect 40639 29124 40684 29152
rect 40678 29112 40684 29124
rect 40736 29112 40742 29164
rect 42812 29152 42840 29183
rect 43364 29164 43392 29260
rect 45097 29257 45109 29260
rect 45143 29288 45155 29291
rect 45278 29288 45284 29300
rect 45143 29260 45284 29288
rect 45143 29257 45155 29260
rect 45097 29251 45155 29257
rect 45278 29248 45284 29260
rect 45336 29248 45342 29300
rect 43257 29155 43315 29161
rect 43257 29152 43269 29155
rect 42812 29124 43269 29152
rect 43257 29121 43269 29124
rect 43303 29121 43315 29155
rect 43257 29115 43315 29121
rect 43346 29112 43352 29164
rect 43404 29152 43410 29164
rect 43533 29155 43591 29161
rect 43404 29124 43449 29152
rect 43404 29112 43410 29124
rect 43533 29121 43545 29155
rect 43579 29121 43591 29155
rect 43533 29115 43591 29121
rect 44453 29155 44511 29161
rect 44453 29121 44465 29155
rect 44499 29121 44511 29155
rect 44453 29115 44511 29121
rect 44913 29155 44971 29161
rect 44913 29121 44925 29155
rect 44959 29152 44971 29155
rect 45002 29152 45008 29164
rect 44959 29124 45008 29152
rect 44959 29121 44971 29124
rect 44913 29115 44971 29121
rect 38746 29044 38752 29096
rect 38804 29084 38810 29096
rect 39577 29087 39635 29093
rect 39577 29084 39589 29087
rect 38804 29056 38849 29084
rect 39040 29056 39589 29084
rect 38804 29044 38810 29056
rect 39040 29025 39068 29056
rect 39577 29053 39589 29056
rect 39623 29053 39635 29087
rect 39577 29047 39635 29053
rect 40310 29044 40316 29096
rect 40368 29084 40374 29096
rect 40589 29087 40647 29093
rect 40589 29084 40601 29087
rect 40368 29056 40601 29084
rect 40368 29044 40374 29056
rect 40589 29053 40601 29056
rect 40635 29053 40647 29087
rect 40589 29047 40647 29053
rect 42794 29044 42800 29096
rect 42852 29084 42858 29096
rect 43548 29084 43576 29115
rect 42852 29056 43576 29084
rect 44468 29084 44496 29115
rect 45002 29112 45008 29124
rect 45060 29112 45066 29164
rect 45922 29084 45928 29096
rect 44468 29056 45928 29084
rect 42852 29044 42858 29056
rect 45922 29044 45928 29056
rect 45980 29044 45986 29096
rect 36311 28988 38700 29016
rect 39025 29019 39083 29025
rect 36311 28985 36323 28988
rect 36265 28979 36323 28985
rect 39025 28985 39037 29019
rect 39071 28985 39083 29019
rect 39025 28979 39083 28985
rect 43622 28976 43628 29028
rect 43680 29016 43686 29028
rect 43717 29019 43775 29025
rect 43717 29016 43729 29019
rect 43680 28988 43729 29016
rect 43680 28976 43686 28988
rect 43717 28985 43729 28988
rect 43763 28985 43775 29019
rect 43717 28979 43775 28985
rect 19978 28948 19984 28960
rect 18800 28920 19984 28948
rect 19978 28908 19984 28920
rect 20036 28908 20042 28960
rect 21913 28951 21971 28957
rect 21913 28917 21925 28951
rect 21959 28948 21971 28951
rect 22002 28948 22008 28960
rect 21959 28920 22008 28948
rect 21959 28917 21971 28920
rect 21913 28911 21971 28917
rect 22002 28908 22008 28920
rect 22060 28908 22066 28960
rect 24670 28908 24676 28960
rect 24728 28948 24734 28960
rect 24765 28951 24823 28957
rect 24765 28948 24777 28951
rect 24728 28920 24777 28948
rect 24728 28908 24734 28920
rect 24765 28917 24777 28920
rect 24811 28917 24823 28951
rect 30190 28948 30196 28960
rect 30151 28920 30196 28948
rect 24765 28911 24823 28917
rect 30190 28908 30196 28920
rect 30248 28908 30254 28960
rect 43438 28908 43444 28960
rect 43496 28948 43502 28960
rect 44266 28948 44272 28960
rect 43496 28920 44272 28948
rect 43496 28908 43502 28920
rect 44266 28908 44272 28920
rect 44324 28908 44330 28960
rect 1104 28858 68816 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 65654 28858
rect 65706 28806 65718 28858
rect 65770 28806 65782 28858
rect 65834 28806 65846 28858
rect 65898 28806 65910 28858
rect 65962 28806 68816 28858
rect 1104 28784 68816 28806
rect 8941 28747 8999 28753
rect 8941 28713 8953 28747
rect 8987 28744 8999 28747
rect 9122 28744 9128 28756
rect 8987 28716 9128 28744
rect 8987 28713 8999 28716
rect 8941 28707 8999 28713
rect 9122 28704 9128 28716
rect 9180 28704 9186 28756
rect 10137 28747 10195 28753
rect 10137 28713 10149 28747
rect 10183 28744 10195 28747
rect 10318 28744 10324 28756
rect 10183 28716 10324 28744
rect 10183 28713 10195 28716
rect 10137 28707 10195 28713
rect 9125 28611 9183 28617
rect 9125 28577 9137 28611
rect 9171 28608 9183 28611
rect 9674 28608 9680 28620
rect 9171 28580 9680 28608
rect 9171 28577 9183 28580
rect 9125 28571 9183 28577
rect 9674 28568 9680 28580
rect 9732 28608 9738 28620
rect 10152 28608 10180 28707
rect 10318 28704 10324 28716
rect 10376 28744 10382 28756
rect 10965 28747 11023 28753
rect 10965 28744 10977 28747
rect 10376 28716 10977 28744
rect 10376 28704 10382 28716
rect 10965 28713 10977 28716
rect 11011 28744 11023 28747
rect 12618 28744 12624 28756
rect 11011 28716 12624 28744
rect 11011 28713 11023 28716
rect 10965 28707 11023 28713
rect 12618 28704 12624 28716
rect 12676 28704 12682 28756
rect 12713 28747 12771 28753
rect 12713 28713 12725 28747
rect 12759 28744 12771 28747
rect 12802 28744 12808 28756
rect 12759 28716 12808 28744
rect 12759 28713 12771 28716
rect 12713 28707 12771 28713
rect 12802 28704 12808 28716
rect 12860 28704 12866 28756
rect 14090 28744 14096 28756
rect 14051 28716 14096 28744
rect 14090 28704 14096 28716
rect 14148 28704 14154 28756
rect 14550 28744 14556 28756
rect 14511 28716 14556 28744
rect 14550 28704 14556 28716
rect 14608 28704 14614 28756
rect 19242 28744 19248 28756
rect 19203 28716 19248 28744
rect 19242 28704 19248 28716
rect 19300 28704 19306 28756
rect 30834 28744 30840 28756
rect 30795 28716 30840 28744
rect 30834 28704 30840 28716
rect 30892 28704 30898 28756
rect 36446 28744 36452 28756
rect 35084 28716 36452 28744
rect 11698 28636 11704 28688
rect 11756 28636 11762 28688
rect 16666 28676 16672 28688
rect 12176 28648 16672 28676
rect 9732 28580 10180 28608
rect 11716 28608 11744 28636
rect 11716 28580 11928 28608
rect 9732 28568 9738 28580
rect 9217 28543 9275 28549
rect 9217 28509 9229 28543
rect 9263 28540 9275 28543
rect 9582 28540 9588 28552
rect 9263 28512 9588 28540
rect 9263 28509 9275 28512
rect 9217 28503 9275 28509
rect 9582 28500 9588 28512
rect 9640 28500 9646 28552
rect 11606 28540 11612 28552
rect 11567 28512 11612 28540
rect 11606 28500 11612 28512
rect 11664 28500 11670 28552
rect 11900 28549 11928 28580
rect 11702 28543 11760 28549
rect 11702 28509 11714 28543
rect 11748 28509 11760 28543
rect 11702 28503 11760 28509
rect 11885 28543 11943 28549
rect 11885 28509 11897 28543
rect 11931 28509 11943 28543
rect 11885 28503 11943 28509
rect 11146 28432 11152 28484
rect 11204 28472 11210 28484
rect 11716 28472 11744 28503
rect 12066 28500 12072 28552
rect 12124 28549 12130 28552
rect 12124 28540 12132 28549
rect 12176 28540 12204 28648
rect 16666 28636 16672 28648
rect 16724 28636 16730 28688
rect 25406 28636 25412 28688
rect 25464 28676 25470 28688
rect 25464 28648 30420 28676
rect 25464 28636 25470 28648
rect 12618 28568 12624 28620
rect 12676 28608 12682 28620
rect 14182 28608 14188 28620
rect 12676 28580 13216 28608
rect 14143 28580 14188 28608
rect 12676 28568 12682 28580
rect 13188 28549 13216 28580
rect 14182 28568 14188 28580
rect 14240 28568 14246 28620
rect 14734 28568 14740 28620
rect 14792 28608 14798 28620
rect 16485 28611 16543 28617
rect 16485 28608 16497 28611
rect 14792 28580 16497 28608
rect 14792 28568 14798 28580
rect 16485 28577 16497 28580
rect 16531 28577 16543 28611
rect 16485 28571 16543 28577
rect 19889 28611 19947 28617
rect 19889 28577 19901 28611
rect 19935 28608 19947 28611
rect 20254 28608 20260 28620
rect 19935 28580 20260 28608
rect 19935 28577 19947 28580
rect 19889 28571 19947 28577
rect 20254 28568 20260 28580
rect 20312 28568 20318 28620
rect 21726 28608 21732 28620
rect 21687 28580 21732 28608
rect 21726 28568 21732 28580
rect 21784 28568 21790 28620
rect 27801 28611 27859 28617
rect 27801 28577 27813 28611
rect 27847 28577 27859 28611
rect 27801 28571 27859 28577
rect 12897 28543 12955 28549
rect 12897 28540 12909 28543
rect 12124 28512 12204 28540
rect 12268 28512 12909 28540
rect 12124 28503 12132 28512
rect 12124 28500 12130 28503
rect 11204 28444 11744 28472
rect 11204 28432 11210 28444
rect 11974 28432 11980 28484
rect 12032 28472 12038 28484
rect 12032 28444 12077 28472
rect 12032 28432 12038 28444
rect 9306 28364 9312 28416
rect 9364 28404 9370 28416
rect 12268 28413 12296 28512
rect 12897 28509 12909 28512
rect 12943 28509 12955 28543
rect 12897 28503 12955 28509
rect 13173 28543 13231 28549
rect 13173 28509 13185 28543
rect 13219 28540 13231 28543
rect 13538 28540 13544 28552
rect 13219 28512 13544 28540
rect 13219 28509 13231 28512
rect 13173 28503 13231 28509
rect 13538 28500 13544 28512
rect 13596 28500 13602 28552
rect 13998 28500 14004 28552
rect 14056 28540 14062 28552
rect 14093 28543 14151 28549
rect 14093 28540 14105 28543
rect 14056 28512 14105 28540
rect 14056 28500 14062 28512
rect 14093 28509 14105 28512
rect 14139 28509 14151 28543
rect 14366 28540 14372 28552
rect 14327 28512 14372 28540
rect 14093 28503 14151 28509
rect 14366 28500 14372 28512
rect 14424 28500 14430 28552
rect 15194 28540 15200 28552
rect 15155 28512 15200 28540
rect 15194 28500 15200 28512
rect 15252 28500 15258 28552
rect 16025 28543 16083 28549
rect 16025 28509 16037 28543
rect 16071 28540 16083 28543
rect 16758 28540 16764 28552
rect 16071 28512 16764 28540
rect 16071 28509 16083 28512
rect 16025 28503 16083 28509
rect 16758 28500 16764 28512
rect 16816 28500 16822 28552
rect 17773 28543 17831 28549
rect 17773 28509 17785 28543
rect 17819 28540 17831 28543
rect 18322 28540 18328 28552
rect 17819 28512 18328 28540
rect 17819 28509 17831 28512
rect 17773 28503 17831 28509
rect 18322 28500 18328 28512
rect 18380 28500 18386 28552
rect 19058 28500 19064 28552
rect 19116 28540 19122 28552
rect 19705 28543 19763 28549
rect 19705 28540 19717 28543
rect 19116 28512 19717 28540
rect 19116 28500 19122 28512
rect 19705 28509 19717 28512
rect 19751 28540 19763 28543
rect 20070 28540 20076 28552
rect 19751 28512 20076 28540
rect 19751 28509 19763 28512
rect 19705 28503 19763 28509
rect 20070 28500 20076 28512
rect 20128 28500 20134 28552
rect 22002 28549 22008 28552
rect 21996 28540 22008 28549
rect 21963 28512 22008 28540
rect 21996 28503 22008 28512
rect 22002 28500 22008 28503
rect 22060 28500 22066 28552
rect 24394 28540 24400 28552
rect 24355 28512 24400 28540
rect 24394 28500 24400 28512
rect 24452 28500 24458 28552
rect 24670 28549 24676 28552
rect 24664 28540 24676 28549
rect 24631 28512 24676 28540
rect 24664 28503 24676 28512
rect 24670 28500 24676 28503
rect 24728 28500 24734 28552
rect 12434 28432 12440 28484
rect 12492 28472 12498 28484
rect 13081 28475 13139 28481
rect 13081 28472 13093 28475
rect 12492 28444 13093 28472
rect 12492 28432 12498 28444
rect 13081 28441 13093 28444
rect 13127 28472 13139 28475
rect 17034 28472 17040 28484
rect 13127 28444 15240 28472
rect 16995 28444 17040 28472
rect 13127 28441 13139 28444
rect 13081 28435 13139 28441
rect 9585 28407 9643 28413
rect 9585 28404 9597 28407
rect 9364 28376 9597 28404
rect 9364 28364 9370 28376
rect 9585 28373 9597 28376
rect 9631 28373 9643 28407
rect 9585 28367 9643 28373
rect 12253 28407 12311 28413
rect 12253 28373 12265 28407
rect 12299 28373 12311 28407
rect 15212 28404 15240 28444
rect 17034 28432 17040 28444
rect 17092 28432 17098 28484
rect 19613 28475 19671 28481
rect 19613 28472 19625 28475
rect 17604 28444 19625 28472
rect 16669 28407 16727 28413
rect 16669 28404 16681 28407
rect 15212 28376 16681 28404
rect 12253 28367 12311 28373
rect 16669 28373 16681 28376
rect 16715 28373 16727 28407
rect 16669 28367 16727 28373
rect 16853 28407 16911 28413
rect 16853 28373 16865 28407
rect 16899 28404 16911 28407
rect 17126 28404 17132 28416
rect 16899 28376 17132 28404
rect 16899 28373 16911 28376
rect 16853 28367 16911 28373
rect 17126 28364 17132 28376
rect 17184 28364 17190 28416
rect 17494 28364 17500 28416
rect 17552 28404 17558 28416
rect 17604 28413 17632 28444
rect 19613 28441 19625 28444
rect 19659 28472 19671 28475
rect 20533 28475 20591 28481
rect 19659 28444 20484 28472
rect 19659 28441 19671 28444
rect 19613 28435 19671 28441
rect 17589 28407 17647 28413
rect 17589 28404 17601 28407
rect 17552 28376 17601 28404
rect 17552 28364 17558 28376
rect 17589 28373 17601 28376
rect 17635 28373 17647 28407
rect 17589 28367 17647 28373
rect 18322 28364 18328 28416
rect 18380 28404 18386 28416
rect 18417 28407 18475 28413
rect 18417 28404 18429 28407
rect 18380 28376 18429 28404
rect 18380 28364 18386 28376
rect 18417 28373 18429 28376
rect 18463 28404 18475 28407
rect 19242 28404 19248 28416
rect 18463 28376 19248 28404
rect 18463 28373 18475 28376
rect 18417 28367 18475 28373
rect 19242 28364 19248 28376
rect 19300 28364 19306 28416
rect 20456 28404 20484 28444
rect 20533 28441 20545 28475
rect 20579 28472 20591 28475
rect 21082 28472 21088 28484
rect 20579 28444 21088 28472
rect 20579 28441 20591 28444
rect 20533 28435 20591 28441
rect 21082 28432 21088 28444
rect 21140 28432 21146 28484
rect 21266 28432 21272 28484
rect 21324 28472 21330 28484
rect 27816 28472 27844 28571
rect 27893 28543 27951 28549
rect 27893 28509 27905 28543
rect 27939 28540 27951 28543
rect 29638 28540 29644 28552
rect 27939 28512 29644 28540
rect 27939 28509 27951 28512
rect 27893 28503 27951 28509
rect 29638 28500 29644 28512
rect 29696 28500 29702 28552
rect 28810 28472 28816 28484
rect 21324 28444 28816 28472
rect 21324 28432 21330 28444
rect 28810 28432 28816 28444
rect 28868 28432 28874 28484
rect 30392 28481 30420 28648
rect 30926 28568 30932 28620
rect 30984 28608 30990 28620
rect 31294 28608 31300 28620
rect 30984 28580 31300 28608
rect 30984 28568 30990 28580
rect 31294 28568 31300 28580
rect 31352 28608 31358 28620
rect 31389 28611 31447 28617
rect 31389 28608 31401 28611
rect 31352 28580 31401 28608
rect 31352 28568 31358 28580
rect 31389 28577 31401 28580
rect 31435 28577 31447 28611
rect 31389 28571 31447 28577
rect 31478 28568 31484 28620
rect 31536 28608 31542 28620
rect 35084 28617 35112 28716
rect 36446 28704 36452 28716
rect 36504 28744 36510 28756
rect 37182 28744 37188 28756
rect 36504 28716 37188 28744
rect 36504 28704 36510 28716
rect 37182 28704 37188 28716
rect 37240 28704 37246 28756
rect 38473 28679 38531 28685
rect 38473 28645 38485 28679
rect 38519 28676 38531 28679
rect 40678 28676 40684 28688
rect 38519 28648 40684 28676
rect 38519 28645 38531 28648
rect 38473 28639 38531 28645
rect 40678 28636 40684 28648
rect 40736 28636 40742 28688
rect 32217 28611 32275 28617
rect 32217 28608 32229 28611
rect 31536 28580 32229 28608
rect 31536 28568 31542 28580
rect 32217 28577 32229 28580
rect 32263 28577 32275 28611
rect 32217 28571 32275 28577
rect 35069 28611 35127 28617
rect 35069 28577 35081 28611
rect 35115 28577 35127 28611
rect 35069 28571 35127 28577
rect 35986 28568 35992 28620
rect 36044 28608 36050 28620
rect 36081 28611 36139 28617
rect 36081 28608 36093 28611
rect 36044 28580 36093 28608
rect 36044 28568 36050 28580
rect 36081 28577 36093 28580
rect 36127 28577 36139 28611
rect 36081 28571 36139 28577
rect 37458 28568 37464 28620
rect 37516 28608 37522 28620
rect 38013 28611 38071 28617
rect 38013 28608 38025 28611
rect 37516 28580 38025 28608
rect 37516 28568 37522 28580
rect 38013 28577 38025 28580
rect 38059 28577 38071 28611
rect 43346 28608 43352 28620
rect 38013 28571 38071 28577
rect 42996 28580 43352 28608
rect 32309 28543 32367 28549
rect 32309 28509 32321 28543
rect 32355 28540 32367 28543
rect 32582 28540 32588 28552
rect 32355 28512 32588 28540
rect 32355 28509 32367 28512
rect 32309 28503 32367 28509
rect 32582 28500 32588 28512
rect 32640 28500 32646 28552
rect 35161 28543 35219 28549
rect 35161 28509 35173 28543
rect 35207 28540 35219 28543
rect 36170 28540 36176 28552
rect 35207 28512 36176 28540
rect 35207 28509 35219 28512
rect 35161 28503 35219 28509
rect 36170 28500 36176 28512
rect 36228 28500 36234 28552
rect 36354 28549 36360 28552
rect 36348 28540 36360 28549
rect 36315 28512 36360 28540
rect 36348 28503 36360 28512
rect 36354 28500 36360 28503
rect 36412 28500 36418 28552
rect 38102 28540 38108 28552
rect 38063 28512 38108 28540
rect 38102 28500 38108 28512
rect 38160 28540 38166 28552
rect 38933 28543 38991 28549
rect 38933 28540 38945 28543
rect 38160 28512 38945 28540
rect 38160 28500 38166 28512
rect 38933 28509 38945 28512
rect 38979 28509 38991 28543
rect 42242 28540 42248 28552
rect 42203 28512 42248 28540
rect 38933 28503 38991 28509
rect 42242 28500 42248 28512
rect 42300 28540 42306 28552
rect 42794 28540 42800 28552
rect 42300 28512 42800 28540
rect 42300 28500 42306 28512
rect 42794 28500 42800 28512
rect 42852 28500 42858 28552
rect 42996 28549 43024 28580
rect 43346 28568 43352 28580
rect 43404 28568 43410 28620
rect 44266 28568 44272 28620
rect 44324 28608 44330 28620
rect 45005 28611 45063 28617
rect 45005 28608 45017 28611
rect 44324 28580 45017 28608
rect 44324 28568 44330 28580
rect 45005 28577 45017 28580
rect 45051 28577 45063 28611
rect 45005 28571 45063 28577
rect 42981 28543 43039 28549
rect 42981 28509 42993 28543
rect 43027 28509 43039 28543
rect 43438 28540 43444 28552
rect 43399 28512 43444 28540
rect 42981 28503 43039 28509
rect 43438 28500 43444 28512
rect 43496 28500 43502 28552
rect 43717 28543 43775 28549
rect 43717 28509 43729 28543
rect 43763 28509 43775 28543
rect 45278 28540 45284 28552
rect 45239 28512 45284 28540
rect 43717 28503 43775 28509
rect 30377 28475 30435 28481
rect 30377 28441 30389 28475
rect 30423 28472 30435 28475
rect 31205 28475 31263 28481
rect 31205 28472 31217 28475
rect 30423 28444 31217 28472
rect 30423 28441 30435 28444
rect 30377 28435 30435 28441
rect 31205 28441 31217 28444
rect 31251 28472 31263 28475
rect 36078 28472 36084 28484
rect 31251 28444 36084 28472
rect 31251 28441 31263 28444
rect 31205 28435 31263 28441
rect 36078 28432 36084 28444
rect 36136 28432 36142 28484
rect 42889 28475 42947 28481
rect 42889 28441 42901 28475
rect 42935 28472 42947 28475
rect 43732 28472 43760 28503
rect 45278 28500 45284 28512
rect 45336 28500 45342 28552
rect 46109 28543 46167 28549
rect 46109 28509 46121 28543
rect 46155 28540 46167 28543
rect 54570 28540 54576 28552
rect 46155 28512 54576 28540
rect 46155 28509 46167 28512
rect 46109 28503 46167 28509
rect 54570 28500 54576 28512
rect 54628 28540 54634 28552
rect 67174 28540 67180 28552
rect 54628 28512 67180 28540
rect 54628 28500 54634 28512
rect 67174 28500 67180 28512
rect 67232 28500 67238 28552
rect 42935 28444 43760 28472
rect 42935 28441 42947 28444
rect 42889 28435 42947 28441
rect 20898 28404 20904 28416
rect 20456 28376 20904 28404
rect 20898 28364 20904 28376
rect 20956 28364 20962 28416
rect 21177 28407 21235 28413
rect 21177 28373 21189 28407
rect 21223 28404 21235 28407
rect 22462 28404 22468 28416
rect 21223 28376 22468 28404
rect 21223 28373 21235 28376
rect 21177 28367 21235 28373
rect 22462 28364 22468 28376
rect 22520 28364 22526 28416
rect 23106 28404 23112 28416
rect 23067 28376 23112 28404
rect 23106 28364 23112 28376
rect 23164 28364 23170 28416
rect 25038 28364 25044 28416
rect 25096 28404 25102 28416
rect 25777 28407 25835 28413
rect 25777 28404 25789 28407
rect 25096 28376 25789 28404
rect 25096 28364 25102 28376
rect 25777 28373 25789 28376
rect 25823 28373 25835 28407
rect 28258 28404 28264 28416
rect 28219 28376 28264 28404
rect 25777 28367 25835 28373
rect 28258 28364 28264 28376
rect 28316 28364 28322 28416
rect 31297 28407 31355 28413
rect 31297 28373 31309 28407
rect 31343 28404 31355 28407
rect 31386 28404 31392 28416
rect 31343 28376 31392 28404
rect 31343 28373 31355 28376
rect 31297 28367 31355 28373
rect 31386 28364 31392 28376
rect 31444 28364 31450 28416
rect 32677 28407 32735 28413
rect 32677 28373 32689 28407
rect 32723 28404 32735 28407
rect 33410 28404 33416 28416
rect 32723 28376 33416 28404
rect 32723 28373 32735 28376
rect 32677 28367 32735 28373
rect 33410 28364 33416 28376
rect 33468 28364 33474 28416
rect 34790 28364 34796 28416
rect 34848 28404 34854 28416
rect 35253 28407 35311 28413
rect 35253 28404 35265 28407
rect 34848 28376 35265 28404
rect 34848 28364 34854 28376
rect 35253 28373 35265 28376
rect 35299 28373 35311 28407
rect 35618 28404 35624 28416
rect 35579 28376 35624 28404
rect 35253 28367 35311 28373
rect 35618 28364 35624 28376
rect 35676 28364 35682 28416
rect 37458 28404 37464 28416
rect 37419 28376 37464 28404
rect 37458 28364 37464 28376
rect 37516 28364 37522 28416
rect 43990 28364 43996 28416
rect 44048 28404 44054 28416
rect 44453 28407 44511 28413
rect 44453 28404 44465 28407
rect 44048 28376 44465 28404
rect 44048 28364 44054 28376
rect 44453 28373 44465 28376
rect 44499 28373 44511 28407
rect 44453 28367 44511 28373
rect 1104 28314 68816 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 68816 28314
rect 1104 28240 68816 28262
rect 6917 28203 6975 28209
rect 6917 28169 6929 28203
rect 6963 28200 6975 28203
rect 7006 28200 7012 28212
rect 6963 28172 7012 28200
rect 6963 28169 6975 28172
rect 6917 28163 6975 28169
rect 7006 28160 7012 28172
rect 7064 28160 7070 28212
rect 9950 28160 9956 28212
rect 10008 28200 10014 28212
rect 10413 28203 10471 28209
rect 10413 28200 10425 28203
rect 10008 28172 10425 28200
rect 10008 28160 10014 28172
rect 10413 28169 10425 28172
rect 10459 28200 10471 28203
rect 10962 28200 10968 28212
rect 10459 28172 10968 28200
rect 10459 28169 10471 28172
rect 10413 28163 10471 28169
rect 10962 28160 10968 28172
rect 11020 28160 11026 28212
rect 11701 28203 11759 28209
rect 11701 28169 11713 28203
rect 11747 28200 11759 28203
rect 11790 28200 11796 28212
rect 11747 28172 11796 28200
rect 11747 28169 11759 28172
rect 11701 28163 11759 28169
rect 11790 28160 11796 28172
rect 11848 28160 11854 28212
rect 11974 28160 11980 28212
rect 12032 28200 12038 28212
rect 12621 28203 12679 28209
rect 12621 28200 12633 28203
rect 12032 28172 12633 28200
rect 12032 28160 12038 28172
rect 12621 28169 12633 28172
rect 12667 28169 12679 28203
rect 12621 28163 12679 28169
rect 14185 28203 14243 28209
rect 14185 28169 14197 28203
rect 14231 28200 14243 28203
rect 14366 28200 14372 28212
rect 14231 28172 14372 28200
rect 14231 28169 14243 28172
rect 14185 28163 14243 28169
rect 14366 28160 14372 28172
rect 14424 28160 14430 28212
rect 15194 28160 15200 28212
rect 15252 28200 15258 28212
rect 15565 28203 15623 28209
rect 15565 28200 15577 28203
rect 15252 28172 15577 28200
rect 15252 28160 15258 28172
rect 15565 28169 15577 28172
rect 15611 28200 15623 28203
rect 20162 28200 20168 28212
rect 15611 28172 16160 28200
rect 20123 28172 20168 28200
rect 15611 28169 15623 28172
rect 15565 28163 15623 28169
rect 14274 28092 14280 28144
rect 14332 28132 14338 28144
rect 16132 28132 16160 28172
rect 20162 28160 20168 28172
rect 20220 28160 20226 28212
rect 21266 28200 21272 28212
rect 21227 28172 21272 28200
rect 21266 28160 21272 28172
rect 21324 28160 21330 28212
rect 22094 28160 22100 28212
rect 22152 28200 22158 28212
rect 22557 28203 22615 28209
rect 22152 28172 22197 28200
rect 22152 28160 22158 28172
rect 22557 28169 22569 28203
rect 22603 28200 22615 28203
rect 23106 28200 23112 28212
rect 22603 28172 23112 28200
rect 22603 28169 22615 28172
rect 22557 28163 22615 28169
rect 23106 28160 23112 28172
rect 23164 28160 23170 28212
rect 23385 28203 23443 28209
rect 23385 28169 23397 28203
rect 23431 28200 23443 28203
rect 23842 28200 23848 28212
rect 23431 28172 23848 28200
rect 23431 28169 23443 28172
rect 23385 28163 23443 28169
rect 23842 28160 23848 28172
rect 23900 28160 23906 28212
rect 24397 28203 24455 28209
rect 24397 28169 24409 28203
rect 24443 28200 24455 28203
rect 24578 28200 24584 28212
rect 24443 28172 24584 28200
rect 24443 28169 24455 28172
rect 24397 28163 24455 28169
rect 24578 28160 24584 28172
rect 24636 28160 24642 28212
rect 24765 28203 24823 28209
rect 24765 28169 24777 28203
rect 24811 28200 24823 28203
rect 24854 28200 24860 28212
rect 24811 28172 24860 28200
rect 24811 28169 24823 28172
rect 24765 28163 24823 28169
rect 24854 28160 24860 28172
rect 24912 28200 24918 28212
rect 27341 28203 27399 28209
rect 27341 28200 27353 28203
rect 24912 28172 27353 28200
rect 24912 28160 24918 28172
rect 27341 28169 27353 28172
rect 27387 28200 27399 28203
rect 31205 28203 31263 28209
rect 31205 28200 31217 28203
rect 27387 28172 31217 28200
rect 27387 28169 27399 28172
rect 27341 28163 27399 28169
rect 31205 28169 31217 28172
rect 31251 28200 31263 28203
rect 31294 28200 31300 28212
rect 31251 28172 31300 28200
rect 31251 28169 31263 28172
rect 31205 28163 31263 28169
rect 31294 28160 31300 28172
rect 31352 28160 31358 28212
rect 31573 28203 31631 28209
rect 31573 28169 31585 28203
rect 31619 28200 31631 28203
rect 31662 28200 31668 28212
rect 31619 28172 31668 28200
rect 31619 28169 31631 28172
rect 31573 28163 31631 28169
rect 31662 28160 31668 28172
rect 31720 28160 31726 28212
rect 32677 28203 32735 28209
rect 32677 28169 32689 28203
rect 32723 28169 32735 28203
rect 32677 28163 32735 28169
rect 35069 28203 35127 28209
rect 35069 28169 35081 28203
rect 35115 28200 35127 28203
rect 35342 28200 35348 28212
rect 35115 28172 35348 28200
rect 35115 28169 35127 28172
rect 35069 28163 35127 28169
rect 32692 28132 32720 28163
rect 35342 28160 35348 28172
rect 35400 28160 35406 28212
rect 35894 28160 35900 28212
rect 35952 28200 35958 28212
rect 35989 28203 36047 28209
rect 35989 28200 36001 28203
rect 35952 28172 36001 28200
rect 35952 28160 35958 28172
rect 35989 28169 36001 28172
rect 36035 28169 36047 28203
rect 35989 28163 36047 28169
rect 36449 28203 36507 28209
rect 36449 28169 36461 28203
rect 36495 28200 36507 28203
rect 37366 28200 37372 28212
rect 36495 28172 37372 28200
rect 36495 28169 36507 28172
rect 36449 28163 36507 28169
rect 37366 28160 37372 28172
rect 37424 28160 37430 28212
rect 37826 28200 37832 28212
rect 37787 28172 37832 28200
rect 37826 28160 37832 28172
rect 37884 28160 37890 28212
rect 38105 28203 38163 28209
rect 38105 28169 38117 28203
rect 38151 28200 38163 28203
rect 45462 28200 45468 28212
rect 38151 28172 45468 28200
rect 38151 28169 38163 28172
rect 38105 28163 38163 28169
rect 45462 28160 45468 28172
rect 45520 28160 45526 28212
rect 45922 28200 45928 28212
rect 45883 28172 45928 28200
rect 45922 28160 45928 28172
rect 45980 28160 45986 28212
rect 33137 28135 33195 28141
rect 33137 28132 33149 28135
rect 14332 28104 15700 28132
rect 16132 28104 32628 28132
rect 32692 28104 33149 28132
rect 14332 28092 14338 28104
rect 5902 28024 5908 28076
rect 5960 28064 5966 28076
rect 6549 28067 6607 28073
rect 6549 28064 6561 28067
rect 5960 28036 6561 28064
rect 5960 28024 5966 28036
rect 6549 28033 6561 28036
rect 6595 28064 6607 28067
rect 7377 28067 7435 28073
rect 7377 28064 7389 28067
rect 6595 28036 7389 28064
rect 6595 28033 6607 28036
rect 6549 28027 6607 28033
rect 7377 28033 7389 28036
rect 7423 28033 7435 28067
rect 7377 28027 7435 28033
rect 10781 28067 10839 28073
rect 10781 28033 10793 28067
rect 10827 28033 10839 28067
rect 10781 28027 10839 28033
rect 6454 27996 6460 28008
rect 6415 27968 6460 27996
rect 6454 27956 6460 27968
rect 6512 27956 6518 28008
rect 10689 27999 10747 28005
rect 10689 27965 10701 27999
rect 10735 27965 10747 27999
rect 10796 27996 10824 28027
rect 11054 28024 11060 28076
rect 11112 28064 11118 28076
rect 11609 28067 11667 28073
rect 11609 28064 11621 28067
rect 11112 28036 11621 28064
rect 11112 28024 11118 28036
rect 11609 28033 11621 28036
rect 11655 28033 11667 28067
rect 11609 28027 11667 28033
rect 11885 28067 11943 28073
rect 11885 28033 11897 28067
rect 11931 28064 11943 28067
rect 12066 28064 12072 28076
rect 11931 28036 12072 28064
rect 11931 28033 11943 28036
rect 11885 28027 11943 28033
rect 12066 28024 12072 28036
rect 12124 28024 12130 28076
rect 12158 28024 12164 28076
rect 12216 28064 12222 28076
rect 12529 28067 12587 28073
rect 12529 28064 12541 28067
rect 12216 28036 12541 28064
rect 12216 28024 12222 28036
rect 12529 28033 12541 28036
rect 12575 28033 12587 28067
rect 12529 28027 12587 28033
rect 12713 28067 12771 28073
rect 12713 28033 12725 28067
rect 12759 28064 12771 28067
rect 12986 28064 12992 28076
rect 12759 28036 12992 28064
rect 12759 28033 12771 28036
rect 12713 28027 12771 28033
rect 12986 28024 12992 28036
rect 13044 28024 13050 28076
rect 14553 28067 14611 28073
rect 14553 28033 14565 28067
rect 14599 28033 14611 28067
rect 14553 28027 14611 28033
rect 11238 27996 11244 28008
rect 10796 27968 11244 27996
rect 10689 27959 10747 27965
rect 10704 27928 10732 27959
rect 11238 27956 11244 27968
rect 11296 27956 11302 28008
rect 11698 27928 11704 27940
rect 10704 27900 11704 27928
rect 11698 27888 11704 27900
rect 11756 27928 11762 27940
rect 12158 27928 12164 27940
rect 11756 27900 12164 27928
rect 11756 27888 11762 27900
rect 12158 27888 12164 27900
rect 12216 27888 12222 27940
rect 14568 27928 14596 28027
rect 15286 28024 15292 28076
rect 15344 28064 15350 28076
rect 15672 28073 15700 28104
rect 15381 28067 15439 28073
rect 15381 28064 15393 28067
rect 15344 28036 15393 28064
rect 15344 28024 15350 28036
rect 15381 28033 15393 28036
rect 15427 28033 15439 28067
rect 15381 28027 15439 28033
rect 15657 28067 15715 28073
rect 15657 28033 15669 28067
rect 15703 28033 15715 28067
rect 15657 28027 15715 28033
rect 17773 28067 17831 28073
rect 17773 28033 17785 28067
rect 17819 28064 17831 28067
rect 18877 28067 18935 28073
rect 18877 28064 18889 28067
rect 17819 28036 18889 28064
rect 17819 28033 17831 28036
rect 17773 28027 17831 28033
rect 18877 28033 18889 28036
rect 18923 28064 18935 28067
rect 19242 28064 19248 28076
rect 18923 28036 19248 28064
rect 18923 28033 18935 28036
rect 18877 28027 18935 28033
rect 19242 28024 19248 28036
rect 19300 28064 19306 28076
rect 19337 28067 19395 28073
rect 19337 28064 19349 28067
rect 19300 28036 19349 28064
rect 19300 28024 19306 28036
rect 19337 28033 19349 28036
rect 19383 28033 19395 28067
rect 19337 28027 19395 28033
rect 20162 28024 20168 28076
rect 20220 28064 20226 28076
rect 20901 28067 20959 28073
rect 20901 28064 20913 28067
rect 20220 28036 20913 28064
rect 20220 28024 20226 28036
rect 20901 28033 20913 28036
rect 20947 28033 20959 28067
rect 22462 28064 22468 28076
rect 22375 28036 22468 28064
rect 20901 28027 20959 28033
rect 22462 28024 22468 28036
rect 22520 28064 22526 28076
rect 23842 28064 23848 28076
rect 22520 28036 23848 28064
rect 22520 28024 22526 28036
rect 23842 28024 23848 28036
rect 23900 28024 23906 28076
rect 24857 28067 24915 28073
rect 24857 28033 24869 28067
rect 24903 28064 24915 28067
rect 25038 28064 25044 28076
rect 24903 28036 25044 28064
rect 24903 28033 24915 28036
rect 24857 28027 24915 28033
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28064 26295 28067
rect 28350 28064 28356 28076
rect 26283 28036 27016 28064
rect 28311 28036 28356 28064
rect 26283 28033 26295 28036
rect 26237 28027 26295 28033
rect 14645 27999 14703 28005
rect 14645 27965 14657 27999
rect 14691 27996 14703 27999
rect 15197 27999 15255 28005
rect 15197 27996 15209 27999
rect 14691 27968 15209 27996
rect 14691 27965 14703 27968
rect 14645 27959 14703 27965
rect 15197 27965 15209 27968
rect 15243 27965 15255 27999
rect 15197 27959 15255 27965
rect 19426 27956 19432 28008
rect 19484 27996 19490 28008
rect 20809 27999 20867 28005
rect 20809 27996 20821 27999
rect 19484 27968 20821 27996
rect 19484 27956 19490 27968
rect 20809 27965 20821 27968
rect 20855 27965 20867 27999
rect 22738 27996 22744 28008
rect 22651 27968 22744 27996
rect 20809 27959 20867 27965
rect 22738 27956 22744 27968
rect 22796 27996 22802 28008
rect 24210 27996 24216 28008
rect 22796 27968 24216 27996
rect 22796 27956 22802 27968
rect 24210 27956 24216 27968
rect 24268 27996 24274 28008
rect 24949 27999 25007 28005
rect 24949 27996 24961 27999
rect 24268 27968 24961 27996
rect 24268 27956 24274 27968
rect 24949 27965 24961 27968
rect 24995 27965 25007 27999
rect 24949 27959 25007 27965
rect 15562 27928 15568 27940
rect 14568 27900 15568 27928
rect 15562 27888 15568 27900
rect 15620 27888 15626 27940
rect 19521 27931 19579 27937
rect 19521 27897 19533 27931
rect 19567 27928 19579 27931
rect 19978 27928 19984 27940
rect 19567 27900 19984 27928
rect 19567 27897 19579 27900
rect 19521 27891 19579 27897
rect 19978 27888 19984 27900
rect 20036 27928 20042 27940
rect 26988 27937 27016 28036
rect 28350 28024 28356 28036
rect 28408 28024 28414 28076
rect 30009 28067 30067 28073
rect 30009 28033 30021 28067
rect 30055 28064 30067 28067
rect 30190 28064 30196 28076
rect 30055 28036 30196 28064
rect 30055 28033 30067 28036
rect 30009 28027 30067 28033
rect 30190 28024 30196 28036
rect 30248 28064 30254 28076
rect 31113 28067 31171 28073
rect 31113 28064 31125 28067
rect 30248 28036 31125 28064
rect 30248 28024 30254 28036
rect 31113 28033 31125 28036
rect 31159 28033 31171 28067
rect 32306 28064 32312 28076
rect 32267 28036 32312 28064
rect 31113 28027 31171 28033
rect 32306 28024 32312 28036
rect 32364 28024 32370 28076
rect 32600 28064 32628 28104
rect 33137 28101 33149 28104
rect 33183 28101 33195 28135
rect 37277 28135 37335 28141
rect 37277 28132 37289 28135
rect 33137 28095 33195 28101
rect 33244 28104 37289 28132
rect 33244 28064 33272 28104
rect 37277 28101 37289 28104
rect 37323 28132 37335 28135
rect 38013 28135 38071 28141
rect 38013 28132 38025 28135
rect 37323 28104 38025 28132
rect 37323 28101 37335 28104
rect 37277 28095 37335 28101
rect 38013 28101 38025 28104
rect 38059 28101 38071 28135
rect 38013 28095 38071 28101
rect 38565 28135 38623 28141
rect 38565 28101 38577 28135
rect 38611 28132 38623 28135
rect 43990 28132 43996 28144
rect 38611 28104 43576 28132
rect 43951 28104 43996 28132
rect 38611 28101 38623 28104
rect 38565 28095 38623 28101
rect 33410 28064 33416 28076
rect 32600 28036 33272 28064
rect 33371 28036 33416 28064
rect 33410 28024 33416 28036
rect 33468 28024 33474 28076
rect 35253 28067 35311 28073
rect 35253 28033 35265 28067
rect 35299 28064 35311 28067
rect 35618 28064 35624 28076
rect 35299 28036 35624 28064
rect 35299 28033 35311 28036
rect 35253 28027 35311 28033
rect 35618 28024 35624 28036
rect 35676 28024 35682 28076
rect 36078 28024 36084 28076
rect 36136 28064 36142 28076
rect 36357 28067 36415 28073
rect 36357 28064 36369 28067
rect 36136 28036 36369 28064
rect 36136 28024 36142 28036
rect 36357 28033 36369 28036
rect 36403 28064 36415 28067
rect 40865 28067 40923 28073
rect 40865 28064 40877 28067
rect 36403 28036 40877 28064
rect 36403 28033 36415 28036
rect 36357 28027 36415 28033
rect 40865 28033 40877 28036
rect 40911 28064 40923 28067
rect 40911 28036 41414 28064
rect 40911 28033 40923 28036
rect 40865 28027 40923 28033
rect 27338 27956 27344 28008
rect 27396 27996 27402 28008
rect 27433 27999 27491 28005
rect 27433 27996 27445 27999
rect 27396 27968 27445 27996
rect 27396 27956 27402 27968
rect 27433 27965 27445 27968
rect 27479 27965 27491 27999
rect 27433 27959 27491 27965
rect 27522 27956 27528 28008
rect 27580 27996 27586 28008
rect 28258 27996 28264 28008
rect 27580 27968 27625 27996
rect 28219 27968 28264 27996
rect 27580 27956 27586 27968
rect 28258 27956 28264 27968
rect 28316 27956 28322 28008
rect 29638 27956 29644 28008
rect 29696 27996 29702 28008
rect 29917 27999 29975 28005
rect 29917 27996 29929 27999
rect 29696 27968 29929 27996
rect 29696 27956 29702 27968
rect 29917 27965 29929 27968
rect 29963 27965 29975 27999
rect 30926 27996 30932 28008
rect 30887 27968 30932 27996
rect 29917 27959 29975 27965
rect 30926 27956 30932 27968
rect 30984 27956 30990 28008
rect 31018 27956 31024 28008
rect 31076 27996 31082 28008
rect 32217 27999 32275 28005
rect 32217 27996 32229 27999
rect 31076 27968 32229 27996
rect 31076 27956 31082 27968
rect 32217 27965 32229 27968
rect 32263 27965 32275 27999
rect 32217 27959 32275 27965
rect 33229 27999 33287 28005
rect 33229 27965 33241 27999
rect 33275 27965 33287 27999
rect 33229 27959 33287 27965
rect 26973 27931 27031 27937
rect 20036 27900 26924 27928
rect 20036 27888 20042 27900
rect 8294 27820 8300 27872
rect 8352 27860 8358 27872
rect 8849 27863 8907 27869
rect 8849 27860 8861 27863
rect 8352 27832 8861 27860
rect 8352 27820 8358 27832
rect 8849 27829 8861 27832
rect 8895 27829 8907 27863
rect 8849 27823 8907 27829
rect 12069 27863 12127 27869
rect 12069 27829 12081 27863
rect 12115 27860 12127 27863
rect 12802 27860 12808 27872
rect 12115 27832 12808 27860
rect 12115 27829 12127 27832
rect 12069 27823 12127 27829
rect 12802 27820 12808 27832
rect 12860 27820 12866 27872
rect 13357 27863 13415 27869
rect 13357 27829 13369 27863
rect 13403 27860 13415 27863
rect 13538 27860 13544 27872
rect 13403 27832 13544 27860
rect 13403 27829 13415 27832
rect 13357 27823 13415 27829
rect 13538 27820 13544 27832
rect 13596 27820 13602 27872
rect 17126 27820 17132 27872
rect 17184 27860 17190 27872
rect 17221 27863 17279 27869
rect 17221 27860 17233 27863
rect 17184 27832 17233 27860
rect 17184 27820 17190 27832
rect 17221 27829 17233 27832
rect 17267 27860 17279 27863
rect 17678 27860 17684 27872
rect 17267 27832 17684 27860
rect 17267 27829 17279 27832
rect 17221 27823 17279 27829
rect 17678 27820 17684 27832
rect 17736 27820 17742 27872
rect 18325 27863 18383 27869
rect 18325 27829 18337 27863
rect 18371 27860 18383 27863
rect 19058 27860 19064 27872
rect 18371 27832 19064 27860
rect 18371 27829 18383 27832
rect 18325 27823 18383 27829
rect 19058 27820 19064 27832
rect 19116 27820 19122 27872
rect 26053 27863 26111 27869
rect 26053 27829 26065 27863
rect 26099 27860 26111 27863
rect 26234 27860 26240 27872
rect 26099 27832 26240 27860
rect 26099 27829 26111 27832
rect 26053 27823 26111 27829
rect 26234 27820 26240 27832
rect 26292 27820 26298 27872
rect 26896 27860 26924 27900
rect 26973 27897 26985 27931
rect 27019 27897 27031 27931
rect 30282 27928 30288 27940
rect 26973 27891 27031 27897
rect 28552 27900 30288 27928
rect 28552 27860 28580 27900
rect 30282 27888 30288 27900
rect 30340 27888 30346 27940
rect 30377 27931 30435 27937
rect 30377 27897 30389 27931
rect 30423 27928 30435 27931
rect 31202 27928 31208 27940
rect 30423 27900 31208 27928
rect 30423 27897 30435 27900
rect 30377 27891 30435 27897
rect 31202 27888 31208 27900
rect 31260 27888 31266 27940
rect 33244 27928 33272 27959
rect 35526 27956 35532 28008
rect 35584 27996 35590 28008
rect 36541 27999 36599 28005
rect 36541 27996 36553 27999
rect 35584 27968 36553 27996
rect 35584 27956 35590 27968
rect 36541 27965 36553 27968
rect 36587 27965 36599 27999
rect 36541 27959 36599 27965
rect 37366 27956 37372 28008
rect 37424 27996 37430 28008
rect 39298 27996 39304 28008
rect 37424 27968 39304 27996
rect 37424 27956 37430 27968
rect 39298 27956 39304 27968
rect 39356 27956 39362 28008
rect 31312 27900 33272 27928
rect 26896 27832 28580 27860
rect 28629 27863 28687 27869
rect 28629 27829 28641 27863
rect 28675 27860 28687 27863
rect 31312 27860 31340 27900
rect 37918 27888 37924 27940
rect 37976 27928 37982 27940
rect 38565 27931 38623 27937
rect 38565 27928 38577 27931
rect 37976 27900 38577 27928
rect 37976 27888 37982 27900
rect 38565 27897 38577 27900
rect 38611 27897 38623 27931
rect 38565 27891 38623 27897
rect 41386 27872 41414 28036
rect 43548 27996 43576 28104
rect 43990 28092 43996 28104
rect 44048 28092 44054 28144
rect 45830 28132 45836 28144
rect 45218 28104 45836 28132
rect 45830 28092 45836 28104
rect 45888 28092 45894 28144
rect 43714 28064 43720 28076
rect 43675 28036 43720 28064
rect 43714 28024 43720 28036
rect 43772 28024 43778 28076
rect 45462 28024 45468 28076
rect 45520 28064 45526 28076
rect 46109 28067 46167 28073
rect 46109 28064 46121 28067
rect 45520 28036 46121 28064
rect 45520 28024 45526 28036
rect 46109 28033 46121 28036
rect 46155 28033 46167 28067
rect 46109 28027 46167 28033
rect 45186 27996 45192 28008
rect 43548 27968 45192 27996
rect 45186 27956 45192 27968
rect 45244 27996 45250 28008
rect 46293 27999 46351 28005
rect 46293 27996 46305 27999
rect 45244 27968 46305 27996
rect 45244 27956 45250 27968
rect 46293 27965 46305 27968
rect 46339 27965 46351 27999
rect 46293 27959 46351 27965
rect 28675 27832 31340 27860
rect 28675 27829 28687 27832
rect 28629 27823 28687 27829
rect 32398 27820 32404 27872
rect 32456 27860 32462 27872
rect 33137 27863 33195 27869
rect 33137 27860 33149 27863
rect 32456 27832 33149 27860
rect 32456 27820 32462 27832
rect 33137 27829 33149 27832
rect 33183 27829 33195 27863
rect 33594 27860 33600 27872
rect 33555 27832 33600 27860
rect 33137 27823 33195 27829
rect 33594 27820 33600 27832
rect 33652 27820 33658 27872
rect 41386 27832 41420 27872
rect 41414 27820 41420 27832
rect 41472 27820 41478 27872
rect 1104 27770 68816 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 65654 27770
rect 65706 27718 65718 27770
rect 65770 27718 65782 27770
rect 65834 27718 65846 27770
rect 65898 27718 65910 27770
rect 65962 27718 68816 27770
rect 1104 27696 68816 27718
rect 6454 27656 6460 27668
rect 6415 27628 6460 27656
rect 6454 27616 6460 27628
rect 6512 27616 6518 27668
rect 11606 27616 11612 27668
rect 11664 27656 11670 27668
rect 11701 27659 11759 27665
rect 11701 27656 11713 27659
rect 11664 27628 11713 27656
rect 11664 27616 11670 27628
rect 11701 27625 11713 27628
rect 11747 27625 11759 27659
rect 11701 27619 11759 27625
rect 19242 27616 19248 27668
rect 19300 27656 19306 27668
rect 22554 27656 22560 27668
rect 19300 27628 22560 27656
rect 19300 27616 19306 27628
rect 22554 27616 22560 27628
rect 22612 27616 22618 27668
rect 27893 27659 27951 27665
rect 27893 27625 27905 27659
rect 27939 27656 27951 27659
rect 28350 27656 28356 27668
rect 27939 27628 28356 27656
rect 27939 27625 27951 27628
rect 27893 27619 27951 27625
rect 28350 27616 28356 27628
rect 28408 27616 28414 27668
rect 31294 27616 31300 27668
rect 31352 27656 31358 27668
rect 34606 27656 34612 27668
rect 31352 27628 34612 27656
rect 31352 27616 31358 27628
rect 34606 27616 34612 27628
rect 34664 27656 34670 27668
rect 34790 27656 34796 27668
rect 34664 27628 34796 27656
rect 34664 27616 34670 27628
rect 34790 27616 34796 27628
rect 34848 27616 34854 27668
rect 35897 27659 35955 27665
rect 35897 27625 35909 27659
rect 35943 27656 35955 27659
rect 36078 27656 36084 27668
rect 35943 27628 36084 27656
rect 35943 27625 35955 27628
rect 35897 27619 35955 27625
rect 36078 27616 36084 27628
rect 36136 27616 36142 27668
rect 37918 27656 37924 27668
rect 37879 27628 37924 27656
rect 37918 27616 37924 27628
rect 37976 27616 37982 27668
rect 9217 27591 9275 27597
rect 9217 27557 9229 27591
rect 9263 27588 9275 27591
rect 11146 27588 11152 27600
rect 9263 27560 11152 27588
rect 9263 27557 9275 27560
rect 9217 27551 9275 27557
rect 11146 27548 11152 27560
rect 11204 27548 11210 27600
rect 18601 27591 18659 27597
rect 18601 27557 18613 27591
rect 18647 27588 18659 27591
rect 19426 27588 19432 27600
rect 18647 27560 19432 27588
rect 18647 27557 18659 27560
rect 18601 27551 18659 27557
rect 19426 27548 19432 27560
rect 19484 27548 19490 27600
rect 20346 27548 20352 27600
rect 20404 27588 20410 27600
rect 20717 27591 20775 27597
rect 20717 27588 20729 27591
rect 20404 27560 20729 27588
rect 20404 27548 20410 27560
rect 20717 27557 20729 27560
rect 20763 27557 20775 27591
rect 20717 27551 20775 27557
rect 20901 27591 20959 27597
rect 20901 27557 20913 27591
rect 20947 27588 20959 27591
rect 20947 27560 22508 27588
rect 20947 27557 20959 27560
rect 20901 27551 20959 27557
rect 9950 27520 9956 27532
rect 9911 27492 9956 27520
rect 9950 27480 9956 27492
rect 10008 27480 10014 27532
rect 15013 27523 15071 27529
rect 15013 27489 15025 27523
rect 15059 27520 15071 27523
rect 15102 27520 15108 27532
rect 15059 27492 15108 27520
rect 15059 27489 15071 27492
rect 15013 27483 15071 27489
rect 15102 27480 15108 27492
rect 15160 27480 15166 27532
rect 4433 27455 4491 27461
rect 4433 27421 4445 27455
rect 4479 27452 4491 27455
rect 4798 27452 4804 27464
rect 4479 27424 4804 27452
rect 4479 27421 4491 27424
rect 4433 27415 4491 27421
rect 4798 27412 4804 27424
rect 4856 27412 4862 27464
rect 5074 27452 5080 27464
rect 5035 27424 5080 27452
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 7101 27455 7159 27461
rect 7101 27421 7113 27455
rect 7147 27452 7159 27455
rect 7374 27452 7380 27464
rect 7147 27424 7380 27452
rect 7147 27421 7159 27424
rect 7101 27415 7159 27421
rect 7374 27412 7380 27424
rect 7432 27412 7438 27464
rect 8754 27412 8760 27464
rect 8812 27452 8818 27464
rect 8941 27455 8999 27461
rect 8941 27452 8953 27455
rect 8812 27424 8953 27452
rect 8812 27412 8818 27424
rect 8941 27421 8953 27424
rect 8987 27421 8999 27455
rect 9861 27455 9919 27461
rect 9861 27452 9873 27455
rect 8941 27415 8999 27421
rect 9048 27424 9873 27452
rect 5344 27387 5402 27393
rect 5344 27353 5356 27387
rect 5390 27384 5402 27387
rect 5994 27384 6000 27396
rect 5390 27356 6000 27384
rect 5390 27353 5402 27356
rect 5344 27347 5402 27353
rect 5994 27344 6000 27356
rect 6052 27344 6058 27396
rect 7742 27344 7748 27396
rect 7800 27384 7806 27396
rect 9048 27384 9076 27424
rect 9861 27421 9873 27424
rect 9907 27421 9919 27455
rect 9861 27415 9919 27421
rect 11054 27412 11060 27464
rect 11112 27452 11118 27464
rect 11517 27455 11575 27461
rect 11517 27452 11529 27455
rect 11112 27424 11529 27452
rect 11112 27412 11118 27424
rect 11517 27421 11529 27424
rect 11563 27421 11575 27455
rect 11698 27452 11704 27464
rect 11659 27424 11704 27452
rect 11517 27415 11575 27421
rect 9214 27384 9220 27396
rect 7800 27356 9076 27384
rect 9175 27356 9220 27384
rect 7800 27344 7806 27356
rect 9214 27344 9220 27356
rect 9272 27344 9278 27396
rect 11532 27384 11560 27415
rect 11698 27412 11704 27424
rect 11756 27412 11762 27464
rect 14734 27452 14740 27464
rect 14695 27424 14740 27452
rect 14734 27412 14740 27424
rect 14792 27412 14798 27464
rect 14921 27455 14979 27461
rect 14921 27421 14933 27455
rect 14967 27452 14979 27455
rect 15194 27452 15200 27464
rect 14967 27424 15200 27452
rect 14967 27421 14979 27424
rect 14921 27415 14979 27421
rect 15194 27412 15200 27424
rect 15252 27412 15258 27464
rect 17221 27455 17279 27461
rect 17221 27421 17233 27455
rect 17267 27452 17279 27455
rect 18230 27452 18236 27464
rect 17267 27424 18236 27452
rect 17267 27421 17279 27424
rect 17221 27415 17279 27421
rect 18230 27412 18236 27424
rect 18288 27412 18294 27464
rect 19444 27452 19472 27548
rect 19797 27523 19855 27529
rect 19797 27489 19809 27523
rect 19843 27520 19855 27523
rect 20438 27520 20444 27532
rect 19843 27492 20444 27520
rect 19843 27489 19855 27492
rect 19797 27483 19855 27489
rect 20438 27480 20444 27492
rect 20496 27480 20502 27532
rect 21729 27523 21787 27529
rect 21729 27489 21741 27523
rect 21775 27520 21787 27523
rect 22002 27520 22008 27532
rect 21775 27492 22008 27520
rect 21775 27489 21787 27492
rect 21729 27483 21787 27489
rect 22002 27480 22008 27492
rect 22060 27480 22066 27532
rect 19705 27455 19763 27461
rect 19705 27452 19717 27455
rect 19444 27424 19717 27452
rect 19705 27421 19717 27424
rect 19751 27421 19763 27455
rect 19705 27415 19763 27421
rect 20898 27412 20904 27464
rect 20956 27452 20962 27464
rect 22480 27461 22508 27560
rect 24394 27548 24400 27600
rect 24452 27588 24458 27600
rect 30101 27591 30159 27597
rect 24452 27560 26004 27588
rect 24452 27548 24458 27560
rect 23198 27480 23204 27532
rect 23256 27520 23262 27532
rect 25976 27529 26004 27560
rect 30101 27557 30113 27591
rect 30147 27588 30159 27591
rect 31018 27588 31024 27600
rect 30147 27560 31024 27588
rect 30147 27557 30159 27560
rect 30101 27551 30159 27557
rect 31018 27548 31024 27560
rect 31076 27548 31082 27600
rect 31665 27591 31723 27597
rect 31665 27557 31677 27591
rect 31711 27588 31723 27591
rect 32398 27588 32404 27600
rect 31711 27560 32404 27588
rect 31711 27557 31723 27560
rect 31665 27551 31723 27557
rect 32398 27548 32404 27560
rect 32456 27548 32462 27600
rect 36446 27548 36452 27600
rect 36504 27588 36510 27600
rect 40310 27588 40316 27600
rect 36504 27560 39988 27588
rect 40271 27560 40316 27588
rect 36504 27548 36510 27560
rect 24581 27523 24639 27529
rect 24581 27520 24593 27523
rect 23256 27492 24593 27520
rect 23256 27480 23262 27492
rect 24581 27489 24593 27492
rect 24627 27489 24639 27523
rect 25961 27523 26019 27529
rect 24581 27483 24639 27489
rect 24688 27492 24900 27520
rect 21637 27455 21695 27461
rect 21637 27452 21649 27455
rect 20956 27424 21649 27452
rect 20956 27412 20962 27424
rect 21637 27421 21649 27424
rect 21683 27421 21695 27455
rect 21637 27415 21695 27421
rect 22465 27455 22523 27461
rect 22465 27421 22477 27455
rect 22511 27421 22523 27455
rect 22465 27415 22523 27421
rect 22646 27412 22652 27464
rect 22704 27452 22710 27464
rect 24688 27452 24716 27492
rect 24762 27461 24768 27464
rect 22704 27424 24716 27452
rect 24751 27455 24768 27461
rect 22704 27412 22710 27424
rect 24751 27421 24763 27455
rect 24751 27415 24768 27421
rect 24762 27412 24768 27415
rect 24820 27412 24826 27464
rect 24872 27452 24900 27492
rect 25961 27489 25973 27523
rect 26007 27489 26019 27523
rect 29362 27520 29368 27532
rect 25961 27483 26019 27489
rect 28368 27492 29368 27520
rect 28368 27461 28396 27492
rect 29362 27480 29368 27492
rect 29420 27520 29426 27532
rect 29641 27523 29699 27529
rect 29641 27520 29653 27523
rect 29420 27492 29653 27520
rect 29420 27480 29426 27492
rect 29641 27489 29653 27492
rect 29687 27489 29699 27523
rect 31202 27520 31208 27532
rect 31163 27492 31208 27520
rect 29641 27483 29699 27489
rect 31202 27480 31208 27492
rect 31260 27480 31266 27532
rect 39206 27480 39212 27532
rect 39264 27520 39270 27532
rect 39960 27520 39988 27560
rect 40310 27548 40316 27560
rect 40368 27548 40374 27600
rect 45002 27588 45008 27600
rect 44963 27560 45008 27588
rect 45002 27548 45008 27560
rect 45060 27548 45066 27600
rect 45186 27588 45192 27600
rect 45147 27560 45192 27588
rect 45186 27548 45192 27560
rect 45244 27548 45250 27600
rect 41141 27523 41199 27529
rect 41141 27520 41153 27523
rect 39264 27492 39896 27520
rect 39960 27492 41153 27520
rect 39264 27480 39270 27492
rect 28077 27455 28135 27461
rect 28077 27452 28089 27455
rect 24872 27424 28089 27452
rect 28077 27421 28089 27424
rect 28123 27421 28135 27455
rect 28077 27415 28135 27421
rect 28353 27455 28411 27461
rect 28353 27421 28365 27455
rect 28399 27421 28411 27455
rect 28810 27452 28816 27464
rect 28771 27424 28816 27452
rect 28353 27415 28411 27421
rect 28810 27412 28816 27424
rect 28868 27412 28874 27464
rect 28997 27455 29055 27461
rect 28997 27421 29009 27455
rect 29043 27452 29055 27455
rect 29733 27455 29791 27461
rect 29733 27452 29745 27455
rect 29043 27424 29745 27452
rect 29043 27421 29055 27424
rect 28997 27415 29055 27421
rect 29733 27421 29745 27424
rect 29779 27421 29791 27455
rect 31294 27452 31300 27464
rect 31255 27424 31300 27452
rect 29733 27415 29791 27421
rect 12253 27387 12311 27393
rect 12253 27384 12265 27387
rect 11532 27356 12265 27384
rect 12253 27353 12265 27356
rect 12299 27384 12311 27387
rect 17034 27384 17040 27396
rect 12299 27356 17040 27384
rect 12299 27353 12311 27356
rect 12253 27347 12311 27353
rect 17034 27344 17040 27356
rect 17092 27344 17098 27396
rect 17310 27344 17316 27396
rect 17368 27384 17374 27396
rect 17466 27387 17524 27393
rect 17466 27384 17478 27387
rect 17368 27356 17478 27384
rect 17368 27344 17374 27356
rect 17466 27353 17478 27356
rect 17512 27353 17524 27387
rect 19334 27384 19340 27396
rect 19295 27356 19340 27384
rect 17466 27347 17524 27353
rect 19334 27344 19340 27356
rect 19392 27344 19398 27396
rect 19429 27387 19487 27393
rect 19429 27353 19441 27387
rect 19475 27384 19487 27387
rect 19518 27384 19524 27396
rect 19475 27356 19524 27384
rect 19475 27353 19487 27356
rect 19429 27347 19487 27353
rect 19518 27344 19524 27356
rect 19576 27384 19582 27396
rect 20162 27384 20168 27396
rect 19576 27356 20168 27384
rect 19576 27344 19582 27356
rect 20162 27344 20168 27356
rect 20220 27344 20226 27396
rect 20441 27387 20499 27393
rect 20441 27353 20453 27387
rect 20487 27384 20499 27387
rect 20806 27384 20812 27396
rect 20487 27356 20812 27384
rect 20487 27353 20499 27356
rect 20441 27347 20499 27353
rect 20806 27344 20812 27356
rect 20864 27344 20870 27396
rect 26234 27393 26240 27396
rect 22557 27387 22615 27393
rect 22557 27353 22569 27387
rect 22603 27384 22615 27387
rect 22603 27356 26188 27384
rect 22603 27353 22615 27356
rect 22557 27347 22615 27353
rect 4617 27319 4675 27325
rect 4617 27285 4629 27319
rect 4663 27316 4675 27319
rect 4706 27316 4712 27328
rect 4663 27288 4712 27316
rect 4663 27285 4675 27288
rect 4617 27279 4675 27285
rect 4706 27276 4712 27288
rect 4764 27276 4770 27328
rect 6914 27316 6920 27328
rect 6875 27288 6920 27316
rect 6914 27276 6920 27288
rect 6972 27276 6978 27328
rect 9033 27319 9091 27325
rect 9033 27285 9045 27319
rect 9079 27316 9091 27319
rect 9306 27316 9312 27328
rect 9079 27288 9312 27316
rect 9079 27285 9091 27288
rect 9033 27279 9091 27285
rect 9306 27276 9312 27288
rect 9364 27276 9370 27328
rect 10226 27316 10232 27328
rect 10187 27288 10232 27316
rect 10226 27276 10232 27288
rect 10284 27276 10290 27328
rect 11057 27319 11115 27325
rect 11057 27285 11069 27319
rect 11103 27316 11115 27319
rect 11238 27316 11244 27328
rect 11103 27288 11244 27316
rect 11103 27285 11115 27288
rect 11057 27279 11115 27285
rect 11238 27276 11244 27288
rect 11296 27276 11302 27328
rect 12897 27319 12955 27325
rect 12897 27285 12909 27319
rect 12943 27316 12955 27319
rect 12986 27316 12992 27328
rect 12943 27288 12992 27316
rect 12943 27285 12955 27288
rect 12897 27279 12955 27285
rect 12986 27276 12992 27288
rect 13044 27276 13050 27328
rect 15562 27316 15568 27328
rect 15475 27288 15568 27316
rect 15562 27276 15568 27288
rect 15620 27316 15626 27328
rect 18414 27316 18420 27328
rect 15620 27288 18420 27316
rect 15620 27276 15626 27288
rect 18414 27276 18420 27288
rect 18472 27276 18478 27328
rect 19978 27316 19984 27328
rect 19939 27288 19984 27316
rect 19978 27276 19984 27288
rect 20036 27276 20042 27328
rect 22005 27319 22063 27325
rect 22005 27285 22017 27319
rect 22051 27316 22063 27319
rect 23290 27316 23296 27328
rect 22051 27288 23296 27316
rect 22051 27285 22063 27288
rect 22005 27279 22063 27285
rect 23290 27276 23296 27288
rect 23348 27276 23354 27328
rect 23385 27319 23443 27325
rect 23385 27285 23397 27319
rect 23431 27316 23443 27319
rect 23658 27316 23664 27328
rect 23431 27288 23664 27316
rect 23431 27285 23443 27288
rect 23385 27279 23443 27285
rect 23658 27276 23664 27288
rect 23716 27276 23722 27328
rect 25041 27319 25099 27325
rect 25041 27285 25053 27319
rect 25087 27316 25099 27319
rect 25406 27316 25412 27328
rect 25087 27288 25412 27316
rect 25087 27285 25099 27288
rect 25041 27279 25099 27285
rect 25406 27276 25412 27288
rect 25464 27276 25470 27328
rect 26160 27316 26188 27356
rect 26228 27347 26240 27393
rect 26292 27384 26298 27396
rect 28261 27387 28319 27393
rect 28261 27384 28273 27387
rect 26292 27356 26328 27384
rect 27172 27356 28273 27384
rect 26234 27344 26240 27347
rect 26292 27344 26298 27356
rect 27172 27316 27200 27356
rect 28261 27353 28273 27356
rect 28307 27384 28319 27387
rect 29012 27384 29040 27415
rect 31294 27412 31300 27424
rect 31352 27412 31358 27464
rect 36633 27455 36691 27461
rect 36633 27421 36645 27455
rect 36679 27421 36691 27455
rect 36633 27415 36691 27421
rect 36817 27455 36875 27461
rect 36817 27421 36829 27455
rect 36863 27452 36875 27455
rect 37458 27452 37464 27464
rect 36863 27424 37464 27452
rect 36863 27421 36875 27424
rect 36817 27415 36875 27421
rect 28307 27356 29040 27384
rect 28307 27353 28319 27356
rect 28261 27347 28319 27353
rect 30282 27344 30288 27396
rect 30340 27384 30346 27396
rect 36648 27384 36676 27415
rect 37458 27412 37464 27424
rect 37516 27412 37522 27464
rect 39117 27455 39175 27461
rect 39117 27452 39129 27455
rect 38672 27424 39129 27452
rect 37277 27387 37335 27393
rect 37277 27384 37289 27387
rect 30340 27356 37289 27384
rect 30340 27344 30346 27356
rect 37277 27353 37289 27356
rect 37323 27353 37335 27387
rect 37277 27347 37335 27353
rect 38672 27328 38700 27424
rect 39117 27421 39129 27424
rect 39163 27421 39175 27455
rect 39298 27452 39304 27464
rect 39259 27424 39304 27452
rect 39117 27415 39175 27421
rect 39298 27412 39304 27424
rect 39356 27412 39362 27464
rect 39868 27461 39896 27492
rect 41141 27489 41153 27492
rect 41187 27520 41199 27523
rect 41506 27520 41512 27532
rect 41187 27492 41512 27520
rect 41187 27489 41199 27492
rect 41141 27483 41199 27489
rect 41506 27480 41512 27492
rect 41564 27480 41570 27532
rect 43438 27520 43444 27532
rect 43399 27492 43444 27520
rect 43438 27480 43444 27492
rect 43496 27480 43502 27532
rect 45462 27520 45468 27532
rect 45423 27492 45468 27520
rect 45462 27480 45468 27492
rect 45520 27480 45526 27532
rect 39853 27455 39911 27461
rect 39853 27421 39865 27455
rect 39899 27421 39911 27455
rect 39853 27415 39911 27421
rect 40129 27455 40187 27461
rect 40129 27421 40141 27455
rect 40175 27421 40187 27455
rect 41414 27452 41420 27464
rect 41375 27424 41420 27452
rect 40129 27415 40187 27421
rect 39758 27344 39764 27396
rect 39816 27384 39822 27396
rect 40144 27384 40172 27415
rect 41414 27412 41420 27424
rect 41472 27412 41478 27464
rect 42245 27455 42303 27461
rect 42245 27452 42257 27455
rect 41800 27424 42257 27452
rect 39816 27356 40172 27384
rect 39816 27344 39822 27356
rect 27338 27316 27344 27328
rect 26160 27288 27200 27316
rect 27299 27288 27344 27316
rect 27338 27276 27344 27288
rect 27396 27276 27402 27328
rect 28994 27316 29000 27328
rect 28907 27288 29000 27316
rect 28994 27276 29000 27288
rect 29052 27316 29058 27328
rect 35526 27316 35532 27328
rect 29052 27288 35532 27316
rect 29052 27276 29058 27288
rect 35526 27276 35532 27288
rect 35584 27276 35590 27328
rect 36722 27316 36728 27328
rect 36683 27288 36728 27316
rect 36722 27276 36728 27288
rect 36780 27276 36786 27328
rect 38654 27316 38660 27328
rect 38615 27288 38660 27316
rect 38654 27276 38660 27288
rect 38712 27276 38718 27328
rect 39209 27319 39267 27325
rect 39209 27285 39221 27319
rect 39255 27316 39267 27319
rect 39574 27316 39580 27328
rect 39255 27288 39580 27316
rect 39255 27285 39267 27288
rect 39209 27279 39267 27285
rect 39574 27276 39580 27288
rect 39632 27276 39638 27328
rect 39945 27319 40003 27325
rect 39945 27285 39957 27319
rect 39991 27316 40003 27319
rect 40218 27316 40224 27328
rect 39991 27288 40224 27316
rect 39991 27285 40003 27288
rect 39945 27279 40003 27285
rect 40218 27276 40224 27288
rect 40276 27276 40282 27328
rect 41322 27316 41328 27328
rect 41283 27288 41328 27316
rect 41322 27276 41328 27288
rect 41380 27276 41386 27328
rect 41800 27325 41828 27424
rect 42245 27421 42257 27424
rect 42291 27421 42303 27455
rect 42245 27415 42303 27421
rect 43622 27412 43628 27464
rect 43680 27452 43686 27464
rect 43717 27455 43775 27461
rect 43717 27452 43729 27455
rect 43680 27424 43729 27452
rect 43680 27412 43686 27424
rect 43717 27421 43729 27424
rect 43763 27421 43775 27455
rect 43717 27415 43775 27421
rect 41785 27319 41843 27325
rect 41785 27285 41797 27319
rect 41831 27285 41843 27319
rect 42426 27316 42432 27328
rect 42387 27288 42432 27316
rect 41785 27279 41843 27285
rect 42426 27276 42432 27288
rect 42484 27276 42490 27328
rect 43898 27276 43904 27328
rect 43956 27316 43962 27328
rect 44453 27319 44511 27325
rect 44453 27316 44465 27319
rect 43956 27288 44465 27316
rect 43956 27276 43962 27288
rect 44453 27285 44465 27288
rect 44499 27285 44511 27319
rect 44453 27279 44511 27285
rect 1104 27226 68816 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 68816 27226
rect 1104 27152 68816 27174
rect 7742 27112 7748 27124
rect 7703 27084 7748 27112
rect 7742 27072 7748 27084
rect 7800 27072 7806 27124
rect 8754 27112 8760 27124
rect 8715 27084 8760 27112
rect 8754 27072 8760 27084
rect 8812 27072 8818 27124
rect 12621 27115 12679 27121
rect 12621 27081 12633 27115
rect 12667 27081 12679 27115
rect 12621 27075 12679 27081
rect 13633 27115 13691 27121
rect 13633 27081 13645 27115
rect 13679 27112 13691 27115
rect 14090 27112 14096 27124
rect 13679 27084 14096 27112
rect 13679 27081 13691 27084
rect 13633 27075 13691 27081
rect 4614 27044 4620 27056
rect 4448 27016 4620 27044
rect 4448 26985 4476 27016
rect 4614 27004 4620 27016
rect 4672 27044 4678 27056
rect 6632 27047 6690 27053
rect 4672 27016 5120 27044
rect 4672 27004 4678 27016
rect 5092 26988 5120 27016
rect 6632 27013 6644 27047
rect 6678 27044 6690 27047
rect 6914 27044 6920 27056
rect 6678 27016 6920 27044
rect 6678 27013 6690 27016
rect 6632 27007 6690 27013
rect 6914 27004 6920 27016
rect 6972 27004 6978 27056
rect 9674 27044 9680 27056
rect 9324 27016 9680 27044
rect 4706 26985 4712 26988
rect 4433 26979 4491 26985
rect 4433 26945 4445 26979
rect 4479 26945 4491 26979
rect 4700 26976 4712 26985
rect 4667 26948 4712 26976
rect 4433 26939 4491 26945
rect 4700 26939 4712 26948
rect 4706 26936 4712 26939
rect 4764 26936 4770 26988
rect 5074 26936 5080 26988
rect 5132 26976 5138 26988
rect 8294 26976 8300 26988
rect 5132 26948 6408 26976
rect 8255 26948 8300 26976
rect 5132 26936 5138 26948
rect 6380 26920 6408 26948
rect 8294 26936 8300 26948
rect 8352 26936 8358 26988
rect 6362 26908 6368 26920
rect 6323 26880 6368 26908
rect 6362 26868 6368 26880
rect 6420 26868 6426 26920
rect 9324 26917 9352 27016
rect 9674 27004 9680 27016
rect 9732 27004 9738 27056
rect 10226 27004 10232 27056
rect 10284 27044 10290 27056
rect 10284 27016 12572 27044
rect 10284 27004 10290 27016
rect 9401 26979 9459 26985
rect 9401 26945 9413 26979
rect 9447 26976 9459 26979
rect 9582 26976 9588 26988
rect 9447 26948 9588 26976
rect 9447 26945 9459 26948
rect 9401 26939 9459 26945
rect 9582 26936 9588 26948
rect 9640 26936 9646 26988
rect 12360 26985 12388 27016
rect 10597 26979 10655 26985
rect 10597 26976 10609 26979
rect 9692 26948 10609 26976
rect 9309 26911 9367 26917
rect 9309 26877 9321 26911
rect 9355 26877 9367 26911
rect 9309 26871 9367 26877
rect 9692 26840 9720 26948
rect 10597 26945 10609 26948
rect 10643 26945 10655 26979
rect 10597 26939 10655 26945
rect 12345 26979 12403 26985
rect 12345 26945 12357 26979
rect 12391 26976 12403 26979
rect 12391 26948 12425 26976
rect 12391 26945 12403 26948
rect 12345 26939 12403 26945
rect 10686 26908 10692 26920
rect 10647 26880 10692 26908
rect 10686 26868 10692 26880
rect 10744 26868 10750 26920
rect 10873 26911 10931 26917
rect 10873 26877 10885 26911
rect 10919 26908 10931 26911
rect 11977 26911 12035 26917
rect 10919 26880 11652 26908
rect 10919 26877 10931 26880
rect 10873 26871 10931 26877
rect 9140 26812 9720 26840
rect 9140 26784 9168 26812
rect 5166 26732 5172 26784
rect 5224 26772 5230 26784
rect 5813 26775 5871 26781
rect 5813 26772 5825 26775
rect 5224 26744 5825 26772
rect 5224 26732 5230 26744
rect 5813 26741 5825 26744
rect 5859 26741 5871 26775
rect 5813 26735 5871 26741
rect 6546 26732 6552 26784
rect 6604 26772 6610 26784
rect 8389 26775 8447 26781
rect 8389 26772 8401 26775
rect 6604 26744 8401 26772
rect 6604 26732 6610 26744
rect 8389 26741 8401 26744
rect 8435 26772 8447 26775
rect 9122 26772 9128 26784
rect 8435 26744 9128 26772
rect 8435 26741 8447 26744
rect 8389 26735 8447 26741
rect 9122 26732 9128 26744
rect 9180 26732 9186 26784
rect 9766 26772 9772 26784
rect 9727 26744 9772 26772
rect 9766 26732 9772 26744
rect 9824 26732 9830 26784
rect 10226 26772 10232 26784
rect 10187 26744 10232 26772
rect 10226 26732 10232 26744
rect 10284 26732 10290 26784
rect 11624 26772 11652 26880
rect 11977 26877 11989 26911
rect 12023 26877 12035 26911
rect 11977 26871 12035 26877
rect 12069 26911 12127 26917
rect 12069 26877 12081 26911
rect 12115 26908 12127 26911
rect 12250 26908 12256 26920
rect 12115 26880 12256 26908
rect 12115 26877 12127 26880
rect 12069 26871 12127 26877
rect 11992 26840 12020 26871
rect 12250 26868 12256 26880
rect 12308 26868 12314 26920
rect 12437 26911 12495 26917
rect 12437 26877 12449 26911
rect 12483 26877 12495 26911
rect 12544 26908 12572 27016
rect 12636 26976 12664 27075
rect 14090 27072 14096 27084
rect 14148 27072 14154 27124
rect 17310 27112 17316 27124
rect 17271 27084 17316 27112
rect 17310 27072 17316 27084
rect 17368 27072 17374 27124
rect 19429 27115 19487 27121
rect 19429 27081 19441 27115
rect 19475 27112 19487 27115
rect 20346 27112 20352 27124
rect 19475 27084 20352 27112
rect 19475 27081 19487 27084
rect 19429 27075 19487 27081
rect 20346 27072 20352 27084
rect 20404 27072 20410 27124
rect 23198 27112 23204 27124
rect 23159 27084 23204 27112
rect 23198 27072 23204 27084
rect 23256 27072 23262 27124
rect 24210 27112 24216 27124
rect 24171 27084 24216 27112
rect 24210 27072 24216 27084
rect 24268 27072 24274 27124
rect 25409 27115 25467 27121
rect 25409 27081 25421 27115
rect 25455 27112 25467 27115
rect 25774 27112 25780 27124
rect 25455 27084 25780 27112
rect 25455 27081 25467 27084
rect 25409 27075 25467 27081
rect 25774 27072 25780 27084
rect 25832 27072 25838 27124
rect 27433 27115 27491 27121
rect 27433 27081 27445 27115
rect 27479 27112 27491 27115
rect 27522 27112 27528 27124
rect 27479 27084 27528 27112
rect 27479 27081 27491 27084
rect 27433 27075 27491 27081
rect 27522 27072 27528 27084
rect 27580 27072 27586 27124
rect 36265 27115 36323 27121
rect 36265 27081 36277 27115
rect 36311 27081 36323 27115
rect 36265 27075 36323 27081
rect 39117 27115 39175 27121
rect 39117 27081 39129 27115
rect 39163 27112 39175 27115
rect 40218 27112 40224 27124
rect 39163 27084 40224 27112
rect 39163 27081 39175 27084
rect 39117 27075 39175 27081
rect 12802 27004 12808 27056
rect 12860 27044 12866 27056
rect 12860 27016 13400 27044
rect 12860 27004 12866 27016
rect 13081 26979 13139 26985
rect 13081 26976 13093 26979
rect 12636 26948 13093 26976
rect 13081 26945 13093 26948
rect 13127 26945 13139 26979
rect 13081 26939 13139 26945
rect 13170 26936 13176 26988
rect 13228 26976 13234 26988
rect 13372 26985 13400 27016
rect 17034 27004 17040 27056
rect 17092 27044 17098 27056
rect 17092 27016 19104 27044
rect 17092 27004 17098 27016
rect 13357 26979 13415 26985
rect 13228 26948 13273 26976
rect 13228 26936 13234 26948
rect 13357 26945 13369 26979
rect 13403 26945 13415 26979
rect 13357 26939 13415 26945
rect 13449 26979 13507 26985
rect 13449 26945 13461 26979
rect 13495 26945 13507 26979
rect 17126 26976 17132 26988
rect 17087 26948 17132 26976
rect 13449 26939 13507 26945
rect 13464 26908 13492 26939
rect 17126 26936 17132 26948
rect 17184 26936 17190 26988
rect 18322 26985 18328 26988
rect 18316 26939 18328 26985
rect 18380 26976 18386 26988
rect 18380 26948 18416 26976
rect 18322 26936 18328 26939
rect 18380 26936 18386 26948
rect 12544 26880 13492 26908
rect 12437 26871 12495 26877
rect 12342 26840 12348 26852
rect 11992 26812 12348 26840
rect 12342 26800 12348 26812
rect 12400 26800 12406 26852
rect 12452 26840 12480 26871
rect 17862 26868 17868 26920
rect 17920 26908 17926 26920
rect 18049 26911 18107 26917
rect 18049 26908 18061 26911
rect 17920 26880 18061 26908
rect 17920 26868 17926 26880
rect 18049 26877 18061 26880
rect 18095 26877 18107 26911
rect 18049 26871 18107 26877
rect 12802 26840 12808 26852
rect 12452 26812 12808 26840
rect 12802 26800 12808 26812
rect 12860 26800 12866 26852
rect 19076 26840 19104 27016
rect 19978 27004 19984 27056
rect 20036 27044 20042 27056
rect 29546 27044 29552 27056
rect 20036 27016 29552 27044
rect 20036 27004 20042 27016
rect 29546 27004 29552 27016
rect 29604 27004 29610 27056
rect 30926 27004 30932 27056
rect 30984 27044 30990 27056
rect 31205 27047 31263 27053
rect 31205 27044 31217 27047
rect 30984 27016 31217 27044
rect 30984 27004 30990 27016
rect 31205 27013 31217 27016
rect 31251 27013 31263 27047
rect 36280 27044 36308 27075
rect 40218 27072 40224 27084
rect 40276 27072 40282 27124
rect 40494 27072 40500 27124
rect 40552 27112 40558 27124
rect 40681 27115 40739 27121
rect 40681 27112 40693 27115
rect 40552 27084 40693 27112
rect 40552 27072 40558 27084
rect 40681 27081 40693 27084
rect 40727 27081 40739 27115
rect 40681 27075 40739 27081
rect 45186 27072 45192 27124
rect 45244 27112 45250 27124
rect 45373 27115 45431 27121
rect 45373 27112 45385 27115
rect 45244 27084 45385 27112
rect 45244 27072 45250 27084
rect 45373 27081 45385 27084
rect 45419 27081 45431 27115
rect 45373 27075 45431 27081
rect 45830 27072 45836 27124
rect 45888 27112 45894 27124
rect 45925 27115 45983 27121
rect 45925 27112 45937 27115
rect 45888 27084 45937 27112
rect 45888 27072 45894 27084
rect 45925 27081 45937 27084
rect 45971 27081 45983 27115
rect 45925 27075 45983 27081
rect 38746 27044 38752 27056
rect 36280 27016 38752 27044
rect 31205 27007 31263 27013
rect 38746 27004 38752 27016
rect 38804 27044 38810 27056
rect 39853 27047 39911 27053
rect 38804 27016 38976 27044
rect 38804 27004 38810 27016
rect 20257 26979 20315 26985
rect 20257 26945 20269 26979
rect 20303 26976 20315 26979
rect 20622 26976 20628 26988
rect 20303 26948 20628 26976
rect 20303 26945 20315 26948
rect 20257 26939 20315 26945
rect 20622 26936 20628 26948
rect 20680 26976 20686 26988
rect 21085 26979 21143 26985
rect 21085 26976 21097 26979
rect 20680 26948 21097 26976
rect 20680 26936 20686 26948
rect 21085 26945 21097 26948
rect 21131 26945 21143 26979
rect 21085 26939 21143 26945
rect 22833 26979 22891 26985
rect 22833 26945 22845 26979
rect 22879 26976 22891 26979
rect 23658 26976 23664 26988
rect 22879 26948 23664 26976
rect 22879 26945 22891 26948
rect 22833 26939 22891 26945
rect 23658 26936 23664 26948
rect 23716 26936 23722 26988
rect 24305 26979 24363 26985
rect 24305 26945 24317 26979
rect 24351 26945 24363 26979
rect 24305 26939 24363 26945
rect 25041 26979 25099 26985
rect 25041 26945 25053 26979
rect 25087 26976 25099 26979
rect 25130 26976 25136 26988
rect 25087 26948 25136 26976
rect 25087 26945 25099 26948
rect 25041 26939 25099 26945
rect 20533 26911 20591 26917
rect 20533 26877 20545 26911
rect 20579 26908 20591 26911
rect 20714 26908 20720 26920
rect 20579 26880 20720 26908
rect 20579 26877 20591 26880
rect 20533 26871 20591 26877
rect 20714 26868 20720 26880
rect 20772 26868 20778 26920
rect 22925 26911 22983 26917
rect 22925 26877 22937 26911
rect 22971 26908 22983 26911
rect 23106 26908 23112 26920
rect 22971 26880 23112 26908
rect 22971 26877 22983 26880
rect 22925 26871 22983 26877
rect 23106 26868 23112 26880
rect 23164 26868 23170 26920
rect 22738 26840 22744 26852
rect 19076 26812 22744 26840
rect 22738 26800 22744 26812
rect 22796 26800 22802 26852
rect 24320 26840 24348 26939
rect 25130 26936 25136 26948
rect 25188 26936 25194 26988
rect 27430 26936 27436 26988
rect 27488 26976 27494 26988
rect 27525 26979 27583 26985
rect 27525 26976 27537 26979
rect 27488 26948 27537 26976
rect 27488 26936 27494 26948
rect 27525 26945 27537 26948
rect 27571 26945 27583 26979
rect 27525 26939 27583 26945
rect 30745 26979 30803 26985
rect 30745 26945 30757 26979
rect 30791 26976 30803 26979
rect 31389 26979 31447 26985
rect 31389 26976 31401 26979
rect 30791 26948 31401 26976
rect 30791 26945 30803 26948
rect 30745 26939 30803 26945
rect 31389 26945 31401 26948
rect 31435 26976 31447 26979
rect 32122 26976 32128 26988
rect 31435 26948 31754 26976
rect 32083 26948 32128 26976
rect 31435 26945 31447 26948
rect 31389 26939 31447 26945
rect 24946 26908 24952 26920
rect 24907 26880 24952 26908
rect 24946 26868 24952 26880
rect 25004 26868 25010 26920
rect 31726 26908 31754 26948
rect 32122 26936 32128 26948
rect 32180 26936 32186 26988
rect 34514 26976 34520 26988
rect 34475 26948 34520 26976
rect 34514 26936 34520 26948
rect 34572 26936 34578 26988
rect 35618 26936 35624 26988
rect 35676 26976 35682 26988
rect 35897 26979 35955 26985
rect 35897 26976 35909 26979
rect 35676 26948 35909 26976
rect 35676 26936 35682 26948
rect 35897 26945 35909 26948
rect 35943 26945 35955 26979
rect 38838 26976 38844 26988
rect 38799 26948 38844 26976
rect 35897 26939 35955 26945
rect 38838 26936 38844 26948
rect 38896 26936 38902 26988
rect 38948 26985 38976 27016
rect 39853 27013 39865 27047
rect 39899 27044 39911 27047
rect 40770 27044 40776 27056
rect 39899 27016 40776 27044
rect 39899 27013 39911 27016
rect 39853 27007 39911 27013
rect 40770 27004 40776 27016
rect 40828 27004 40834 27056
rect 43898 27044 43904 27056
rect 43859 27016 43904 27044
rect 43898 27004 43904 27016
rect 43956 27004 43962 27056
rect 38933 26979 38991 26985
rect 38933 26945 38945 26979
rect 38979 26945 38991 26979
rect 39574 26976 39580 26988
rect 39535 26948 39580 26976
rect 38933 26939 38991 26945
rect 39574 26936 39580 26948
rect 39632 26936 39638 26988
rect 39670 26979 39728 26985
rect 39670 26945 39682 26979
rect 39716 26976 39728 26979
rect 39758 26976 39764 26988
rect 39716 26948 39764 26976
rect 39716 26945 39728 26948
rect 39670 26939 39728 26945
rect 34422 26908 34428 26920
rect 31726 26880 34428 26908
rect 34422 26868 34428 26880
rect 34480 26868 34486 26920
rect 35989 26911 36047 26917
rect 35989 26877 36001 26911
rect 36035 26908 36047 26911
rect 36078 26908 36084 26920
rect 36035 26880 36084 26908
rect 36035 26877 36047 26880
rect 35989 26871 36047 26877
rect 36078 26868 36084 26880
rect 36136 26868 36142 26920
rect 38194 26868 38200 26920
rect 38252 26908 38258 26920
rect 39684 26908 39712 26939
rect 39758 26936 39764 26948
rect 39816 26936 39822 26988
rect 39945 26979 40003 26985
rect 39945 26976 39957 26979
rect 39868 26948 39957 26976
rect 39868 26920 39896 26948
rect 39945 26945 39957 26948
rect 39991 26945 40003 26979
rect 39945 26939 40003 26945
rect 40042 26979 40100 26985
rect 40042 26945 40054 26979
rect 40088 26945 40100 26979
rect 40865 26979 40923 26985
rect 40865 26976 40877 26979
rect 40042 26939 40100 26945
rect 40236 26948 40877 26976
rect 38252 26880 39712 26908
rect 38252 26868 38258 26880
rect 39850 26868 39856 26920
rect 39908 26868 39914 26920
rect 40052 26852 40080 26939
rect 25866 26840 25872 26852
rect 24320 26812 25872 26840
rect 25866 26800 25872 26812
rect 25924 26800 25930 26852
rect 36722 26800 36728 26852
rect 36780 26840 36786 26852
rect 40034 26840 40040 26852
rect 36780 26812 40040 26840
rect 36780 26800 36786 26812
rect 40034 26800 40040 26812
rect 40092 26800 40098 26852
rect 40236 26849 40264 26948
rect 40865 26945 40877 26948
rect 40911 26945 40923 26979
rect 41046 26976 41052 26988
rect 41007 26948 41052 26976
rect 40865 26939 40923 26945
rect 41046 26936 41052 26948
rect 41104 26936 41110 26988
rect 41141 26979 41199 26985
rect 41141 26945 41153 26979
rect 41187 26945 41199 26979
rect 43622 26976 43628 26988
rect 43583 26948 43628 26976
rect 41141 26939 41199 26945
rect 41156 26908 41184 26939
rect 43622 26936 43628 26948
rect 43680 26936 43686 26988
rect 45002 26936 45008 26988
rect 45060 26936 45066 26988
rect 45278 26936 45284 26988
rect 45336 26976 45342 26988
rect 45833 26979 45891 26985
rect 45833 26976 45845 26979
rect 45336 26948 45845 26976
rect 45336 26936 45342 26948
rect 45833 26945 45845 26948
rect 45879 26945 45891 26979
rect 45833 26939 45891 26945
rect 41064 26880 41184 26908
rect 40221 26843 40279 26849
rect 40221 26809 40233 26843
rect 40267 26809 40279 26843
rect 40221 26803 40279 26809
rect 13814 26772 13820 26784
rect 11624 26744 13820 26772
rect 13814 26732 13820 26744
rect 13872 26772 13878 26784
rect 13998 26772 14004 26784
rect 13872 26744 14004 26772
rect 13872 26732 13878 26744
rect 13998 26732 14004 26744
rect 14056 26732 14062 26784
rect 14274 26772 14280 26784
rect 14235 26744 14280 26772
rect 14274 26732 14280 26744
rect 14332 26772 14338 26784
rect 14829 26775 14887 26781
rect 14829 26772 14841 26775
rect 14332 26744 14841 26772
rect 14332 26732 14338 26744
rect 14829 26741 14841 26744
rect 14875 26741 14887 26775
rect 15562 26772 15568 26784
rect 15523 26744 15568 26772
rect 14829 26735 14887 26741
rect 15562 26732 15568 26744
rect 15620 26732 15626 26784
rect 19889 26775 19947 26781
rect 19889 26741 19901 26775
rect 19935 26772 19947 26775
rect 19978 26772 19984 26784
rect 19935 26744 19984 26772
rect 19935 26741 19947 26744
rect 19889 26735 19947 26741
rect 19978 26732 19984 26744
rect 20036 26732 20042 26784
rect 32309 26775 32367 26781
rect 32309 26741 32321 26775
rect 32355 26772 32367 26775
rect 33226 26772 33232 26784
rect 32355 26744 33232 26772
rect 32355 26741 32367 26744
rect 32309 26735 32367 26741
rect 33226 26732 33232 26744
rect 33284 26732 33290 26784
rect 34701 26775 34759 26781
rect 34701 26741 34713 26775
rect 34747 26772 34759 26775
rect 34790 26772 34796 26784
rect 34747 26744 34796 26772
rect 34747 26741 34759 26744
rect 34701 26735 34759 26741
rect 34790 26732 34796 26744
rect 34848 26732 34854 26784
rect 35253 26775 35311 26781
rect 35253 26741 35265 26775
rect 35299 26772 35311 26775
rect 35618 26772 35624 26784
rect 35299 26744 35624 26772
rect 35299 26741 35311 26744
rect 35253 26735 35311 26741
rect 35618 26732 35624 26744
rect 35676 26732 35682 26784
rect 39206 26732 39212 26784
rect 39264 26772 39270 26784
rect 41064 26772 41092 26880
rect 39264 26744 41092 26772
rect 39264 26732 39270 26744
rect 1104 26682 68816 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 65654 26682
rect 65706 26630 65718 26682
rect 65770 26630 65782 26682
rect 65834 26630 65846 26682
rect 65898 26630 65910 26682
rect 65962 26630 68816 26682
rect 1104 26608 68816 26630
rect 4798 26568 4804 26580
rect 4759 26540 4804 26568
rect 4798 26528 4804 26540
rect 4856 26528 4862 26580
rect 5994 26568 6000 26580
rect 5955 26540 6000 26568
rect 5994 26528 6000 26540
rect 6052 26528 6058 26580
rect 7374 26568 7380 26580
rect 7335 26540 7380 26568
rect 7374 26528 7380 26540
rect 7432 26528 7438 26580
rect 9033 26571 9091 26577
rect 9033 26537 9045 26571
rect 9079 26568 9091 26571
rect 9214 26568 9220 26580
rect 9079 26540 9220 26568
rect 9079 26537 9091 26540
rect 9033 26531 9091 26537
rect 9214 26528 9220 26540
rect 9272 26528 9278 26580
rect 9674 26528 9680 26580
rect 9732 26568 9738 26580
rect 9953 26571 10011 26577
rect 9953 26568 9965 26571
rect 9732 26540 9965 26568
rect 9732 26528 9738 26540
rect 9953 26537 9965 26540
rect 9999 26537 10011 26571
rect 9953 26531 10011 26537
rect 10686 26528 10692 26580
rect 10744 26568 10750 26580
rect 11057 26571 11115 26577
rect 11057 26568 11069 26571
rect 10744 26540 11069 26568
rect 10744 26528 10750 26540
rect 11057 26537 11069 26540
rect 11103 26568 11115 26571
rect 11974 26568 11980 26580
rect 11103 26540 11980 26568
rect 11103 26537 11115 26540
rect 11057 26531 11115 26537
rect 11974 26528 11980 26540
rect 12032 26528 12038 26580
rect 12250 26568 12256 26580
rect 12211 26540 12256 26568
rect 12250 26528 12256 26540
rect 12308 26528 12314 26580
rect 12342 26528 12348 26580
rect 12400 26568 12406 26580
rect 12805 26571 12863 26577
rect 12805 26568 12817 26571
rect 12400 26540 12817 26568
rect 12400 26528 12406 26540
rect 12805 26537 12817 26540
rect 12851 26537 12863 26571
rect 12805 26531 12863 26537
rect 12986 26528 12992 26580
rect 13044 26568 13050 26580
rect 14737 26571 14795 26577
rect 13044 26540 14688 26568
rect 13044 26528 13050 26540
rect 5718 26500 5724 26512
rect 5276 26472 5724 26500
rect 5276 26441 5304 26472
rect 5718 26460 5724 26472
rect 5776 26500 5782 26512
rect 7282 26500 7288 26512
rect 5776 26472 7288 26500
rect 5776 26460 5782 26472
rect 7282 26460 7288 26472
rect 7340 26460 7346 26512
rect 9122 26500 9128 26512
rect 9083 26472 9128 26500
rect 9122 26460 9128 26472
rect 9180 26460 9186 26512
rect 14274 26460 14280 26512
rect 14332 26500 14338 26512
rect 14553 26503 14611 26509
rect 14553 26500 14565 26503
rect 14332 26472 14565 26500
rect 14332 26460 14338 26472
rect 14553 26469 14565 26472
rect 14599 26469 14611 26503
rect 14660 26500 14688 26540
rect 14737 26537 14749 26571
rect 14783 26568 14795 26571
rect 15194 26568 15200 26580
rect 14783 26540 15200 26568
rect 14783 26537 14795 26540
rect 14737 26531 14795 26537
rect 15194 26528 15200 26540
rect 15252 26528 15258 26580
rect 20993 26571 21051 26577
rect 15304 26540 20944 26568
rect 15304 26500 15332 26540
rect 17954 26500 17960 26512
rect 14660 26472 15332 26500
rect 17915 26472 17960 26500
rect 14553 26463 14611 26469
rect 17954 26460 17960 26472
rect 18012 26460 18018 26512
rect 20806 26500 20812 26512
rect 20719 26472 20812 26500
rect 20806 26460 20812 26472
rect 20864 26460 20870 26512
rect 20916 26500 20944 26540
rect 20993 26537 21005 26571
rect 21039 26568 21051 26571
rect 22646 26568 22652 26580
rect 21039 26540 22652 26568
rect 21039 26537 21051 26540
rect 20993 26531 21051 26537
rect 22646 26528 22652 26540
rect 22704 26528 22710 26580
rect 27430 26528 27436 26580
rect 27488 26568 27494 26580
rect 31846 26568 31852 26580
rect 27488 26540 31852 26568
rect 27488 26528 27494 26540
rect 31846 26528 31852 26540
rect 31904 26528 31910 26580
rect 36446 26528 36452 26580
rect 36504 26568 36510 26580
rect 36725 26571 36783 26577
rect 36725 26568 36737 26571
rect 36504 26540 36737 26568
rect 36504 26528 36510 26540
rect 36725 26537 36737 26540
rect 36771 26537 36783 26571
rect 38194 26568 38200 26580
rect 38155 26540 38200 26568
rect 36725 26531 36783 26537
rect 38194 26528 38200 26540
rect 38252 26528 38258 26580
rect 39301 26571 39359 26577
rect 39301 26537 39313 26571
rect 39347 26568 39359 26571
rect 39666 26568 39672 26580
rect 39347 26540 39672 26568
rect 39347 26537 39359 26540
rect 39301 26531 39359 26537
rect 39666 26528 39672 26540
rect 39724 26528 39730 26580
rect 40770 26568 40776 26580
rect 40731 26540 40776 26568
rect 40770 26528 40776 26540
rect 40828 26528 40834 26580
rect 45002 26528 45008 26580
rect 45060 26568 45066 26580
rect 45097 26571 45155 26577
rect 45097 26568 45109 26571
rect 45060 26540 45109 26568
rect 45060 26528 45066 26540
rect 45097 26537 45109 26540
rect 45143 26537 45155 26571
rect 45097 26531 45155 26537
rect 23566 26500 23572 26512
rect 20916 26472 23572 26500
rect 23566 26460 23572 26472
rect 23624 26460 23630 26512
rect 29362 26460 29368 26512
rect 29420 26500 29426 26512
rect 31665 26503 31723 26509
rect 29420 26472 30144 26500
rect 29420 26460 29426 26472
rect 5261 26435 5319 26441
rect 5261 26401 5273 26435
rect 5307 26401 5319 26435
rect 5442 26432 5448 26444
rect 5403 26404 5448 26432
rect 5261 26395 5319 26401
rect 5442 26392 5448 26404
rect 5500 26392 5506 26444
rect 6825 26435 6883 26441
rect 6825 26401 6837 26435
rect 6871 26432 6883 26435
rect 7098 26432 7104 26444
rect 6871 26404 7104 26432
rect 6871 26401 6883 26404
rect 6825 26395 6883 26401
rect 7098 26392 7104 26404
rect 7156 26432 7162 26444
rect 7558 26432 7564 26444
rect 7156 26404 7564 26432
rect 7156 26392 7162 26404
rect 7558 26392 7564 26404
rect 7616 26392 7622 26444
rect 9766 26392 9772 26444
rect 9824 26432 9830 26444
rect 15378 26432 15384 26444
rect 9824 26404 12940 26432
rect 15339 26404 15384 26432
rect 9824 26392 9830 26404
rect 5166 26364 5172 26376
rect 5127 26336 5172 26364
rect 5166 26324 5172 26336
rect 5224 26324 5230 26376
rect 6181 26367 6239 26373
rect 6181 26333 6193 26367
rect 6227 26364 6239 26367
rect 10226 26364 10232 26376
rect 6227 26336 10232 26364
rect 6227 26333 6239 26336
rect 6181 26327 6239 26333
rect 10226 26324 10232 26336
rect 10284 26324 10290 26376
rect 11900 26373 11928 26404
rect 11885 26367 11943 26373
rect 11885 26333 11897 26367
rect 11931 26333 11943 26367
rect 11885 26327 11943 26333
rect 11974 26324 11980 26376
rect 12032 26364 12038 26376
rect 12032 26336 12204 26364
rect 12032 26324 12038 26336
rect 6914 26296 6920 26308
rect 6875 26268 6920 26296
rect 6914 26256 6920 26268
rect 6972 26256 6978 26308
rect 7009 26299 7067 26305
rect 7009 26265 7021 26299
rect 7055 26296 7067 26299
rect 7742 26296 7748 26308
rect 7055 26268 7748 26296
rect 7055 26265 7067 26268
rect 7009 26259 7067 26265
rect 7742 26256 7748 26268
rect 7800 26256 7806 26308
rect 8294 26256 8300 26308
rect 8352 26296 8358 26308
rect 9493 26299 9551 26305
rect 9493 26296 9505 26299
rect 8352 26268 9505 26296
rect 8352 26256 8358 26268
rect 9493 26265 9505 26268
rect 9539 26296 9551 26299
rect 10594 26296 10600 26308
rect 9539 26268 10600 26296
rect 9539 26265 9551 26268
rect 9493 26259 9551 26265
rect 10594 26256 10600 26268
rect 10652 26256 10658 26308
rect 12066 26296 12072 26308
rect 12027 26268 12072 26296
rect 12066 26256 12072 26268
rect 12124 26256 12130 26308
rect 12176 26296 12204 26336
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12912 26373 12940 26404
rect 15378 26392 15384 26404
rect 15436 26392 15442 26444
rect 19150 26392 19156 26444
rect 19208 26432 19214 26444
rect 19245 26435 19303 26441
rect 19245 26432 19257 26435
rect 19208 26404 19257 26432
rect 19208 26392 19214 26404
rect 19245 26401 19257 26404
rect 19291 26401 19303 26435
rect 19245 26395 19303 26401
rect 20346 26392 20352 26444
rect 20404 26432 20410 26444
rect 20533 26435 20591 26441
rect 20533 26432 20545 26435
rect 20404 26404 20545 26432
rect 20404 26392 20410 26404
rect 20533 26401 20545 26404
rect 20579 26401 20591 26435
rect 20533 26395 20591 26401
rect 12713 26367 12771 26373
rect 12713 26364 12725 26367
rect 12308 26336 12725 26364
rect 12308 26324 12314 26336
rect 12713 26333 12725 26336
rect 12759 26333 12771 26367
rect 12713 26327 12771 26333
rect 12897 26367 12955 26373
rect 12897 26333 12909 26367
rect 12943 26333 12955 26367
rect 17954 26364 17960 26376
rect 16790 26336 17960 26364
rect 12897 26327 12955 26333
rect 17954 26324 17960 26336
rect 18012 26324 18018 26376
rect 18874 26324 18880 26376
rect 18932 26364 18938 26376
rect 19521 26367 19579 26373
rect 19521 26364 19533 26367
rect 18932 26336 19533 26364
rect 18932 26324 18938 26336
rect 19521 26333 19533 26336
rect 19567 26364 19579 26367
rect 20824 26364 20852 26460
rect 23198 26392 23204 26444
rect 23256 26432 23262 26444
rect 23477 26435 23535 26441
rect 23477 26432 23489 26435
rect 23256 26404 23489 26432
rect 23256 26392 23262 26404
rect 23477 26401 23489 26404
rect 23523 26401 23535 26435
rect 23477 26395 23535 26401
rect 24854 26392 24860 26444
rect 24912 26432 24918 26444
rect 24949 26435 25007 26441
rect 24949 26432 24961 26435
rect 24912 26404 24961 26432
rect 24912 26392 24918 26404
rect 24949 26401 24961 26404
rect 24995 26401 25007 26435
rect 25130 26432 25136 26444
rect 24949 26395 25007 26401
rect 25056 26404 25136 26432
rect 19567 26336 20852 26364
rect 19567 26333 19579 26336
rect 19521 26327 19579 26333
rect 23290 26324 23296 26376
rect 23348 26364 23354 26376
rect 23661 26367 23719 26373
rect 23661 26364 23673 26367
rect 23348 26336 23673 26364
rect 23348 26324 23354 26336
rect 23661 26333 23673 26336
rect 23707 26364 23719 26367
rect 25056 26364 25084 26404
rect 25130 26392 25136 26404
rect 25188 26392 25194 26444
rect 30116 26441 30144 26472
rect 31665 26469 31677 26503
rect 31711 26469 31723 26503
rect 31665 26463 31723 26469
rect 39853 26503 39911 26509
rect 39853 26469 39865 26503
rect 39899 26500 39911 26503
rect 40402 26500 40408 26512
rect 39899 26472 40408 26500
rect 39899 26469 39911 26472
rect 39853 26463 39911 26469
rect 28905 26435 28963 26441
rect 28905 26401 28917 26435
rect 28951 26432 28963 26435
rect 30101 26435 30159 26441
rect 28951 26404 29960 26432
rect 28951 26401 28963 26404
rect 28905 26395 28963 26401
rect 25222 26364 25228 26376
rect 23707 26336 25084 26364
rect 25183 26336 25228 26364
rect 23707 26333 23719 26336
rect 23661 26327 23719 26333
rect 25222 26324 25228 26336
rect 25280 26364 25286 26376
rect 25685 26367 25743 26373
rect 25685 26364 25697 26367
rect 25280 26336 25697 26364
rect 25280 26324 25286 26336
rect 25685 26333 25697 26336
rect 25731 26333 25743 26367
rect 28994 26364 29000 26376
rect 28955 26336 29000 26364
rect 25685 26327 25743 26333
rect 28994 26324 29000 26336
rect 29052 26324 29058 26376
rect 29546 26364 29552 26376
rect 29507 26336 29552 26364
rect 29546 26324 29552 26336
rect 29604 26324 29610 26376
rect 29932 26373 29960 26404
rect 30101 26401 30113 26435
rect 30147 26401 30159 26435
rect 30101 26395 30159 26401
rect 31110 26392 31116 26444
rect 31168 26432 31174 26444
rect 31205 26435 31263 26441
rect 31205 26432 31217 26435
rect 31168 26404 31217 26432
rect 31168 26392 31174 26404
rect 31205 26401 31217 26404
rect 31251 26432 31263 26435
rect 31680 26432 31708 26463
rect 40402 26460 40408 26472
rect 40460 26460 40466 26512
rect 40586 26460 40592 26512
rect 40644 26500 40650 26512
rect 41322 26500 41328 26512
rect 40644 26472 41328 26500
rect 40644 26460 40650 26472
rect 41322 26460 41328 26472
rect 41380 26500 41386 26512
rect 41601 26503 41659 26509
rect 41601 26500 41613 26503
rect 41380 26472 41613 26500
rect 41380 26460 41386 26472
rect 41601 26469 41613 26472
rect 41647 26469 41659 26503
rect 68002 26500 68008 26512
rect 67963 26472 68008 26500
rect 41601 26463 41659 26469
rect 68002 26460 68008 26472
rect 68060 26460 68066 26512
rect 32217 26435 32275 26441
rect 32217 26432 32229 26435
rect 31251 26404 31432 26432
rect 31680 26404 32229 26432
rect 31251 26401 31263 26404
rect 31205 26395 31263 26401
rect 29917 26367 29975 26373
rect 29917 26333 29929 26367
rect 29963 26333 29975 26367
rect 29917 26327 29975 26333
rect 31297 26367 31355 26373
rect 31297 26333 31309 26367
rect 31343 26333 31355 26367
rect 31404 26364 31432 26404
rect 32217 26401 32229 26404
rect 32263 26401 32275 26435
rect 32217 26395 32275 26401
rect 42981 26435 43039 26441
rect 42981 26401 42993 26435
rect 43027 26432 43039 26435
rect 43622 26432 43628 26444
rect 43027 26404 43628 26432
rect 43027 26401 43039 26404
rect 42981 26395 43039 26401
rect 43622 26392 43628 26404
rect 43680 26392 43686 26444
rect 32306 26364 32312 26376
rect 31404 26336 32168 26364
rect 32267 26336 32312 26364
rect 31297 26327 31355 26333
rect 13078 26296 13084 26308
rect 12176 26268 13084 26296
rect 13078 26256 13084 26268
rect 13136 26256 13142 26308
rect 13170 26256 13176 26308
rect 13228 26296 13234 26308
rect 13630 26296 13636 26308
rect 13228 26268 13636 26296
rect 13228 26256 13234 26268
rect 13630 26256 13636 26268
rect 13688 26256 13694 26308
rect 13814 26256 13820 26308
rect 13872 26296 13878 26308
rect 14277 26299 14335 26305
rect 14277 26296 14289 26299
rect 13872 26268 14289 26296
rect 13872 26256 13878 26268
rect 14277 26265 14289 26268
rect 14323 26265 14335 26299
rect 15654 26296 15660 26308
rect 15615 26268 15660 26296
rect 14277 26259 14335 26265
rect 15654 26256 15660 26268
rect 15712 26256 15718 26308
rect 17405 26299 17463 26305
rect 17405 26296 17417 26299
rect 16960 26268 17417 26296
rect 15562 26188 15568 26240
rect 15620 26228 15626 26240
rect 16960 26228 16988 26268
rect 17405 26265 17417 26268
rect 17451 26296 17463 26299
rect 20070 26296 20076 26308
rect 17451 26268 20076 26296
rect 17451 26265 17463 26268
rect 17405 26259 17463 26265
rect 20070 26256 20076 26268
rect 20128 26256 20134 26308
rect 29641 26299 29699 26305
rect 29641 26265 29653 26299
rect 29687 26296 29699 26299
rect 30742 26296 30748 26308
rect 29687 26268 30748 26296
rect 29687 26265 29699 26268
rect 29641 26259 29699 26265
rect 30742 26256 30748 26268
rect 30800 26256 30806 26308
rect 31312 26296 31340 26327
rect 31938 26296 31944 26308
rect 31312 26268 31944 26296
rect 31938 26256 31944 26268
rect 31996 26256 32002 26308
rect 32140 26296 32168 26336
rect 32306 26324 32312 26336
rect 32364 26324 32370 26376
rect 34698 26364 34704 26376
rect 34659 26336 34704 26364
rect 34698 26324 34704 26336
rect 34756 26324 34762 26376
rect 34790 26324 34796 26376
rect 34848 26364 34854 26376
rect 34957 26367 35015 26373
rect 34957 26364 34969 26367
rect 34848 26336 34969 26364
rect 34848 26324 34854 26336
rect 34957 26333 34969 26336
rect 35003 26333 35015 26367
rect 37918 26364 37924 26376
rect 37879 26336 37924 26364
rect 34957 26327 35015 26333
rect 37918 26324 37924 26336
rect 37976 26324 37982 26376
rect 38657 26367 38715 26373
rect 38657 26364 38669 26367
rect 38028 26336 38669 26364
rect 38028 26308 38056 26336
rect 38657 26333 38669 26336
rect 38703 26333 38715 26367
rect 38657 26327 38715 26333
rect 38838 26324 38844 26376
rect 38896 26364 38902 26376
rect 39025 26367 39083 26373
rect 39025 26364 39037 26367
rect 38896 26336 39037 26364
rect 38896 26324 38902 26336
rect 39025 26333 39037 26336
rect 39071 26333 39083 26367
rect 39025 26327 39083 26333
rect 39117 26367 39175 26373
rect 39117 26333 39129 26367
rect 39163 26364 39175 26367
rect 39206 26364 39212 26376
rect 39163 26336 39212 26364
rect 39163 26333 39175 26336
rect 39117 26327 39175 26333
rect 39206 26324 39212 26336
rect 39264 26324 39270 26376
rect 40034 26364 40040 26376
rect 39995 26336 40040 26364
rect 40034 26324 40040 26336
rect 40092 26324 40098 26376
rect 40310 26364 40316 26376
rect 40271 26336 40316 26364
rect 40310 26324 40316 26336
rect 40368 26324 40374 26376
rect 40678 26324 40684 26376
rect 40736 26364 40742 26376
rect 40957 26367 41015 26373
rect 40957 26364 40969 26367
rect 40736 26336 40969 26364
rect 40736 26324 40742 26336
rect 40957 26333 40969 26336
rect 41003 26333 41015 26367
rect 41138 26364 41144 26376
rect 41099 26336 41144 26364
rect 40957 26327 41015 26333
rect 41138 26324 41144 26336
rect 41196 26324 41202 26376
rect 42426 26324 42432 26376
rect 42484 26364 42490 26376
rect 42714 26367 42772 26373
rect 42714 26364 42726 26367
rect 42484 26336 42726 26364
rect 42484 26324 42490 26336
rect 42714 26333 42726 26336
rect 42760 26333 42772 26367
rect 42714 26327 42772 26333
rect 45189 26367 45247 26373
rect 45189 26333 45201 26367
rect 45235 26364 45247 26367
rect 45278 26364 45284 26376
rect 45235 26336 45284 26364
rect 45235 26333 45247 26336
rect 45189 26327 45247 26333
rect 45278 26324 45284 26336
rect 45336 26324 45342 26376
rect 67818 26364 67824 26376
rect 67779 26336 67824 26364
rect 67818 26324 67824 26336
rect 67876 26324 67882 26376
rect 32582 26296 32588 26308
rect 32140 26268 32588 26296
rect 32582 26256 32588 26268
rect 32640 26256 32646 26308
rect 36446 26256 36452 26308
rect 36504 26296 36510 26308
rect 36633 26299 36691 26305
rect 36633 26296 36645 26299
rect 36504 26268 36645 26296
rect 36504 26256 36510 26268
rect 36633 26265 36645 26268
rect 36679 26265 36691 26299
rect 38010 26296 38016 26308
rect 37971 26268 38016 26296
rect 36633 26259 36691 26265
rect 38010 26256 38016 26268
rect 38068 26256 38074 26308
rect 38194 26296 38200 26308
rect 38155 26268 38200 26296
rect 38194 26256 38200 26268
rect 38252 26256 38258 26308
rect 40696 26296 40724 26324
rect 40420 26268 40724 26296
rect 15620 26200 16988 26228
rect 23845 26231 23903 26237
rect 15620 26188 15626 26200
rect 23845 26197 23857 26231
rect 23891 26228 23903 26231
rect 24486 26228 24492 26240
rect 23891 26200 24492 26228
rect 23891 26197 23903 26200
rect 23845 26191 23903 26197
rect 24486 26188 24492 26200
rect 24544 26188 24550 26240
rect 32674 26228 32680 26240
rect 32635 26200 32680 26228
rect 32674 26188 32680 26200
rect 32732 26188 32738 26240
rect 36078 26228 36084 26240
rect 36039 26200 36084 26228
rect 36078 26188 36084 26200
rect 36136 26188 36142 26240
rect 37369 26231 37427 26237
rect 37369 26197 37381 26231
rect 37415 26228 37427 26231
rect 37458 26228 37464 26240
rect 37415 26200 37464 26228
rect 37415 26197 37427 26200
rect 37369 26191 37427 26197
rect 37458 26188 37464 26200
rect 37516 26188 37522 26240
rect 40221 26231 40279 26237
rect 40221 26197 40233 26231
rect 40267 26228 40279 26231
rect 40420 26228 40448 26268
rect 40267 26200 40448 26228
rect 40267 26197 40279 26200
rect 40221 26191 40279 26197
rect 1104 26138 68816 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 68816 26138
rect 1104 26064 68816 26086
rect 5718 26024 5724 26036
rect 5679 25996 5724 26024
rect 5718 25984 5724 25996
rect 5776 25984 5782 26036
rect 7285 26027 7343 26033
rect 7285 25993 7297 26027
rect 7331 26024 7343 26027
rect 7926 26024 7932 26036
rect 7331 25996 7932 26024
rect 7331 25993 7343 25996
rect 7285 25987 7343 25993
rect 7926 25984 7932 25996
rect 7984 25984 7990 26036
rect 10502 25984 10508 26036
rect 10560 26024 10566 26036
rect 10597 26027 10655 26033
rect 10597 26024 10609 26027
rect 10560 25996 10609 26024
rect 10560 25984 10566 25996
rect 10597 25993 10609 25996
rect 10643 26024 10655 26027
rect 12434 26024 12440 26036
rect 10643 25996 12440 26024
rect 10643 25993 10655 25996
rect 10597 25987 10655 25993
rect 12434 25984 12440 25996
rect 12492 25984 12498 26036
rect 15378 26024 15384 26036
rect 12636 25996 15384 26024
rect 6362 25916 6368 25968
rect 6420 25956 6426 25968
rect 12636 25965 12664 25996
rect 15378 25984 15384 25996
rect 15436 25984 15442 26036
rect 15654 25984 15660 26036
rect 15712 26024 15718 26036
rect 15933 26027 15991 26033
rect 15933 26024 15945 26027
rect 15712 25996 15945 26024
rect 15712 25984 15718 25996
rect 15933 25993 15945 25996
rect 15979 25993 15991 26027
rect 15933 25987 15991 25993
rect 16945 26027 17003 26033
rect 16945 25993 16957 26027
rect 16991 26024 17003 26027
rect 17126 26024 17132 26036
rect 16991 25996 17132 26024
rect 16991 25993 17003 25996
rect 16945 25987 17003 25993
rect 17126 25984 17132 25996
rect 17184 25984 17190 26036
rect 17405 26027 17463 26033
rect 17405 25993 17417 26027
rect 17451 26024 17463 26027
rect 19426 26024 19432 26036
rect 17451 25996 19432 26024
rect 17451 25993 17463 25996
rect 17405 25987 17463 25993
rect 19426 25984 19432 25996
rect 19484 26024 19490 26036
rect 19794 26024 19800 26036
rect 19484 25996 19800 26024
rect 19484 25984 19490 25996
rect 19794 25984 19800 25996
rect 19852 25984 19858 26036
rect 21913 26027 21971 26033
rect 21913 25993 21925 26027
rect 21959 26024 21971 26027
rect 32125 26027 32183 26033
rect 21959 25996 24716 26024
rect 21959 25993 21971 25996
rect 21913 25987 21971 25993
rect 12621 25959 12679 25965
rect 12621 25956 12633 25959
rect 6420 25928 12633 25956
rect 6420 25916 6426 25928
rect 4890 25888 4896 25900
rect 4851 25860 4896 25888
rect 4890 25848 4896 25860
rect 4948 25848 4954 25900
rect 9232 25897 9260 25928
rect 12621 25925 12633 25928
rect 12667 25925 12679 25959
rect 12621 25919 12679 25925
rect 17034 25916 17040 25968
rect 17092 25956 17098 25968
rect 17313 25959 17371 25965
rect 17313 25956 17325 25959
rect 17092 25928 17325 25956
rect 17092 25916 17098 25928
rect 17313 25925 17325 25928
rect 17359 25956 17371 25959
rect 18046 25956 18052 25968
rect 17359 25928 18052 25956
rect 17359 25925 17371 25928
rect 17313 25919 17371 25925
rect 18046 25916 18052 25928
rect 18104 25916 18110 25968
rect 18230 25956 18236 25968
rect 18191 25928 18236 25956
rect 18230 25916 18236 25928
rect 18288 25916 18294 25968
rect 19521 25959 19579 25965
rect 19521 25925 19533 25959
rect 19567 25956 19579 25959
rect 20346 25956 20352 25968
rect 19567 25928 20352 25956
rect 19567 25925 19579 25928
rect 19521 25919 19579 25925
rect 20346 25916 20352 25928
rect 20404 25916 20410 25968
rect 22738 25956 22744 25968
rect 22699 25928 22744 25956
rect 22738 25916 22744 25928
rect 22796 25916 22802 25968
rect 23385 25959 23443 25965
rect 23385 25925 23397 25959
rect 23431 25956 23443 25959
rect 24581 25959 24639 25965
rect 24581 25956 24593 25959
rect 23431 25928 24593 25956
rect 23431 25925 23443 25928
rect 23385 25919 23443 25925
rect 24581 25925 24593 25928
rect 24627 25925 24639 25959
rect 24581 25919 24639 25925
rect 24688 25900 24716 25996
rect 32125 25993 32137 26027
rect 32171 26024 32183 26027
rect 32306 26024 32312 26036
rect 32171 25996 32312 26024
rect 32171 25993 32183 25996
rect 32125 25987 32183 25993
rect 32306 25984 32312 25996
rect 32364 25984 32370 26036
rect 34514 25984 34520 26036
rect 34572 26024 34578 26036
rect 34701 26027 34759 26033
rect 34701 26024 34713 26027
rect 34572 25996 34713 26024
rect 34572 25984 34578 25996
rect 34701 25993 34713 25996
rect 34747 25993 34759 26027
rect 34701 25987 34759 25993
rect 37921 26027 37979 26033
rect 37921 25993 37933 26027
rect 37967 26024 37979 26027
rect 38194 26024 38200 26036
rect 37967 25996 38200 26024
rect 37967 25993 37979 25996
rect 37921 25987 37979 25993
rect 38194 25984 38200 25996
rect 38252 25984 38258 26036
rect 39485 26027 39543 26033
rect 39485 25993 39497 26027
rect 39531 26024 39543 26027
rect 39850 26024 39856 26036
rect 39531 25996 39856 26024
rect 39531 25993 39543 25996
rect 39485 25987 39543 25993
rect 39850 25984 39856 25996
rect 39908 25984 39914 26036
rect 40589 26027 40647 26033
rect 40589 25993 40601 26027
rect 40635 26024 40647 26027
rect 41046 26024 41052 26036
rect 40635 25996 41052 26024
rect 40635 25993 40647 25996
rect 40589 25987 40647 25993
rect 41046 25984 41052 25996
rect 41104 25984 41110 26036
rect 33226 25916 33232 25968
rect 33284 25965 33290 25968
rect 33284 25956 33296 25965
rect 33284 25928 33329 25956
rect 33284 25919 33296 25928
rect 33284 25916 33290 25919
rect 34606 25916 34612 25968
rect 34664 25956 34670 25968
rect 35069 25959 35127 25965
rect 35069 25956 35081 25959
rect 34664 25928 35081 25956
rect 34664 25916 34670 25928
rect 35069 25925 35081 25928
rect 35115 25925 35127 25959
rect 35069 25919 35127 25925
rect 9490 25897 9496 25900
rect 9217 25891 9275 25897
rect 9217 25857 9229 25891
rect 9263 25857 9275 25891
rect 9217 25851 9275 25857
rect 9484 25851 9496 25897
rect 9548 25888 9554 25900
rect 9548 25860 9584 25888
rect 9490 25848 9496 25851
rect 9548 25848 9554 25860
rect 10594 25848 10600 25900
rect 10652 25888 10658 25900
rect 13170 25888 13176 25900
rect 10652 25860 13176 25888
rect 10652 25848 10658 25860
rect 13170 25848 13176 25860
rect 13228 25848 13234 25900
rect 13357 25891 13415 25897
rect 13357 25857 13369 25891
rect 13403 25888 13415 25891
rect 14090 25888 14096 25900
rect 13403 25860 14096 25888
rect 13403 25857 13415 25860
rect 13357 25851 13415 25857
rect 14090 25848 14096 25860
rect 14148 25848 14154 25900
rect 15381 25891 15439 25897
rect 15381 25857 15393 25891
rect 15427 25888 15439 25891
rect 15562 25888 15568 25900
rect 15427 25860 15568 25888
rect 15427 25857 15439 25860
rect 15381 25851 15439 25857
rect 15562 25848 15568 25860
rect 15620 25848 15626 25900
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25888 16175 25891
rect 16574 25888 16580 25900
rect 16163 25860 16580 25888
rect 16163 25857 16175 25860
rect 16117 25851 16175 25857
rect 16574 25848 16580 25860
rect 16632 25848 16638 25900
rect 19061 25891 19119 25897
rect 19061 25857 19073 25891
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 14274 25820 14280 25832
rect 14235 25792 14280 25820
rect 14274 25780 14280 25792
rect 14332 25780 14338 25832
rect 14734 25820 14740 25832
rect 14695 25792 14740 25820
rect 14734 25780 14740 25792
rect 14792 25780 14798 25832
rect 16482 25780 16488 25832
rect 16540 25820 16546 25832
rect 17497 25823 17555 25829
rect 17497 25820 17509 25823
rect 16540 25792 17509 25820
rect 16540 25780 16546 25792
rect 17497 25789 17509 25792
rect 17543 25789 17555 25823
rect 19076 25820 19104 25851
rect 19426 25848 19432 25900
rect 19484 25888 19490 25900
rect 19705 25891 19763 25897
rect 19705 25888 19717 25891
rect 19484 25860 19717 25888
rect 19484 25848 19490 25860
rect 19705 25857 19717 25860
rect 19751 25857 19763 25891
rect 19705 25851 19763 25857
rect 19794 25848 19800 25900
rect 19852 25888 19858 25900
rect 19852 25860 19897 25888
rect 19852 25848 19858 25860
rect 20530 25848 20536 25900
rect 20588 25888 20594 25900
rect 21821 25891 21879 25897
rect 21821 25888 21833 25891
rect 20588 25860 21833 25888
rect 20588 25848 20594 25860
rect 21821 25857 21833 25860
rect 21867 25857 21879 25891
rect 22002 25888 22008 25900
rect 21963 25860 22008 25888
rect 21821 25851 21879 25857
rect 22002 25848 22008 25860
rect 22060 25848 22066 25900
rect 23106 25848 23112 25900
rect 23164 25888 23170 25900
rect 23293 25891 23351 25897
rect 23293 25888 23305 25891
rect 23164 25860 23305 25888
rect 23164 25848 23170 25860
rect 23293 25857 23305 25860
rect 23339 25857 23351 25891
rect 23293 25851 23351 25857
rect 23477 25891 23535 25897
rect 23477 25857 23489 25891
rect 23523 25857 23535 25891
rect 24210 25888 24216 25900
rect 24171 25860 24216 25888
rect 23477 25851 23535 25857
rect 19076 25792 20392 25820
rect 17497 25783 17555 25789
rect 13814 25712 13820 25764
rect 13872 25752 13878 25764
rect 14553 25755 14611 25761
rect 14553 25752 14565 25755
rect 13872 25724 14565 25752
rect 13872 25712 13878 25724
rect 14553 25721 14565 25724
rect 14599 25721 14611 25755
rect 14553 25715 14611 25721
rect 19334 25712 19340 25764
rect 19392 25752 19398 25764
rect 19521 25755 19579 25761
rect 19521 25752 19533 25755
rect 19392 25724 19533 25752
rect 19392 25712 19398 25724
rect 19521 25721 19533 25724
rect 19567 25721 19579 25755
rect 19521 25715 19579 25721
rect 4706 25684 4712 25696
rect 4667 25656 4712 25684
rect 4706 25644 4712 25656
rect 4764 25644 4770 25696
rect 14918 25644 14924 25696
rect 14976 25684 14982 25696
rect 20364 25693 20392 25792
rect 22738 25780 22744 25832
rect 22796 25820 22802 25832
rect 23492 25820 23520 25851
rect 24210 25848 24216 25860
rect 24268 25848 24274 25900
rect 24361 25891 24419 25897
rect 24361 25857 24373 25891
rect 24407 25888 24419 25891
rect 24407 25857 24440 25888
rect 24361 25851 24440 25857
rect 22796 25792 23520 25820
rect 22796 25780 22802 25792
rect 24412 25752 24440 25851
rect 24486 25848 24492 25900
rect 24544 25888 24550 25900
rect 24544 25860 24589 25888
rect 24544 25848 24550 25860
rect 24670 25848 24676 25900
rect 24728 25897 24734 25900
rect 24728 25888 24736 25897
rect 25498 25888 25504 25900
rect 24728 25860 24821 25888
rect 25459 25860 25504 25888
rect 24728 25851 24736 25860
rect 24728 25848 24734 25851
rect 25498 25848 25504 25860
rect 25556 25848 25562 25900
rect 30561 25891 30619 25897
rect 30561 25857 30573 25891
rect 30607 25888 30619 25891
rect 31205 25891 31263 25897
rect 31205 25888 31217 25891
rect 30607 25860 31217 25888
rect 30607 25857 30619 25860
rect 30561 25851 30619 25857
rect 31205 25857 31217 25860
rect 31251 25888 31263 25891
rect 32766 25888 32772 25900
rect 31251 25860 32772 25888
rect 31251 25857 31263 25860
rect 31205 25851 31263 25857
rect 32766 25848 32772 25860
rect 32824 25848 32830 25900
rect 39298 25888 39304 25900
rect 39259 25860 39304 25888
rect 39298 25848 39304 25860
rect 39356 25848 39362 25900
rect 39485 25891 39543 25897
rect 39485 25857 39497 25891
rect 39531 25857 39543 25891
rect 40218 25888 40224 25900
rect 40179 25860 40224 25888
rect 39485 25851 39543 25857
rect 25406 25820 25412 25832
rect 25367 25792 25412 25820
rect 25406 25780 25412 25792
rect 25464 25780 25470 25832
rect 31297 25823 31355 25829
rect 31297 25789 31309 25823
rect 31343 25820 31355 25823
rect 32030 25820 32036 25832
rect 31343 25792 32036 25820
rect 31343 25789 31355 25792
rect 31297 25783 31355 25789
rect 32030 25780 32036 25792
rect 32088 25780 32094 25832
rect 33502 25820 33508 25832
rect 33463 25792 33508 25820
rect 33502 25780 33508 25792
rect 33560 25780 33566 25832
rect 35161 25823 35219 25829
rect 35161 25789 35173 25823
rect 35207 25789 35219 25823
rect 35161 25783 35219 25789
rect 35345 25823 35403 25829
rect 35345 25789 35357 25823
rect 35391 25820 35403 25823
rect 35434 25820 35440 25832
rect 35391 25792 35440 25820
rect 35391 25789 35403 25792
rect 35345 25783 35403 25789
rect 25590 25752 25596 25764
rect 24412 25724 25596 25752
rect 25590 25712 25596 25724
rect 25648 25712 25654 25764
rect 25869 25755 25927 25761
rect 25869 25721 25881 25755
rect 25915 25752 25927 25755
rect 27522 25752 27528 25764
rect 25915 25724 27528 25752
rect 25915 25721 25927 25724
rect 25869 25715 25927 25721
rect 27522 25712 27528 25724
rect 27580 25712 27586 25764
rect 35176 25752 35204 25783
rect 35434 25780 35440 25792
rect 35492 25780 35498 25832
rect 37458 25820 37464 25832
rect 37419 25792 37464 25820
rect 37458 25780 37464 25792
rect 37516 25780 37522 25832
rect 39500 25820 39528 25851
rect 40218 25848 40224 25860
rect 40276 25848 40282 25900
rect 40405 25891 40463 25897
rect 40405 25857 40417 25891
rect 40451 25888 40463 25891
rect 40770 25888 40776 25900
rect 40451 25860 40776 25888
rect 40451 25857 40463 25860
rect 40405 25851 40463 25857
rect 40770 25848 40776 25860
rect 40828 25848 40834 25900
rect 38764 25792 39528 25820
rect 36078 25752 36084 25764
rect 35176 25724 36084 25752
rect 36078 25712 36084 25724
rect 36136 25752 36142 25764
rect 37734 25752 37740 25764
rect 36136 25724 37740 25752
rect 36136 25712 36142 25724
rect 37734 25712 37740 25724
rect 37792 25712 37798 25764
rect 38764 25696 38792 25792
rect 15289 25687 15347 25693
rect 15289 25684 15301 25687
rect 14976 25656 15301 25684
rect 14976 25644 14982 25656
rect 15289 25653 15301 25656
rect 15335 25653 15347 25687
rect 15289 25647 15347 25653
rect 20349 25687 20407 25693
rect 20349 25653 20361 25687
rect 20395 25684 20407 25687
rect 20438 25684 20444 25696
rect 20395 25656 20444 25684
rect 20395 25653 20407 25656
rect 20349 25647 20407 25653
rect 20438 25644 20444 25656
rect 20496 25644 20502 25696
rect 24854 25684 24860 25696
rect 24815 25656 24860 25684
rect 24854 25644 24860 25656
rect 24912 25644 24918 25696
rect 31481 25687 31539 25693
rect 31481 25653 31493 25687
rect 31527 25684 31539 25687
rect 33226 25684 33232 25696
rect 31527 25656 33232 25684
rect 31527 25653 31539 25656
rect 31481 25647 31539 25653
rect 33226 25644 33232 25656
rect 33284 25644 33290 25696
rect 36446 25684 36452 25696
rect 36407 25656 36452 25684
rect 36446 25644 36452 25656
rect 36504 25644 36510 25696
rect 38746 25684 38752 25696
rect 38707 25656 38752 25684
rect 38746 25644 38752 25656
rect 38804 25644 38810 25696
rect 41046 25644 41052 25696
rect 41104 25684 41110 25696
rect 41506 25684 41512 25696
rect 41104 25656 41512 25684
rect 41104 25644 41110 25656
rect 41506 25644 41512 25656
rect 41564 25644 41570 25696
rect 1104 25594 68816 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 65654 25594
rect 65706 25542 65718 25594
rect 65770 25542 65782 25594
rect 65834 25542 65846 25594
rect 65898 25542 65910 25594
rect 65962 25542 68816 25594
rect 1104 25520 68816 25542
rect 4890 25440 4896 25492
rect 4948 25480 4954 25492
rect 6365 25483 6423 25489
rect 6365 25480 6377 25483
rect 4948 25452 6377 25480
rect 4948 25440 4954 25452
rect 6365 25449 6377 25452
rect 6411 25449 6423 25483
rect 6365 25443 6423 25449
rect 9490 25440 9496 25492
rect 9548 25480 9554 25492
rect 9677 25483 9735 25489
rect 9677 25480 9689 25483
rect 9548 25452 9689 25480
rect 9548 25440 9554 25452
rect 9677 25449 9689 25452
rect 9723 25449 9735 25483
rect 9677 25443 9735 25449
rect 12805 25483 12863 25489
rect 12805 25449 12817 25483
rect 12851 25480 12863 25483
rect 12894 25480 12900 25492
rect 12851 25452 12900 25480
rect 12851 25449 12863 25452
rect 12805 25443 12863 25449
rect 12894 25440 12900 25452
rect 12952 25440 12958 25492
rect 13998 25440 14004 25492
rect 14056 25480 14062 25492
rect 14369 25483 14427 25489
rect 14369 25480 14381 25483
rect 14056 25452 14381 25480
rect 14056 25440 14062 25452
rect 14369 25449 14381 25452
rect 14415 25449 14427 25483
rect 14369 25443 14427 25449
rect 16669 25483 16727 25489
rect 16669 25449 16681 25483
rect 16715 25480 16727 25483
rect 16850 25480 16856 25492
rect 16715 25452 16856 25480
rect 16715 25449 16727 25452
rect 16669 25443 16727 25449
rect 16850 25440 16856 25452
rect 16908 25440 16914 25492
rect 18233 25483 18291 25489
rect 18233 25449 18245 25483
rect 18279 25480 18291 25483
rect 18322 25480 18328 25492
rect 18279 25452 18328 25480
rect 18279 25449 18291 25452
rect 18233 25443 18291 25449
rect 18322 25440 18328 25452
rect 18380 25440 18386 25492
rect 22738 25480 22744 25492
rect 22699 25452 22744 25480
rect 22738 25440 22744 25452
rect 22796 25440 22802 25492
rect 23293 25483 23351 25489
rect 23293 25449 23305 25483
rect 23339 25480 23351 25483
rect 24210 25480 24216 25492
rect 23339 25452 24216 25480
rect 23339 25449 23351 25452
rect 23293 25443 23351 25449
rect 24210 25440 24216 25452
rect 24268 25440 24274 25492
rect 24489 25483 24547 25489
rect 24489 25449 24501 25483
rect 24535 25480 24547 25483
rect 25498 25480 25504 25492
rect 24535 25452 25504 25480
rect 24535 25449 24547 25452
rect 24489 25443 24547 25449
rect 25498 25440 25504 25452
rect 25556 25440 25562 25492
rect 27157 25483 27215 25489
rect 27157 25449 27169 25483
rect 27203 25480 27215 25483
rect 27246 25480 27252 25492
rect 27203 25452 27252 25480
rect 27203 25449 27215 25452
rect 27157 25443 27215 25449
rect 27246 25440 27252 25452
rect 27304 25440 27310 25492
rect 32122 25440 32128 25492
rect 32180 25480 32186 25492
rect 32493 25483 32551 25489
rect 32493 25480 32505 25483
rect 32180 25452 32505 25480
rect 32180 25440 32186 25452
rect 32493 25449 32505 25452
rect 32539 25449 32551 25483
rect 32950 25480 32956 25492
rect 32911 25452 32956 25480
rect 32493 25443 32551 25449
rect 32950 25440 32956 25452
rect 33008 25440 33014 25492
rect 37734 25480 37740 25492
rect 37695 25452 37740 25480
rect 37734 25440 37740 25452
rect 37792 25440 37798 25492
rect 37918 25480 37924 25492
rect 37879 25452 37924 25480
rect 37918 25440 37924 25452
rect 37976 25440 37982 25492
rect 7558 25412 7564 25424
rect 7519 25384 7564 25412
rect 7558 25372 7564 25384
rect 7616 25372 7622 25424
rect 13170 25372 13176 25424
rect 13228 25412 13234 25424
rect 13228 25384 22094 25412
rect 13228 25372 13234 25384
rect 5534 25304 5540 25356
rect 5592 25344 5598 25356
rect 6917 25347 6975 25353
rect 6917 25344 6929 25347
rect 5592 25316 6929 25344
rect 5592 25304 5598 25316
rect 6917 25313 6929 25316
rect 6963 25313 6975 25347
rect 6917 25307 6975 25313
rect 15197 25347 15255 25353
rect 15197 25313 15209 25347
rect 15243 25344 15255 25347
rect 16482 25344 16488 25356
rect 15243 25316 16488 25344
rect 15243 25313 15255 25316
rect 15197 25307 15255 25313
rect 16482 25304 16488 25316
rect 16540 25304 16546 25356
rect 19978 25344 19984 25356
rect 18432 25316 19984 25344
rect 4525 25279 4583 25285
rect 4525 25245 4537 25279
rect 4571 25276 4583 25279
rect 4614 25276 4620 25288
rect 4571 25248 4620 25276
rect 4571 25245 4583 25248
rect 4525 25239 4583 25245
rect 4614 25236 4620 25248
rect 4672 25236 4678 25288
rect 4792 25279 4850 25285
rect 4792 25245 4804 25279
rect 4838 25245 4850 25279
rect 4792 25239 4850 25245
rect 6825 25279 6883 25285
rect 6825 25245 6837 25279
rect 6871 25276 6883 25279
rect 7926 25276 7932 25288
rect 6871 25248 7932 25276
rect 6871 25245 6883 25248
rect 6825 25239 6883 25245
rect 4706 25168 4712 25220
rect 4764 25208 4770 25220
rect 4816 25208 4844 25239
rect 7926 25236 7932 25248
rect 7984 25236 7990 25288
rect 9858 25276 9864 25288
rect 9819 25248 9864 25276
rect 9858 25236 9864 25248
rect 9916 25236 9922 25288
rect 16850 25236 16856 25288
rect 16908 25276 16914 25288
rect 18432 25285 18460 25316
rect 19978 25304 19984 25316
rect 20036 25304 20042 25356
rect 17221 25279 17279 25285
rect 17221 25276 17233 25279
rect 16908 25248 17233 25276
rect 16908 25236 16914 25248
rect 17221 25245 17233 25248
rect 17267 25245 17279 25279
rect 17221 25239 17279 25245
rect 18417 25279 18475 25285
rect 18417 25245 18429 25279
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 18690 25236 18696 25288
rect 18748 25276 18754 25288
rect 19429 25279 19487 25285
rect 19429 25276 19441 25279
rect 18748 25248 19441 25276
rect 18748 25236 18754 25248
rect 19429 25245 19441 25248
rect 19475 25276 19487 25279
rect 20070 25276 20076 25288
rect 19475 25248 20076 25276
rect 19475 25245 19487 25248
rect 19429 25239 19487 25245
rect 20070 25236 20076 25248
rect 20128 25236 20134 25288
rect 22066 25276 22094 25384
rect 22756 25344 22784 25440
rect 30745 25415 30803 25421
rect 30745 25381 30757 25415
rect 30791 25412 30803 25415
rect 31478 25412 31484 25424
rect 30791 25384 31484 25412
rect 30791 25381 30803 25384
rect 30745 25375 30803 25381
rect 31478 25372 31484 25384
rect 31536 25372 31542 25424
rect 22830 25344 22836 25356
rect 22743 25316 22836 25344
rect 22830 25304 22836 25316
rect 22888 25344 22894 25356
rect 22888 25316 23520 25344
rect 22888 25304 22894 25316
rect 23014 25276 23020 25288
rect 22066 25248 23020 25276
rect 23014 25236 23020 25248
rect 23072 25236 23078 25288
rect 23106 25236 23112 25288
rect 23164 25276 23170 25288
rect 23492 25285 23520 25316
rect 24854 25304 24860 25356
rect 24912 25344 24918 25356
rect 24912 25316 27016 25344
rect 24912 25304 24918 25316
rect 23293 25279 23351 25285
rect 23293 25276 23305 25279
rect 23164 25248 23305 25276
rect 23164 25236 23170 25248
rect 23293 25245 23305 25248
rect 23339 25245 23351 25279
rect 23293 25239 23351 25245
rect 23477 25279 23535 25285
rect 23477 25245 23489 25279
rect 23523 25245 23535 25279
rect 24670 25276 24676 25288
rect 24631 25248 24676 25276
rect 23477 25239 23535 25245
rect 24670 25236 24676 25248
rect 24728 25236 24734 25288
rect 24946 25276 24952 25288
rect 24907 25248 24952 25276
rect 24946 25236 24952 25248
rect 25004 25276 25010 25288
rect 25409 25279 25467 25285
rect 25409 25276 25421 25279
rect 25004 25248 25421 25276
rect 25004 25236 25010 25248
rect 25409 25245 25421 25248
rect 25455 25245 25467 25279
rect 25590 25276 25596 25288
rect 25551 25248 25596 25276
rect 25409 25239 25467 25245
rect 25590 25236 25596 25248
rect 25648 25236 25654 25288
rect 25869 25279 25927 25285
rect 25869 25245 25881 25279
rect 25915 25276 25927 25279
rect 26694 25276 26700 25288
rect 25915 25248 26700 25276
rect 25915 25245 25927 25248
rect 25869 25239 25927 25245
rect 26694 25236 26700 25248
rect 26752 25236 26758 25288
rect 26988 25285 27016 25316
rect 30006 25304 30012 25356
rect 30064 25344 30070 25356
rect 30285 25347 30343 25353
rect 30285 25344 30297 25347
rect 30064 25316 30297 25344
rect 30064 25304 30070 25316
rect 30285 25313 30297 25316
rect 30331 25313 30343 25347
rect 31846 25344 31852 25356
rect 31807 25316 31852 25344
rect 30285 25307 30343 25313
rect 31846 25304 31852 25316
rect 31904 25304 31910 25356
rect 32033 25347 32091 25353
rect 32033 25313 32045 25347
rect 32079 25344 32091 25347
rect 32306 25344 32312 25356
rect 32079 25316 32312 25344
rect 32079 25313 32091 25316
rect 32033 25307 32091 25313
rect 32306 25304 32312 25316
rect 32364 25304 32370 25356
rect 33134 25344 33140 25356
rect 33095 25316 33140 25344
rect 33134 25304 33140 25316
rect 33192 25304 33198 25356
rect 26973 25279 27031 25285
rect 26973 25245 26985 25279
rect 27019 25245 27031 25279
rect 26973 25239 27031 25245
rect 29914 25236 29920 25288
rect 29972 25276 29978 25288
rect 30377 25279 30435 25285
rect 30377 25276 30389 25279
rect 29972 25248 30389 25276
rect 29972 25236 29978 25248
rect 30377 25245 30389 25248
rect 30423 25245 30435 25279
rect 30377 25239 30435 25245
rect 32674 25236 32680 25288
rect 32732 25276 32738 25288
rect 32953 25279 33011 25285
rect 32953 25276 32965 25279
rect 32732 25248 32965 25276
rect 32732 25236 32738 25248
rect 32953 25245 32965 25248
rect 32999 25245 33011 25279
rect 33226 25276 33232 25288
rect 33187 25248 33232 25276
rect 32953 25239 33011 25245
rect 33226 25236 33232 25248
rect 33284 25236 33290 25288
rect 37458 25276 37464 25288
rect 36924 25248 37464 25276
rect 4764 25180 4844 25208
rect 7745 25211 7803 25217
rect 4764 25168 4770 25180
rect 7745 25177 7757 25211
rect 7791 25177 7803 25211
rect 14458 25208 14464 25220
rect 14419 25180 14464 25208
rect 7745 25171 7803 25177
rect 5626 25100 5632 25152
rect 5684 25140 5690 25152
rect 5905 25143 5963 25149
rect 5905 25140 5917 25143
rect 5684 25112 5917 25140
rect 5684 25100 5690 25112
rect 5905 25109 5917 25112
rect 5951 25140 5963 25143
rect 6733 25143 6791 25149
rect 6733 25140 6745 25143
rect 5951 25112 6745 25140
rect 5951 25109 5963 25112
rect 5905 25103 5963 25109
rect 6733 25109 6745 25112
rect 6779 25109 6791 25143
rect 7760 25140 7788 25171
rect 14458 25168 14464 25180
rect 14516 25168 14522 25220
rect 17405 25211 17463 25217
rect 17405 25208 17417 25211
rect 16868 25180 17417 25208
rect 16868 25152 16896 25180
rect 17405 25177 17417 25180
rect 17451 25208 17463 25211
rect 20530 25208 20536 25220
rect 17451 25180 20536 25208
rect 17451 25177 17463 25180
rect 17405 25171 17463 25177
rect 20530 25168 20536 25180
rect 20588 25168 20594 25220
rect 24857 25211 24915 25217
rect 24857 25177 24869 25211
rect 24903 25208 24915 25211
rect 25130 25208 25136 25220
rect 24903 25180 25136 25208
rect 24903 25177 24915 25180
rect 24857 25171 24915 25177
rect 25130 25168 25136 25180
rect 25188 25168 25194 25220
rect 32125 25211 32183 25217
rect 32125 25208 32137 25211
rect 31220 25180 32137 25208
rect 31220 25152 31248 25180
rect 32125 25177 32137 25180
rect 32171 25208 32183 25211
rect 34514 25208 34520 25220
rect 32171 25180 34520 25208
rect 32171 25177 32183 25180
rect 32125 25171 32183 25177
rect 34514 25168 34520 25180
rect 34572 25168 34578 25220
rect 8389 25143 8447 25149
rect 8389 25140 8401 25143
rect 7760 25112 8401 25140
rect 6733 25103 6791 25109
rect 8389 25109 8401 25112
rect 8435 25140 8447 25143
rect 11241 25143 11299 25149
rect 11241 25140 11253 25143
rect 8435 25112 11253 25140
rect 8435 25109 8447 25112
rect 8389 25103 8447 25109
rect 11241 25109 11253 25112
rect 11287 25140 11299 25143
rect 11606 25140 11612 25152
rect 11287 25112 11612 25140
rect 11287 25109 11299 25112
rect 11241 25103 11299 25109
rect 11606 25100 11612 25112
rect 11664 25100 11670 25152
rect 11793 25143 11851 25149
rect 11793 25109 11805 25143
rect 11839 25140 11851 25143
rect 11882 25140 11888 25152
rect 11839 25112 11888 25140
rect 11839 25109 11851 25112
rect 11793 25103 11851 25109
rect 11882 25100 11888 25112
rect 11940 25100 11946 25152
rect 13541 25143 13599 25149
rect 13541 25109 13553 25143
rect 13587 25140 13599 25143
rect 14090 25140 14096 25152
rect 13587 25112 14096 25140
rect 13587 25109 13599 25112
rect 13541 25103 13599 25109
rect 14090 25100 14096 25112
rect 14148 25100 14154 25152
rect 15286 25140 15292 25152
rect 15247 25112 15292 25140
rect 15286 25100 15292 25112
rect 15344 25100 15350 25152
rect 15378 25100 15384 25152
rect 15436 25140 15442 25152
rect 15749 25143 15807 25149
rect 15436 25112 15481 25140
rect 15436 25100 15442 25112
rect 15749 25109 15761 25143
rect 15795 25140 15807 25143
rect 15930 25140 15936 25152
rect 15795 25112 15936 25140
rect 15795 25109 15807 25112
rect 15749 25103 15807 25109
rect 15930 25100 15936 25112
rect 15988 25100 15994 25152
rect 16850 25100 16856 25152
rect 16908 25100 16914 25152
rect 19337 25143 19395 25149
rect 19337 25109 19349 25143
rect 19383 25140 19395 25143
rect 19426 25140 19432 25152
rect 19383 25112 19432 25140
rect 19383 25109 19395 25112
rect 19337 25103 19395 25109
rect 19426 25100 19432 25112
rect 19484 25100 19490 25152
rect 25682 25100 25688 25152
rect 25740 25140 25746 25152
rect 25777 25143 25835 25149
rect 25777 25140 25789 25143
rect 25740 25112 25789 25140
rect 25740 25100 25746 25112
rect 25777 25109 25789 25112
rect 25823 25109 25835 25143
rect 25777 25103 25835 25109
rect 26789 25143 26847 25149
rect 26789 25109 26801 25143
rect 26835 25140 26847 25143
rect 27706 25140 27712 25152
rect 26835 25112 27712 25140
rect 26835 25109 26847 25112
rect 26789 25103 26847 25109
rect 27706 25100 27712 25112
rect 27764 25100 27770 25152
rect 31202 25140 31208 25152
rect 31163 25112 31208 25140
rect 31202 25100 31208 25112
rect 31260 25100 31266 25152
rect 33410 25140 33416 25152
rect 33371 25112 33416 25140
rect 33410 25100 33416 25112
rect 33468 25100 33474 25152
rect 35894 25100 35900 25152
rect 35952 25140 35958 25152
rect 36924 25149 36952 25248
rect 37458 25236 37464 25248
rect 37516 25236 37522 25288
rect 60550 25276 60556 25288
rect 60511 25248 60556 25276
rect 60550 25236 60556 25248
rect 60608 25276 60614 25288
rect 61197 25279 61255 25285
rect 61197 25276 61209 25279
rect 60608 25248 61209 25276
rect 60608 25236 60614 25248
rect 61197 25245 61209 25248
rect 61243 25245 61255 25279
rect 61197 25239 61255 25245
rect 67818 25208 67824 25220
rect 60752 25180 67824 25208
rect 60752 25149 60780 25180
rect 67818 25168 67824 25180
rect 67876 25168 67882 25220
rect 36909 25143 36967 25149
rect 36909 25140 36921 25143
rect 35952 25112 36921 25140
rect 35952 25100 35958 25112
rect 36909 25109 36921 25112
rect 36955 25109 36967 25143
rect 36909 25103 36967 25109
rect 60737 25143 60795 25149
rect 60737 25109 60749 25143
rect 60783 25109 60795 25143
rect 60737 25103 60795 25109
rect 1104 25050 68816 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 68816 25050
rect 1104 24976 68816 24998
rect 9858 24896 9864 24948
rect 9916 24936 9922 24948
rect 10137 24939 10195 24945
rect 10137 24936 10149 24939
rect 9916 24908 10149 24936
rect 9916 24896 9922 24908
rect 10137 24905 10149 24908
rect 10183 24905 10195 24939
rect 10502 24936 10508 24948
rect 10463 24908 10508 24936
rect 10137 24899 10195 24905
rect 10502 24896 10508 24908
rect 10560 24896 10566 24948
rect 16482 24896 16488 24948
rect 16540 24936 16546 24948
rect 20714 24936 20720 24948
rect 16540 24908 20720 24936
rect 16540 24896 16546 24908
rect 20714 24896 20720 24908
rect 20772 24936 20778 24948
rect 21450 24936 21456 24948
rect 20772 24908 21456 24936
rect 20772 24896 20778 24908
rect 21450 24896 21456 24908
rect 21508 24896 21514 24948
rect 28994 24896 29000 24948
rect 29052 24936 29058 24948
rect 29052 24908 29316 24936
rect 29052 24896 29058 24908
rect 10686 24828 10692 24880
rect 10744 24868 10750 24880
rect 11517 24871 11575 24877
rect 11517 24868 11529 24871
rect 10744 24840 11529 24868
rect 10744 24828 10750 24840
rect 11517 24837 11529 24840
rect 11563 24837 11575 24871
rect 12894 24868 12900 24880
rect 11517 24831 11575 24837
rect 12406 24840 12900 24868
rect 4893 24803 4951 24809
rect 4893 24769 4905 24803
rect 4939 24800 4951 24803
rect 5166 24800 5172 24812
rect 4939 24772 5172 24800
rect 4939 24769 4951 24772
rect 4893 24763 4951 24769
rect 5166 24760 5172 24772
rect 5224 24760 5230 24812
rect 6908 24803 6966 24809
rect 6908 24769 6920 24803
rect 6954 24800 6966 24803
rect 7374 24800 7380 24812
rect 6954 24772 7380 24800
rect 6954 24769 6966 24772
rect 6908 24763 6966 24769
rect 7374 24760 7380 24772
rect 7432 24760 7438 24812
rect 7926 24760 7932 24812
rect 7984 24800 7990 24812
rect 8481 24803 8539 24809
rect 8481 24800 8493 24803
rect 7984 24772 8493 24800
rect 7984 24760 7990 24772
rect 8481 24769 8493 24772
rect 8527 24769 8539 24803
rect 8481 24763 8539 24769
rect 10597 24803 10655 24809
rect 10597 24769 10609 24803
rect 10643 24800 10655 24803
rect 11882 24800 11888 24812
rect 10643 24772 11888 24800
rect 10643 24769 10655 24772
rect 10597 24763 10655 24769
rect 11882 24760 11888 24772
rect 11940 24760 11946 24812
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 12406 24800 12434 24840
rect 12894 24828 12900 24840
rect 12952 24828 12958 24880
rect 13188 24840 13400 24868
rect 12299 24772 12434 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 12802 24760 12808 24812
rect 12860 24800 12866 24812
rect 13081 24803 13139 24809
rect 13081 24800 13093 24803
rect 12860 24772 13093 24800
rect 12860 24760 12866 24772
rect 13081 24769 13093 24772
rect 13127 24769 13139 24803
rect 13081 24763 13139 24769
rect 4985 24735 5043 24741
rect 4985 24701 4997 24735
rect 5031 24701 5043 24735
rect 6638 24732 6644 24744
rect 6599 24704 6644 24732
rect 4985 24695 5043 24701
rect 4617 24599 4675 24605
rect 4617 24565 4629 24599
rect 4663 24596 4675 24599
rect 4706 24596 4712 24608
rect 4663 24568 4712 24596
rect 4663 24565 4675 24568
rect 4617 24559 4675 24565
rect 4706 24556 4712 24568
rect 4764 24556 4770 24608
rect 5000 24596 5028 24695
rect 6638 24692 6644 24704
rect 6696 24692 6702 24744
rect 10781 24735 10839 24741
rect 10781 24701 10793 24735
rect 10827 24732 10839 24735
rect 11422 24732 11428 24744
rect 10827 24704 11428 24732
rect 10827 24701 10839 24704
rect 10781 24695 10839 24701
rect 11422 24692 11428 24704
rect 11480 24692 11486 24744
rect 12437 24735 12495 24741
rect 12437 24701 12449 24735
rect 12483 24732 12495 24735
rect 12894 24732 12900 24744
rect 12483 24704 12900 24732
rect 12483 24701 12495 24704
rect 12437 24695 12495 24701
rect 12894 24692 12900 24704
rect 12952 24732 12958 24744
rect 13188 24732 13216 24840
rect 13372 24809 13400 24840
rect 13722 24828 13728 24880
rect 13780 24868 13786 24880
rect 17034 24868 17040 24880
rect 13780 24840 17040 24868
rect 13780 24828 13786 24840
rect 17034 24828 17040 24840
rect 17092 24828 17098 24880
rect 19426 24868 19432 24880
rect 19366 24840 19432 24868
rect 19426 24828 19432 24840
rect 19484 24828 19490 24880
rect 29178 24868 29184 24880
rect 28920 24840 29184 24868
rect 13265 24803 13323 24809
rect 13265 24769 13277 24803
rect 13311 24769 13323 24803
rect 13265 24763 13323 24769
rect 13357 24803 13415 24809
rect 13357 24769 13369 24803
rect 13403 24769 13415 24803
rect 13357 24763 13415 24769
rect 14176 24803 14234 24809
rect 14176 24769 14188 24803
rect 14222 24800 14234 24803
rect 15930 24800 15936 24812
rect 14222 24772 15792 24800
rect 15891 24772 15936 24800
rect 14222 24769 14234 24772
rect 14176 24763 14234 24769
rect 12952 24704 13216 24732
rect 13280 24732 13308 24763
rect 13906 24732 13912 24744
rect 13280 24704 13400 24732
rect 13867 24704 13912 24732
rect 12952 24692 12958 24704
rect 9766 24664 9772 24676
rect 7944 24636 9772 24664
rect 7944 24596 7972 24636
rect 9766 24624 9772 24636
rect 9824 24624 9830 24676
rect 5000 24568 7972 24596
rect 8021 24599 8079 24605
rect 8021 24565 8033 24599
rect 8067 24596 8079 24599
rect 9122 24596 9128 24608
rect 8067 24568 9128 24596
rect 8067 24565 8079 24568
rect 8021 24559 8079 24565
rect 9122 24556 9128 24568
rect 9180 24556 9186 24608
rect 13078 24596 13084 24608
rect 13039 24568 13084 24596
rect 13078 24556 13084 24568
rect 13136 24556 13142 24608
rect 13372 24596 13400 24704
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 15764 24673 15792 24772
rect 15930 24760 15936 24772
rect 15988 24760 15994 24812
rect 17218 24800 17224 24812
rect 17179 24772 17224 24800
rect 17218 24760 17224 24772
rect 17276 24760 17282 24812
rect 17405 24803 17463 24809
rect 17405 24769 17417 24803
rect 17451 24800 17463 24803
rect 17586 24800 17592 24812
rect 17451 24772 17592 24800
rect 17451 24769 17463 24772
rect 17405 24763 17463 24769
rect 17586 24760 17592 24772
rect 17644 24760 17650 24812
rect 20070 24760 20076 24812
rect 20128 24800 20134 24812
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 20128 24772 21833 24800
rect 20128 24760 20134 24772
rect 21821 24769 21833 24772
rect 21867 24800 21879 24803
rect 21910 24800 21916 24812
rect 21867 24772 21916 24800
rect 21867 24769 21879 24772
rect 21821 24763 21879 24769
rect 21910 24760 21916 24772
rect 21968 24760 21974 24812
rect 24486 24760 24492 24812
rect 24544 24800 24550 24812
rect 25961 24803 26019 24809
rect 25961 24800 25973 24803
rect 24544 24772 25973 24800
rect 24544 24760 24550 24772
rect 25961 24769 25973 24772
rect 26007 24769 26019 24803
rect 28261 24803 28319 24809
rect 28261 24800 28273 24803
rect 25961 24763 26019 24769
rect 27632 24772 28273 24800
rect 17862 24732 17868 24744
rect 17823 24704 17868 24732
rect 17862 24692 17868 24704
rect 17920 24692 17926 24744
rect 18141 24735 18199 24741
rect 18141 24701 18153 24735
rect 18187 24732 18199 24735
rect 18598 24732 18604 24744
rect 18187 24704 18604 24732
rect 18187 24701 18199 24704
rect 18141 24695 18199 24701
rect 18598 24692 18604 24704
rect 18656 24692 18662 24744
rect 19150 24692 19156 24744
rect 19208 24732 19214 24744
rect 19613 24735 19671 24741
rect 19613 24732 19625 24735
rect 19208 24704 19625 24732
rect 19208 24692 19214 24704
rect 19613 24701 19625 24704
rect 19659 24701 19671 24735
rect 19613 24695 19671 24701
rect 22554 24692 22560 24744
rect 22612 24692 22618 24744
rect 25682 24692 25688 24744
rect 25740 24732 25746 24744
rect 27632 24741 27660 24772
rect 28261 24769 28273 24772
rect 28307 24800 28319 24803
rect 28920 24800 28948 24840
rect 29178 24828 29184 24840
rect 29236 24828 29242 24880
rect 29288 24812 29316 24908
rect 33410 24896 33416 24948
rect 33468 24936 33474 24948
rect 45186 24936 45192 24948
rect 33468 24908 45192 24936
rect 33468 24896 33474 24908
rect 45186 24896 45192 24908
rect 45244 24896 45250 24948
rect 35820 24840 36676 24868
rect 29086 24800 29092 24812
rect 28307 24772 28948 24800
rect 29047 24772 29092 24800
rect 28307 24769 28319 24772
rect 28261 24763 28319 24769
rect 29086 24760 29092 24772
rect 29144 24760 29150 24812
rect 29270 24760 29276 24812
rect 29328 24800 29334 24812
rect 29730 24800 29736 24812
rect 29328 24772 29736 24800
rect 29328 24760 29334 24772
rect 29730 24760 29736 24772
rect 29788 24760 29794 24812
rect 32030 24760 32036 24812
rect 32088 24800 32094 24812
rect 32125 24803 32183 24809
rect 32125 24800 32137 24803
rect 32088 24772 32137 24800
rect 32088 24760 32094 24772
rect 32125 24769 32137 24772
rect 32171 24769 32183 24803
rect 32306 24800 32312 24812
rect 32267 24772 32312 24800
rect 32125 24763 32183 24769
rect 32306 24760 32312 24772
rect 32364 24760 32370 24812
rect 32493 24803 32551 24809
rect 32493 24769 32505 24803
rect 32539 24769 32551 24803
rect 32493 24763 32551 24769
rect 25777 24735 25835 24741
rect 25777 24732 25789 24735
rect 25740 24704 25789 24732
rect 25740 24692 25746 24704
rect 25777 24701 25789 24704
rect 25823 24701 25835 24735
rect 27617 24735 27675 24741
rect 27617 24732 27629 24735
rect 25777 24695 25835 24701
rect 26068 24704 27629 24732
rect 15749 24667 15807 24673
rect 15749 24633 15761 24667
rect 15795 24633 15807 24667
rect 22572 24664 22600 24692
rect 26068 24664 26096 24704
rect 27617 24701 27629 24704
rect 27663 24701 27675 24735
rect 28166 24732 28172 24744
rect 28127 24704 28172 24732
rect 27617 24695 27675 24701
rect 28166 24692 28172 24704
rect 28224 24692 28230 24744
rect 28718 24692 28724 24744
rect 28776 24732 28782 24744
rect 28776 24704 31754 24732
rect 28776 24692 28782 24704
rect 22572 24636 26096 24664
rect 26145 24667 26203 24673
rect 15749 24627 15807 24633
rect 26145 24633 26157 24667
rect 26191 24664 26203 24667
rect 27706 24664 27712 24676
rect 26191 24636 27712 24664
rect 26191 24633 26203 24636
rect 26145 24627 26203 24633
rect 27706 24624 27712 24636
rect 27764 24624 27770 24676
rect 28629 24667 28687 24673
rect 28629 24633 28641 24667
rect 28675 24664 28687 24667
rect 29914 24664 29920 24676
rect 28675 24636 29920 24664
rect 28675 24633 28687 24636
rect 28629 24627 28687 24633
rect 29914 24624 29920 24636
rect 29972 24624 29978 24676
rect 31726 24664 31754 24704
rect 31938 24692 31944 24744
rect 31996 24732 32002 24744
rect 32508 24732 32536 24763
rect 32582 24760 32588 24812
rect 32640 24800 32646 24812
rect 32640 24772 32685 24800
rect 32640 24760 32646 24772
rect 34514 24760 34520 24812
rect 34572 24800 34578 24812
rect 34701 24803 34759 24809
rect 34701 24800 34713 24803
rect 34572 24772 34713 24800
rect 34572 24760 34578 24772
rect 34701 24769 34713 24772
rect 34747 24800 34759 24803
rect 35529 24803 35587 24809
rect 35529 24800 35541 24803
rect 34747 24772 35541 24800
rect 34747 24769 34759 24772
rect 34701 24763 34759 24769
rect 35529 24769 35541 24772
rect 35575 24800 35587 24803
rect 35710 24800 35716 24812
rect 35575 24772 35716 24800
rect 35575 24769 35587 24772
rect 35529 24763 35587 24769
rect 35710 24760 35716 24772
rect 35768 24760 35774 24812
rect 31996 24704 32536 24732
rect 31996 24692 32002 24704
rect 34606 24692 34612 24744
rect 34664 24732 34670 24744
rect 35253 24735 35311 24741
rect 35253 24732 35265 24735
rect 34664 24704 35265 24732
rect 34664 24692 34670 24704
rect 35253 24701 35265 24704
rect 35299 24701 35311 24735
rect 35434 24732 35440 24744
rect 35395 24704 35440 24732
rect 35253 24695 35311 24701
rect 35434 24692 35440 24704
rect 35492 24692 35498 24744
rect 35820 24732 35848 24840
rect 36541 24803 36599 24809
rect 36541 24800 36553 24803
rect 35636 24704 35848 24732
rect 35912 24772 36553 24800
rect 35636 24664 35664 24704
rect 35912 24673 35940 24772
rect 36541 24769 36553 24772
rect 36587 24769 36599 24803
rect 36648 24800 36676 24840
rect 38013 24803 38071 24809
rect 38013 24800 38025 24803
rect 36648 24772 38025 24800
rect 36541 24763 36599 24769
rect 38013 24769 38025 24772
rect 38059 24800 38071 24803
rect 38749 24803 38807 24809
rect 38749 24800 38761 24803
rect 38059 24772 38761 24800
rect 38059 24769 38071 24772
rect 38013 24763 38071 24769
rect 38749 24769 38761 24772
rect 38795 24769 38807 24803
rect 39298 24800 39304 24812
rect 38749 24763 38807 24769
rect 38856 24772 39304 24800
rect 38856 24741 38884 24772
rect 39298 24760 39304 24772
rect 39356 24760 39362 24812
rect 40586 24800 40592 24812
rect 40547 24772 40592 24800
rect 40586 24760 40592 24772
rect 40644 24760 40650 24812
rect 44637 24803 44695 24809
rect 44637 24769 44649 24803
rect 44683 24800 44695 24803
rect 45002 24800 45008 24812
rect 44683 24772 45008 24800
rect 44683 24769 44695 24772
rect 44637 24763 44695 24769
rect 45002 24760 45008 24772
rect 45060 24760 45066 24812
rect 45278 24760 45284 24812
rect 45336 24800 45342 24812
rect 45557 24803 45615 24809
rect 45557 24800 45569 24803
rect 45336 24772 45569 24800
rect 45336 24760 45342 24772
rect 45557 24769 45569 24772
rect 45603 24769 45615 24803
rect 45557 24763 45615 24769
rect 38841 24735 38899 24741
rect 38841 24701 38853 24735
rect 38887 24701 38899 24735
rect 40681 24735 40739 24741
rect 40681 24732 40693 24735
rect 38841 24695 38899 24701
rect 39132 24704 40693 24732
rect 31726 24636 35664 24664
rect 35897 24667 35955 24673
rect 35897 24633 35909 24667
rect 35943 24633 35955 24667
rect 38746 24664 38752 24676
rect 35897 24627 35955 24633
rect 36188 24636 38752 24664
rect 14918 24596 14924 24608
rect 13372 24568 14924 24596
rect 14918 24556 14924 24568
rect 14976 24556 14982 24608
rect 15286 24596 15292 24608
rect 15247 24568 15292 24596
rect 15286 24556 15292 24568
rect 15344 24556 15350 24608
rect 16758 24556 16764 24608
rect 16816 24596 16822 24608
rect 17037 24599 17095 24605
rect 17037 24596 17049 24599
rect 16816 24568 17049 24596
rect 16816 24556 16822 24568
rect 17037 24565 17049 24568
rect 17083 24565 17095 24599
rect 17037 24559 17095 24565
rect 18506 24556 18512 24608
rect 18564 24596 18570 24608
rect 20162 24596 20168 24608
rect 18564 24568 20168 24596
rect 18564 24556 18570 24568
rect 20162 24556 20168 24568
rect 20220 24556 20226 24608
rect 20438 24596 20444 24608
rect 20399 24568 20444 24596
rect 20438 24556 20444 24568
rect 20496 24556 20502 24608
rect 21818 24556 21824 24608
rect 21876 24596 21882 24608
rect 21913 24599 21971 24605
rect 21913 24596 21925 24599
rect 21876 24568 21925 24596
rect 21876 24556 21882 24568
rect 21913 24565 21925 24568
rect 21959 24565 21971 24599
rect 21913 24559 21971 24565
rect 22557 24599 22615 24605
rect 22557 24565 22569 24599
rect 22603 24596 22615 24599
rect 23290 24596 23296 24608
rect 22603 24568 23296 24596
rect 22603 24565 22615 24568
rect 22557 24559 22615 24565
rect 23290 24556 23296 24568
rect 23348 24556 23354 24608
rect 24762 24556 24768 24608
rect 24820 24596 24826 24608
rect 28994 24596 29000 24608
rect 24820 24568 29000 24596
rect 24820 24556 24826 24568
rect 28994 24556 29000 24568
rect 29052 24556 29058 24608
rect 29089 24599 29147 24605
rect 29089 24565 29101 24599
rect 29135 24596 29147 24599
rect 29546 24596 29552 24608
rect 29135 24568 29552 24596
rect 29135 24565 29147 24568
rect 29089 24559 29147 24565
rect 29546 24556 29552 24568
rect 29604 24556 29610 24608
rect 29730 24556 29736 24608
rect 29788 24596 29794 24608
rect 36188 24596 36216 24636
rect 38746 24624 38752 24636
rect 38804 24624 38810 24676
rect 39132 24673 39160 24704
rect 40681 24701 40693 24704
rect 40727 24732 40739 24735
rect 41138 24732 41144 24744
rect 40727 24704 41144 24732
rect 40727 24701 40739 24704
rect 40681 24695 40739 24701
rect 41138 24692 41144 24704
rect 41196 24692 41202 24744
rect 44913 24735 44971 24741
rect 44913 24701 44925 24735
rect 44959 24732 44971 24735
rect 45830 24732 45836 24744
rect 44959 24704 45836 24732
rect 44959 24701 44971 24704
rect 44913 24695 44971 24701
rect 45830 24692 45836 24704
rect 45888 24692 45894 24744
rect 39117 24667 39175 24673
rect 39117 24633 39129 24667
rect 39163 24633 39175 24667
rect 39117 24627 39175 24633
rect 36354 24596 36360 24608
rect 29788 24568 36216 24596
rect 36315 24568 36360 24596
rect 29788 24556 29794 24568
rect 36354 24556 36360 24568
rect 36412 24556 36418 24608
rect 40313 24599 40371 24605
rect 40313 24565 40325 24599
rect 40359 24596 40371 24599
rect 40402 24596 40408 24608
rect 40359 24568 40408 24596
rect 40359 24565 40371 24568
rect 40313 24559 40371 24565
rect 40402 24556 40408 24568
rect 40460 24556 40466 24608
rect 43901 24599 43959 24605
rect 43901 24565 43913 24599
rect 43947 24596 43959 24599
rect 44174 24596 44180 24608
rect 43947 24568 44180 24596
rect 43947 24565 43959 24568
rect 43901 24559 43959 24565
rect 44174 24556 44180 24568
rect 44232 24556 44238 24608
rect 45462 24596 45468 24608
rect 45423 24568 45468 24596
rect 45462 24556 45468 24568
rect 45520 24556 45526 24608
rect 1104 24506 68816 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 65654 24506
rect 65706 24454 65718 24506
rect 65770 24454 65782 24506
rect 65834 24454 65846 24506
rect 65898 24454 65910 24506
rect 65962 24454 68816 24506
rect 1104 24432 68816 24454
rect 9122 24352 9128 24404
rect 9180 24392 9186 24404
rect 12802 24392 12808 24404
rect 9180 24364 12808 24392
rect 9180 24352 9186 24364
rect 12802 24352 12808 24364
rect 12860 24352 12866 24404
rect 16574 24392 16580 24404
rect 16535 24364 16580 24392
rect 16574 24352 16580 24364
rect 16632 24352 16638 24404
rect 17954 24392 17960 24404
rect 17915 24364 17960 24392
rect 17954 24352 17960 24364
rect 18012 24352 18018 24404
rect 29086 24392 29092 24404
rect 18064 24364 29092 24392
rect 15286 24284 15292 24336
rect 15344 24324 15350 24336
rect 18064 24324 18092 24364
rect 15344 24296 18092 24324
rect 15344 24284 15350 24296
rect 18138 24284 18144 24336
rect 18196 24324 18202 24336
rect 18690 24324 18696 24336
rect 18196 24296 18696 24324
rect 18196 24284 18202 24296
rect 18690 24284 18696 24296
rect 18748 24284 18754 24336
rect 23566 24324 23572 24336
rect 23527 24296 23572 24324
rect 23566 24284 23572 24296
rect 23624 24324 23630 24336
rect 24762 24324 24768 24336
rect 23624 24296 24768 24324
rect 23624 24284 23630 24296
rect 24762 24284 24768 24296
rect 24820 24284 24826 24336
rect 25225 24327 25283 24333
rect 25225 24293 25237 24327
rect 25271 24324 25283 24327
rect 25271 24296 25820 24324
rect 25271 24293 25283 24296
rect 25225 24287 25283 24293
rect 25792 24268 25820 24296
rect 4706 24256 4712 24268
rect 4667 24228 4712 24256
rect 4706 24216 4712 24228
rect 4764 24216 4770 24268
rect 7745 24259 7803 24265
rect 7745 24225 7757 24259
rect 7791 24256 7803 24259
rect 7834 24256 7840 24268
rect 7791 24228 7840 24256
rect 7791 24225 7803 24228
rect 7745 24219 7803 24225
rect 7834 24216 7840 24228
rect 7892 24216 7898 24268
rect 7929 24259 7987 24265
rect 7929 24225 7941 24259
rect 7975 24256 7987 24259
rect 11698 24256 11704 24268
rect 7975 24228 11704 24256
rect 7975 24225 7987 24228
rect 7929 24219 7987 24225
rect 11698 24216 11704 24228
rect 11756 24216 11762 24268
rect 14918 24256 14924 24268
rect 14879 24228 14924 24256
rect 14918 24216 14924 24228
rect 14976 24216 14982 24268
rect 17862 24216 17868 24268
rect 17920 24256 17926 24268
rect 20165 24259 20223 24265
rect 20165 24256 20177 24259
rect 17920 24228 20177 24256
rect 17920 24216 17926 24228
rect 20165 24225 20177 24228
rect 20211 24256 20223 24259
rect 20809 24259 20867 24265
rect 20809 24256 20821 24259
rect 20211 24228 20821 24256
rect 20211 24225 20223 24228
rect 20165 24219 20223 24225
rect 20809 24225 20821 24228
rect 20855 24256 20867 24259
rect 22094 24256 22100 24268
rect 20855 24228 22100 24256
rect 20855 24225 20867 24228
rect 20809 24219 20867 24225
rect 22094 24216 22100 24228
rect 22152 24216 22158 24268
rect 22554 24216 22560 24268
rect 22612 24256 22618 24268
rect 22833 24259 22891 24265
rect 22833 24256 22845 24259
rect 22612 24228 22845 24256
rect 22612 24216 22618 24228
rect 22833 24225 22845 24228
rect 22879 24225 22891 24259
rect 22833 24219 22891 24225
rect 24949 24259 25007 24265
rect 24949 24225 24961 24259
rect 24995 24256 25007 24259
rect 25038 24256 25044 24268
rect 24995 24228 25044 24256
rect 24995 24225 25007 24228
rect 24949 24219 25007 24225
rect 25038 24216 25044 24228
rect 25096 24216 25102 24268
rect 25774 24256 25780 24268
rect 25687 24228 25780 24256
rect 25774 24216 25780 24228
rect 25832 24216 25838 24268
rect 28552 24265 28580 24364
rect 29086 24352 29092 24364
rect 29144 24352 29150 24404
rect 29178 24352 29184 24404
rect 29236 24392 29242 24404
rect 29236 24364 30512 24392
rect 29236 24352 29242 24364
rect 28997 24327 29055 24333
rect 28997 24293 29009 24327
rect 29043 24324 29055 24327
rect 30374 24324 30380 24336
rect 29043 24296 30380 24324
rect 29043 24293 29055 24296
rect 28997 24287 29055 24293
rect 30374 24284 30380 24296
rect 30432 24284 30438 24336
rect 30484 24324 30512 24364
rect 30834 24352 30840 24404
rect 30892 24392 30898 24404
rect 30892 24364 35388 24392
rect 30892 24352 30898 24364
rect 34514 24324 34520 24336
rect 30484 24296 34520 24324
rect 34514 24284 34520 24296
rect 34572 24284 34578 24336
rect 34606 24284 34612 24336
rect 34664 24324 34670 24336
rect 34793 24327 34851 24333
rect 34793 24324 34805 24327
rect 34664 24296 34805 24324
rect 34664 24284 34670 24296
rect 34793 24293 34805 24296
rect 34839 24293 34851 24327
rect 35360 24324 35388 24364
rect 35434 24352 35440 24404
rect 35492 24392 35498 24404
rect 37461 24395 37519 24401
rect 37461 24392 37473 24395
rect 35492 24364 37473 24392
rect 35492 24352 35498 24364
rect 37461 24361 37473 24364
rect 37507 24392 37519 24395
rect 37642 24392 37648 24404
rect 37507 24364 37648 24392
rect 37507 24361 37519 24364
rect 37461 24355 37519 24361
rect 37642 24352 37648 24364
rect 37700 24352 37706 24404
rect 40494 24352 40500 24404
rect 40552 24392 40558 24404
rect 43622 24392 43628 24404
rect 40552 24364 43628 24392
rect 40552 24352 40558 24364
rect 43622 24352 43628 24364
rect 43680 24352 43686 24404
rect 45002 24392 45008 24404
rect 44963 24364 45008 24392
rect 45002 24352 45008 24364
rect 45060 24352 45066 24404
rect 35802 24324 35808 24336
rect 35360 24296 35808 24324
rect 34793 24287 34851 24293
rect 35802 24284 35808 24296
rect 35860 24284 35866 24336
rect 45278 24324 45284 24336
rect 44284 24296 45284 24324
rect 28537 24259 28595 24265
rect 28537 24225 28549 24259
rect 28583 24225 28595 24259
rect 28537 24219 28595 24225
rect 28810 24216 28816 24268
rect 28868 24256 28874 24268
rect 32030 24256 32036 24268
rect 28868 24228 32036 24256
rect 28868 24216 28874 24228
rect 32030 24216 32036 24228
rect 32088 24216 32094 24268
rect 33413 24259 33471 24265
rect 33413 24225 33425 24259
rect 33459 24256 33471 24259
rect 34698 24256 34704 24268
rect 33459 24228 34704 24256
rect 33459 24225 33471 24228
rect 33413 24219 33471 24225
rect 34698 24216 34704 24228
rect 34756 24216 34762 24268
rect 35986 24216 35992 24268
rect 36044 24256 36050 24268
rect 36081 24259 36139 24265
rect 36081 24256 36093 24259
rect 36044 24228 36093 24256
rect 36044 24216 36050 24228
rect 36081 24225 36093 24228
rect 36127 24225 36139 24259
rect 36081 24219 36139 24225
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24188 4675 24191
rect 6089 24191 6147 24197
rect 6089 24188 6101 24191
rect 4663 24160 6101 24188
rect 4663 24157 4675 24160
rect 4617 24151 4675 24157
rect 6089 24157 6101 24160
rect 6135 24157 6147 24191
rect 6089 24151 6147 24157
rect 6273 24191 6331 24197
rect 6273 24157 6285 24191
rect 6319 24157 6331 24191
rect 6546 24188 6552 24200
rect 6507 24160 6552 24188
rect 6273 24151 6331 24157
rect 6288 24120 6316 24151
rect 6546 24148 6552 24160
rect 6604 24148 6610 24200
rect 7653 24191 7711 24197
rect 7653 24157 7665 24191
rect 7699 24188 7711 24191
rect 8018 24188 8024 24200
rect 7699 24160 8024 24188
rect 7699 24157 7711 24160
rect 7653 24151 7711 24157
rect 8018 24148 8024 24160
rect 8076 24188 8082 24200
rect 9122 24188 9128 24200
rect 8076 24160 9128 24188
rect 8076 24148 8082 24160
rect 9122 24148 9128 24160
rect 9180 24148 9186 24200
rect 9309 24191 9367 24197
rect 9309 24157 9321 24191
rect 9355 24157 9367 24191
rect 11146 24188 11152 24200
rect 11107 24160 11152 24188
rect 9309 24151 9367 24157
rect 8110 24120 8116 24132
rect 6288 24092 8116 24120
rect 8110 24080 8116 24092
rect 8168 24080 8174 24132
rect 8294 24080 8300 24132
rect 8352 24120 8358 24132
rect 9324 24120 9352 24151
rect 11146 24148 11152 24160
rect 11204 24148 11210 24200
rect 11514 24148 11520 24200
rect 11572 24188 11578 24200
rect 12161 24191 12219 24197
rect 12161 24188 12173 24191
rect 11572 24160 12173 24188
rect 11572 24148 11578 24160
rect 12161 24157 12173 24160
rect 12207 24188 12219 24191
rect 13906 24188 13912 24200
rect 12207 24160 13912 24188
rect 12207 24157 12219 24160
rect 12161 24151 12219 24157
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 14642 24188 14648 24200
rect 14603 24160 14648 24188
rect 14642 24148 14648 24160
rect 14700 24188 14706 24200
rect 15841 24191 15899 24197
rect 14700 24160 15792 24188
rect 14700 24148 14706 24160
rect 9861 24123 9919 24129
rect 9861 24120 9873 24123
rect 8352 24092 9873 24120
rect 8352 24080 8358 24092
rect 9861 24089 9873 24092
rect 9907 24120 9919 24123
rect 12428 24123 12486 24129
rect 9907 24092 11468 24120
rect 9907 24089 9919 24092
rect 9861 24083 9919 24089
rect 4985 24055 5043 24061
rect 4985 24021 4997 24055
rect 5031 24052 5043 24055
rect 5350 24052 5356 24064
rect 5031 24024 5356 24052
rect 5031 24021 5043 24024
rect 4985 24015 5043 24021
rect 5350 24012 5356 24024
rect 5408 24012 5414 24064
rect 6457 24055 6515 24061
rect 6457 24021 6469 24055
rect 6503 24052 6515 24055
rect 6730 24052 6736 24064
rect 6503 24024 6736 24052
rect 6503 24021 6515 24024
rect 6457 24015 6515 24021
rect 6730 24012 6736 24024
rect 6788 24012 6794 24064
rect 7285 24055 7343 24061
rect 7285 24021 7297 24055
rect 7331 24052 7343 24055
rect 7558 24052 7564 24064
rect 7331 24024 7564 24052
rect 7331 24021 7343 24024
rect 7285 24015 7343 24021
rect 7558 24012 7564 24024
rect 7616 24012 7622 24064
rect 8846 24012 8852 24064
rect 8904 24052 8910 24064
rect 8941 24055 8999 24061
rect 8941 24052 8953 24055
rect 8904 24024 8953 24052
rect 8904 24012 8910 24024
rect 8941 24021 8953 24024
rect 8987 24021 8999 24055
rect 8941 24015 8999 24021
rect 9766 24012 9772 24064
rect 9824 24052 9830 24064
rect 10686 24052 10692 24064
rect 9824 24024 10692 24052
rect 9824 24012 9830 24024
rect 10686 24012 10692 24024
rect 10744 24012 10750 24064
rect 11330 24052 11336 24064
rect 11291 24024 11336 24052
rect 11330 24012 11336 24024
rect 11388 24012 11394 24064
rect 11440 24052 11468 24092
rect 12428 24089 12440 24123
rect 12474 24120 12486 24123
rect 13354 24120 13360 24132
rect 12474 24092 13360 24120
rect 12474 24089 12486 24092
rect 12428 24083 12486 24089
rect 13354 24080 13360 24092
rect 13412 24080 13418 24132
rect 15010 24120 15016 24132
rect 13464 24092 15016 24120
rect 13464 24052 13492 24092
rect 15010 24080 15016 24092
rect 15068 24080 15074 24132
rect 15764 24120 15792 24160
rect 15841 24157 15853 24191
rect 15887 24188 15899 24191
rect 16114 24188 16120 24200
rect 15887 24160 16120 24188
rect 15887 24157 15899 24160
rect 15841 24151 15899 24157
rect 16114 24148 16120 24160
rect 16172 24148 16178 24200
rect 16758 24188 16764 24200
rect 16719 24160 16764 24188
rect 16758 24148 16764 24160
rect 16816 24148 16822 24200
rect 16945 24191 17003 24197
rect 16945 24157 16957 24191
rect 16991 24188 17003 24191
rect 17494 24188 17500 24200
rect 16991 24160 17500 24188
rect 16991 24157 17003 24160
rect 16945 24151 17003 24157
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 18049 24191 18107 24197
rect 18049 24157 18061 24191
rect 18095 24188 18107 24191
rect 18138 24188 18144 24200
rect 18095 24160 18144 24188
rect 18095 24157 18107 24160
rect 18049 24151 18107 24157
rect 18138 24148 18144 24160
rect 18196 24148 18202 24200
rect 18506 24188 18512 24200
rect 18467 24160 18512 24188
rect 18506 24148 18512 24160
rect 18564 24148 18570 24200
rect 18693 24191 18751 24197
rect 18693 24157 18705 24191
rect 18739 24157 18751 24191
rect 19426 24188 19432 24200
rect 19339 24160 19432 24188
rect 18693 24151 18751 24157
rect 16390 24120 16396 24132
rect 15764 24092 16396 24120
rect 16390 24080 16396 24092
rect 16448 24080 16454 24132
rect 18708 24120 18736 24151
rect 19426 24148 19432 24160
rect 19484 24188 19490 24200
rect 20438 24188 20444 24200
rect 19484 24160 20444 24188
rect 19484 24148 19490 24160
rect 20438 24148 20444 24160
rect 20496 24148 20502 24200
rect 24857 24191 24915 24197
rect 24857 24157 24869 24191
rect 24903 24157 24915 24191
rect 24857 24151 24915 24157
rect 25947 24191 26005 24197
rect 25947 24157 25959 24191
rect 25993 24188 26005 24191
rect 27338 24188 27344 24200
rect 25993 24160 27344 24188
rect 25993 24157 26005 24160
rect 25947 24151 26005 24157
rect 19334 24120 19340 24132
rect 18708 24092 19340 24120
rect 19334 24080 19340 24092
rect 19392 24080 19398 24132
rect 21082 24120 21088 24132
rect 21043 24092 21088 24120
rect 21082 24080 21088 24092
rect 21140 24080 21146 24132
rect 21818 24080 21824 24132
rect 21876 24080 21882 24132
rect 23382 24120 23388 24132
rect 23343 24092 23388 24120
rect 23382 24080 23388 24092
rect 23440 24080 23446 24132
rect 24578 24080 24584 24132
rect 24636 24120 24642 24132
rect 24872 24120 24900 24151
rect 27338 24148 27344 24160
rect 27396 24148 27402 24200
rect 28718 24197 28724 24200
rect 27985 24191 28043 24197
rect 27985 24157 27997 24191
rect 28031 24188 28043 24191
rect 28707 24191 28724 24197
rect 28707 24188 28719 24191
rect 28031 24160 28719 24188
rect 28031 24157 28043 24160
rect 27985 24151 28043 24157
rect 28707 24157 28719 24160
rect 28707 24151 28724 24157
rect 24636 24092 27200 24120
rect 24636 24080 24642 24092
rect 11440 24024 13492 24052
rect 13541 24055 13599 24061
rect 13541 24021 13553 24055
rect 13587 24052 13599 24055
rect 13814 24052 13820 24064
rect 13587 24024 13820 24052
rect 13587 24021 13599 24024
rect 13541 24015 13599 24021
rect 13814 24012 13820 24024
rect 13872 24012 13878 24064
rect 15654 24052 15660 24064
rect 15615 24024 15660 24052
rect 15654 24012 15660 24024
rect 15712 24012 15718 24064
rect 18506 24012 18512 24064
rect 18564 24052 18570 24064
rect 18601 24055 18659 24061
rect 18601 24052 18613 24055
rect 18564 24024 18613 24052
rect 18564 24012 18570 24024
rect 18601 24021 18613 24024
rect 18647 24021 18659 24055
rect 18601 24015 18659 24021
rect 26237 24055 26295 24061
rect 26237 24021 26249 24055
rect 26283 24052 26295 24055
rect 27062 24052 27068 24064
rect 26283 24024 27068 24052
rect 26283 24021 26295 24024
rect 26237 24015 26295 24021
rect 27062 24012 27068 24024
rect 27120 24012 27126 24064
rect 27172 24052 27200 24092
rect 27246 24080 27252 24132
rect 27304 24120 27310 24132
rect 28000 24120 28028 24151
rect 28718 24148 28724 24151
rect 28776 24148 28782 24200
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 28828 24160 29561 24188
rect 27304 24092 28028 24120
rect 27304 24080 27310 24092
rect 28166 24080 28172 24132
rect 28224 24120 28230 24132
rect 28828 24120 28856 24160
rect 29549 24157 29561 24160
rect 29595 24157 29607 24191
rect 29549 24151 29607 24157
rect 29733 24191 29791 24197
rect 29733 24157 29745 24191
rect 29779 24188 29791 24191
rect 30282 24188 30288 24200
rect 29779 24160 30288 24188
rect 29779 24157 29791 24160
rect 29733 24151 29791 24157
rect 30282 24148 30288 24160
rect 30340 24148 30346 24200
rect 35894 24188 35900 24200
rect 31726 24160 35900 24188
rect 31726 24120 31754 24160
rect 35894 24148 35900 24160
rect 35952 24148 35958 24200
rect 36096 24188 36124 24219
rect 39758 24216 39764 24268
rect 39816 24256 39822 24268
rect 42705 24259 42763 24265
rect 42705 24256 42717 24259
rect 39816 24228 42717 24256
rect 39816 24216 39822 24228
rect 42705 24225 42717 24228
rect 42751 24225 42763 24259
rect 42705 24219 42763 24225
rect 44284 24200 44312 24296
rect 45278 24284 45284 24296
rect 45336 24284 45342 24336
rect 45830 24284 45836 24336
rect 45888 24324 45894 24336
rect 46842 24324 46848 24336
rect 45888 24296 46848 24324
rect 45888 24284 45894 24296
rect 46842 24284 46848 24296
rect 46900 24324 46906 24336
rect 47121 24327 47179 24333
rect 47121 24324 47133 24327
rect 46900 24296 47133 24324
rect 46900 24284 46906 24296
rect 47121 24293 47133 24296
rect 47167 24293 47179 24327
rect 47121 24287 47179 24293
rect 45186 24256 45192 24268
rect 45147 24228 45192 24256
rect 45186 24216 45192 24228
rect 45244 24216 45250 24268
rect 46014 24216 46020 24268
rect 46072 24256 46078 24268
rect 46072 24228 46336 24256
rect 46072 24216 46078 24228
rect 38562 24188 38568 24200
rect 36096 24160 38568 24188
rect 38562 24148 38568 24160
rect 38620 24188 38626 24200
rect 40494 24188 40500 24200
rect 38620 24160 40500 24188
rect 38620 24148 38626 24160
rect 40494 24148 40500 24160
rect 40552 24148 40558 24200
rect 42981 24191 43039 24197
rect 42981 24157 42993 24191
rect 43027 24157 43039 24191
rect 42981 24151 43039 24157
rect 43809 24191 43867 24197
rect 43809 24157 43821 24191
rect 43855 24157 43867 24191
rect 44266 24188 44272 24200
rect 44179 24160 44272 24188
rect 43809 24151 43867 24157
rect 36354 24129 36360 24132
rect 28224 24092 28856 24120
rect 28920 24092 31754 24120
rect 34149 24123 34207 24129
rect 28224 24080 28230 24092
rect 28920 24052 28948 24092
rect 34149 24089 34161 24123
rect 34195 24089 34207 24123
rect 36348 24120 36360 24129
rect 36315 24092 36360 24120
rect 34149 24083 34207 24089
rect 36348 24083 36360 24092
rect 27172 24024 28948 24052
rect 29641 24055 29699 24061
rect 29641 24021 29653 24055
rect 29687 24052 29699 24055
rect 30098 24052 30104 24064
rect 29687 24024 30104 24052
rect 29687 24021 29699 24024
rect 29641 24015 29699 24021
rect 30098 24012 30104 24024
rect 30156 24012 30162 24064
rect 32769 24055 32827 24061
rect 32769 24021 32781 24055
rect 32815 24052 32827 24055
rect 32858 24052 32864 24064
rect 32815 24024 32864 24052
rect 32815 24021 32827 24024
rect 32769 24015 32827 24021
rect 32858 24012 32864 24024
rect 32916 24052 32922 24064
rect 34164 24052 34192 24083
rect 36354 24080 36360 24083
rect 36412 24080 36418 24132
rect 40770 24120 40776 24132
rect 40731 24092 40776 24120
rect 40770 24080 40776 24092
rect 40828 24080 40834 24132
rect 42518 24120 42524 24132
rect 41998 24092 42524 24120
rect 42518 24080 42524 24092
rect 42576 24080 42582 24132
rect 32916 24024 34192 24052
rect 32916 24012 32922 24024
rect 34514 24012 34520 24064
rect 34572 24052 34578 24064
rect 38102 24052 38108 24064
rect 34572 24024 38108 24052
rect 34572 24012 34578 24024
rect 38102 24012 38108 24024
rect 38160 24012 38166 24064
rect 42242 24052 42248 24064
rect 42203 24024 42248 24052
rect 42242 24012 42248 24024
rect 42300 24012 42306 24064
rect 42334 24012 42340 24064
rect 42392 24052 42398 24064
rect 42996 24052 43024 24151
rect 43824 24120 43852 24151
rect 44266 24148 44272 24160
rect 44324 24148 44330 24200
rect 45278 24148 45284 24200
rect 45336 24188 45342 24200
rect 46308 24197 46336 24228
rect 46201 24191 46259 24197
rect 45336 24160 45381 24188
rect 45336 24148 45342 24160
rect 46201 24157 46213 24191
rect 46247 24157 46259 24191
rect 46201 24151 46259 24157
rect 46293 24191 46351 24197
rect 46293 24157 46305 24191
rect 46339 24157 46351 24191
rect 46293 24151 46351 24157
rect 46477 24191 46535 24197
rect 46477 24157 46489 24191
rect 46523 24188 46535 24191
rect 46937 24191 46995 24197
rect 46937 24188 46949 24191
rect 46523 24160 46949 24188
rect 46523 24157 46535 24160
rect 46477 24151 46535 24157
rect 46937 24157 46949 24160
rect 46983 24157 46995 24191
rect 46937 24151 46995 24157
rect 44082 24120 44088 24132
rect 43824 24092 44088 24120
rect 44082 24080 44088 24092
rect 44140 24120 44146 24132
rect 44726 24120 44732 24132
rect 44140 24092 44732 24120
rect 44140 24080 44146 24092
rect 44726 24080 44732 24092
rect 44784 24080 44790 24132
rect 42392 24024 43024 24052
rect 44361 24055 44419 24061
rect 42392 24012 42398 24024
rect 44361 24021 44373 24055
rect 44407 24052 44419 24055
rect 44634 24052 44640 24064
rect 44407 24024 44640 24052
rect 44407 24021 44419 24024
rect 44361 24015 44419 24021
rect 44634 24012 44640 24024
rect 44692 24012 44698 24064
rect 45646 24052 45652 24064
rect 45607 24024 45652 24052
rect 45646 24012 45652 24024
rect 45704 24012 45710 24064
rect 46216 24052 46244 24151
rect 46934 24052 46940 24064
rect 46216 24024 46940 24052
rect 46934 24012 46940 24024
rect 46992 24012 46998 24064
rect 1104 23962 68816 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 68816 23962
rect 1104 23888 68816 23910
rect 7374 23848 7380 23860
rect 7335 23820 7380 23848
rect 7374 23808 7380 23820
rect 7432 23808 7438 23860
rect 8110 23848 8116 23860
rect 8071 23820 8116 23848
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 9953 23851 10011 23857
rect 9953 23817 9965 23851
rect 9999 23848 10011 23851
rect 10870 23848 10876 23860
rect 9999 23820 10876 23848
rect 9999 23817 10011 23820
rect 9953 23811 10011 23817
rect 10870 23808 10876 23820
rect 10928 23808 10934 23860
rect 12894 23848 12900 23860
rect 12855 23820 12900 23848
rect 12894 23808 12900 23820
rect 12952 23808 12958 23860
rect 13354 23848 13360 23860
rect 13315 23820 13360 23848
rect 13354 23808 13360 23820
rect 13412 23808 13418 23860
rect 14090 23848 14096 23860
rect 14003 23820 14096 23848
rect 14090 23808 14096 23820
rect 14148 23848 14154 23860
rect 19426 23848 19432 23860
rect 14148 23820 19432 23848
rect 14148 23808 14154 23820
rect 19426 23808 19432 23820
rect 19484 23808 19490 23860
rect 20901 23851 20959 23857
rect 20901 23817 20913 23851
rect 20947 23848 20959 23851
rect 21082 23848 21088 23860
rect 20947 23820 21088 23848
rect 20947 23817 20959 23820
rect 20901 23811 20959 23817
rect 21082 23808 21088 23820
rect 21140 23808 21146 23860
rect 22830 23848 22836 23860
rect 22791 23820 22836 23848
rect 22830 23808 22836 23820
rect 22888 23808 22894 23860
rect 23014 23808 23020 23860
rect 23072 23848 23078 23860
rect 23750 23848 23756 23860
rect 23072 23820 23756 23848
rect 23072 23808 23078 23820
rect 23750 23808 23756 23820
rect 23808 23848 23814 23860
rect 24578 23848 24584 23860
rect 23808 23820 24584 23848
rect 23808 23808 23814 23820
rect 24578 23808 24584 23820
rect 24636 23808 24642 23860
rect 25682 23848 25688 23860
rect 25643 23820 25688 23848
rect 25682 23808 25688 23820
rect 25740 23808 25746 23860
rect 26602 23808 26608 23860
rect 26660 23848 26666 23860
rect 28537 23851 28595 23857
rect 26660 23820 28488 23848
rect 26660 23808 26666 23820
rect 5626 23780 5632 23792
rect 5000 23752 5632 23780
rect 5000 23721 5028 23752
rect 5626 23740 5632 23752
rect 5684 23740 5690 23792
rect 8128 23780 8156 23808
rect 8128 23752 8708 23780
rect 4801 23715 4859 23721
rect 4801 23681 4813 23715
rect 4847 23681 4859 23715
rect 4801 23675 4859 23681
rect 4985 23715 5043 23721
rect 4985 23681 4997 23715
rect 5031 23681 5043 23715
rect 4985 23675 5043 23681
rect 5445 23715 5503 23721
rect 5445 23681 5457 23715
rect 5491 23681 5503 23715
rect 6730 23712 6736 23724
rect 6691 23684 6736 23712
rect 5445 23675 5503 23681
rect 4816 23644 4844 23675
rect 5460 23644 5488 23675
rect 6730 23672 6736 23684
rect 6788 23672 6794 23724
rect 7558 23712 7564 23724
rect 7519 23684 7564 23712
rect 7558 23672 7564 23684
rect 7616 23672 7622 23724
rect 8018 23712 8024 23724
rect 7979 23684 8024 23712
rect 8018 23672 8024 23684
rect 8076 23672 8082 23724
rect 8205 23715 8263 23721
rect 8205 23681 8217 23715
rect 8251 23712 8263 23715
rect 8294 23712 8300 23724
rect 8251 23684 8300 23712
rect 8251 23681 8263 23684
rect 8205 23675 8263 23681
rect 8294 23672 8300 23684
rect 8352 23672 8358 23724
rect 8680 23721 8708 23752
rect 10134 23740 10140 23792
rect 10192 23780 10198 23792
rect 10192 23752 10824 23780
rect 10192 23740 10198 23752
rect 8665 23715 8723 23721
rect 8665 23681 8677 23715
rect 8711 23681 8723 23715
rect 8846 23712 8852 23724
rect 8807 23684 8852 23712
rect 8665 23675 8723 23681
rect 8846 23672 8852 23684
rect 8904 23672 8910 23724
rect 9766 23712 9772 23724
rect 9727 23684 9772 23712
rect 9766 23672 9772 23684
rect 9824 23672 9830 23724
rect 10686 23712 10692 23724
rect 9944 23705 10002 23711
rect 9944 23702 9956 23705
rect 9876 23674 9956 23702
rect 6365 23647 6423 23653
rect 6365 23644 6377 23647
rect 4816 23616 6377 23644
rect 6365 23613 6377 23616
rect 6411 23613 6423 23647
rect 6365 23607 6423 23613
rect 6546 23604 6552 23656
rect 6604 23644 6610 23656
rect 6641 23647 6699 23653
rect 6641 23644 6653 23647
rect 6604 23616 6653 23644
rect 6604 23604 6610 23616
rect 6641 23613 6653 23616
rect 6687 23613 6699 23647
rect 6748 23644 6776 23672
rect 8757 23647 8815 23653
rect 8757 23644 8769 23647
rect 6748 23616 8769 23644
rect 6641 23607 6699 23613
rect 8757 23613 8769 23616
rect 8803 23644 8815 23647
rect 8803 23616 9674 23644
rect 8803 23613 8815 23616
rect 8757 23607 8815 23613
rect 4893 23579 4951 23585
rect 4893 23545 4905 23579
rect 4939 23576 4951 23579
rect 5718 23576 5724 23588
rect 4939 23548 5724 23576
rect 4939 23545 4951 23548
rect 4893 23539 4951 23545
rect 5718 23536 5724 23548
rect 5776 23536 5782 23588
rect 6656 23576 6684 23607
rect 9646 23576 9674 23616
rect 9876 23576 9904 23674
rect 9944 23671 9956 23674
rect 9990 23671 10002 23705
rect 10647 23684 10692 23712
rect 10686 23672 10692 23684
rect 10744 23672 10750 23724
rect 10796 23721 10824 23752
rect 11330 23740 11336 23792
rect 11388 23780 11394 23792
rect 11762 23783 11820 23789
rect 11762 23780 11774 23783
rect 11388 23752 11774 23780
rect 11388 23740 11394 23752
rect 11762 23749 11774 23752
rect 11808 23749 11820 23783
rect 11762 23743 11820 23749
rect 11882 23740 11888 23792
rect 11940 23780 11946 23792
rect 17126 23780 17132 23792
rect 11940 23752 17132 23780
rect 11940 23740 11946 23752
rect 17126 23740 17132 23752
rect 17184 23740 17190 23792
rect 17494 23780 17500 23792
rect 17455 23752 17500 23780
rect 17494 23740 17500 23752
rect 17552 23740 17558 23792
rect 18598 23780 18604 23792
rect 18559 23752 18604 23780
rect 18598 23740 18604 23752
rect 18656 23740 18662 23792
rect 22097 23783 22155 23789
rect 22097 23749 22109 23783
rect 22143 23780 22155 23783
rect 22741 23783 22799 23789
rect 22741 23780 22753 23783
rect 22143 23752 22753 23780
rect 22143 23749 22155 23752
rect 22097 23743 22155 23749
rect 22741 23749 22753 23752
rect 22787 23780 22799 23783
rect 23382 23780 23388 23792
rect 22787 23752 23388 23780
rect 22787 23749 22799 23752
rect 22741 23743 22799 23749
rect 23382 23740 23388 23752
rect 23440 23740 23446 23792
rect 27246 23780 27252 23792
rect 23676 23752 27252 23780
rect 10781 23715 10839 23721
rect 10781 23681 10793 23715
rect 10827 23681 10839 23715
rect 10781 23675 10839 23681
rect 10873 23715 10931 23721
rect 10873 23681 10885 23715
rect 10919 23712 10931 23715
rect 12526 23712 12532 23724
rect 10919 23684 12532 23712
rect 10919 23681 10931 23684
rect 10873 23675 10931 23681
rect 12526 23672 12532 23684
rect 12584 23672 12590 23724
rect 13541 23715 13599 23721
rect 13541 23681 13553 23715
rect 13587 23712 13599 23715
rect 13998 23712 14004 23724
rect 13587 23684 14004 23712
rect 13587 23681 13599 23684
rect 13541 23675 13599 23681
rect 13998 23672 14004 23684
rect 14056 23672 14062 23724
rect 15194 23672 15200 23724
rect 15252 23712 15258 23724
rect 15749 23715 15807 23721
rect 15749 23712 15761 23715
rect 15252 23684 15761 23712
rect 15252 23672 15258 23684
rect 15749 23681 15761 23684
rect 15795 23712 15807 23715
rect 15838 23712 15844 23724
rect 15795 23684 15844 23712
rect 15795 23681 15807 23684
rect 15749 23675 15807 23681
rect 15838 23672 15844 23684
rect 15896 23712 15902 23724
rect 16669 23715 16727 23721
rect 16669 23712 16681 23715
rect 15896 23684 16681 23712
rect 15896 23672 15902 23684
rect 16669 23681 16681 23684
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 17218 23672 17224 23724
rect 17276 23712 17282 23724
rect 17405 23715 17463 23721
rect 17405 23712 17417 23715
rect 17276 23684 17417 23712
rect 17276 23672 17282 23684
rect 17405 23681 17417 23684
rect 17451 23681 17463 23715
rect 17586 23712 17592 23724
rect 17547 23684 17592 23712
rect 17405 23675 17463 23681
rect 17586 23672 17592 23684
rect 17644 23672 17650 23724
rect 18506 23712 18512 23724
rect 18467 23684 18512 23712
rect 18506 23672 18512 23684
rect 18564 23672 18570 23724
rect 18693 23715 18751 23721
rect 18693 23681 18705 23715
rect 18739 23681 18751 23715
rect 18693 23675 18751 23681
rect 9944 23665 10002 23671
rect 10597 23647 10655 23653
rect 10597 23613 10609 23647
rect 10643 23613 10655 23647
rect 11514 23644 11520 23656
rect 11475 23616 11520 23644
rect 10597 23607 10655 23613
rect 10134 23576 10140 23588
rect 6656 23548 9168 23576
rect 9646 23548 10140 23576
rect 9140 23520 9168 23548
rect 10134 23536 10140 23548
rect 10192 23536 10198 23588
rect 10612 23576 10640 23607
rect 11514 23604 11520 23616
rect 11572 23604 11578 23656
rect 15565 23647 15623 23653
rect 15565 23613 15577 23647
rect 15611 23613 15623 23647
rect 15565 23607 15623 23613
rect 15657 23647 15715 23653
rect 15657 23613 15669 23647
rect 15703 23644 15715 23647
rect 16758 23644 16764 23656
rect 15703 23616 16764 23644
rect 15703 23613 15715 23616
rect 15657 23607 15715 23613
rect 10244 23548 10640 23576
rect 5810 23508 5816 23520
rect 5771 23480 5816 23508
rect 5810 23468 5816 23480
rect 5868 23468 5874 23520
rect 9122 23468 9128 23520
rect 9180 23508 9186 23520
rect 10244 23508 10272 23548
rect 10410 23508 10416 23520
rect 9180 23480 10272 23508
rect 10371 23480 10416 23508
rect 9180 23468 9186 23480
rect 10410 23468 10416 23480
rect 10468 23468 10474 23520
rect 15580 23508 15608 23607
rect 16758 23604 16764 23616
rect 16816 23604 16822 23656
rect 17604 23644 17632 23672
rect 18046 23644 18052 23656
rect 17604 23616 18052 23644
rect 18046 23604 18052 23616
rect 18104 23644 18110 23656
rect 18708 23644 18736 23675
rect 19978 23672 19984 23724
rect 20036 23712 20042 23724
rect 20530 23712 20536 23724
rect 20036 23684 20536 23712
rect 20036 23672 20042 23684
rect 20530 23672 20536 23684
rect 20588 23672 20594 23724
rect 23676 23721 23704 23752
rect 27246 23740 27252 23752
rect 27304 23740 27310 23792
rect 27522 23740 27528 23792
rect 27580 23780 27586 23792
rect 28077 23783 28135 23789
rect 28077 23780 28089 23783
rect 27580 23752 28089 23780
rect 27580 23740 27586 23752
rect 28077 23749 28089 23752
rect 28123 23749 28135 23783
rect 28077 23743 28135 23749
rect 22189 23715 22247 23721
rect 22189 23681 22201 23715
rect 22235 23712 22247 23715
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 22235 23684 23673 23712
rect 22235 23681 22247 23684
rect 22189 23675 22247 23681
rect 23400 23656 23428 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 25774 23672 25780 23724
rect 25832 23712 25838 23724
rect 25869 23715 25927 23721
rect 25869 23712 25881 23715
rect 25832 23684 25881 23712
rect 25832 23672 25838 23684
rect 25869 23681 25881 23684
rect 25915 23681 25927 23715
rect 27154 23712 27160 23724
rect 27115 23684 27160 23712
rect 25869 23675 25927 23681
rect 27154 23672 27160 23684
rect 27212 23672 27218 23724
rect 28353 23715 28411 23721
rect 28353 23712 28365 23715
rect 27540 23684 28365 23712
rect 19242 23644 19248 23656
rect 18104 23616 19248 23644
rect 18104 23604 18110 23616
rect 19242 23604 19248 23616
rect 19300 23604 19306 23656
rect 20441 23647 20499 23653
rect 20441 23613 20453 23647
rect 20487 23613 20499 23647
rect 20441 23607 20499 23613
rect 16114 23576 16120 23588
rect 16075 23548 16120 23576
rect 16114 23536 16120 23548
rect 16172 23536 16178 23588
rect 16390 23536 16396 23588
rect 16448 23576 16454 23588
rect 19150 23576 19156 23588
rect 16448 23548 19156 23576
rect 16448 23536 16454 23548
rect 19150 23536 19156 23548
rect 19208 23536 19214 23588
rect 20456 23576 20484 23607
rect 23382 23604 23388 23656
rect 23440 23604 23446 23656
rect 26050 23644 26056 23656
rect 26011 23616 26056 23644
rect 26050 23604 26056 23616
rect 26108 23604 26114 23656
rect 27062 23644 27068 23656
rect 27023 23616 27068 23644
rect 27062 23604 27068 23616
rect 27120 23604 27126 23656
rect 20530 23576 20536 23588
rect 20456 23548 20536 23576
rect 20530 23536 20536 23548
rect 20588 23536 20594 23588
rect 27540 23585 27568 23684
rect 28353 23681 28365 23684
rect 28399 23681 28411 23715
rect 28460 23712 28488 23820
rect 28537 23817 28549 23851
rect 28583 23848 28595 23851
rect 32950 23848 32956 23860
rect 28583 23820 32956 23848
rect 28583 23817 28595 23820
rect 28537 23811 28595 23817
rect 32950 23808 32956 23820
rect 33008 23808 33014 23860
rect 34149 23851 34207 23857
rect 33244 23820 34100 23848
rect 28828 23752 30604 23780
rect 28828 23712 28856 23752
rect 28460 23684 28856 23712
rect 28997 23715 29055 23721
rect 28353 23675 28411 23681
rect 28997 23681 29009 23715
rect 29043 23712 29055 23715
rect 29086 23712 29092 23724
rect 29043 23684 29092 23712
rect 29043 23681 29055 23684
rect 28997 23675 29055 23681
rect 29086 23672 29092 23684
rect 29144 23672 29150 23724
rect 29181 23715 29239 23721
rect 29181 23681 29193 23715
rect 29227 23712 29239 23715
rect 29270 23712 29276 23724
rect 29227 23684 29276 23712
rect 29227 23681 29239 23684
rect 29181 23675 29239 23681
rect 29270 23672 29276 23684
rect 29328 23672 29334 23724
rect 29914 23712 29920 23724
rect 29875 23684 29920 23712
rect 29914 23672 29920 23684
rect 29972 23712 29978 23724
rect 30282 23712 30288 23724
rect 29972 23684 30288 23712
rect 29972 23672 29978 23684
rect 30282 23672 30288 23684
rect 30340 23672 30346 23724
rect 28169 23647 28227 23653
rect 28169 23613 28181 23647
rect 28215 23644 28227 23647
rect 28810 23644 28816 23656
rect 28215 23616 28816 23644
rect 28215 23613 28227 23616
rect 28169 23607 28227 23613
rect 28810 23604 28816 23616
rect 28868 23604 28874 23656
rect 29733 23647 29791 23653
rect 29733 23613 29745 23647
rect 29779 23644 29791 23647
rect 30374 23644 30380 23656
rect 29779 23616 30380 23644
rect 29779 23613 29791 23616
rect 29733 23607 29791 23613
rect 30374 23604 30380 23616
rect 30432 23604 30438 23656
rect 30576 23653 30604 23752
rect 31938 23740 31944 23792
rect 31996 23780 32002 23792
rect 32309 23783 32367 23789
rect 32309 23780 32321 23783
rect 31996 23752 32321 23780
rect 31996 23740 32002 23752
rect 32309 23749 32321 23752
rect 32355 23780 32367 23783
rect 32355 23752 32904 23780
rect 32355 23749 32367 23752
rect 32309 23743 32367 23749
rect 30742 23712 30748 23724
rect 30703 23684 30748 23712
rect 30742 23672 30748 23684
rect 30800 23672 30806 23724
rect 30834 23672 30840 23724
rect 30892 23712 30898 23724
rect 32214 23712 32220 23724
rect 30892 23684 30937 23712
rect 32175 23684 32220 23712
rect 30892 23672 30898 23684
rect 32214 23672 32220 23684
rect 32272 23672 32278 23724
rect 32876 23721 32904 23752
rect 32401 23715 32459 23721
rect 32401 23681 32413 23715
rect 32447 23681 32459 23715
rect 32401 23675 32459 23681
rect 32861 23715 32919 23721
rect 32861 23681 32873 23715
rect 32907 23681 32919 23715
rect 33042 23712 33048 23724
rect 33003 23684 33048 23712
rect 32861 23675 32919 23681
rect 30561 23647 30619 23653
rect 30561 23613 30573 23647
rect 30607 23613 30619 23647
rect 30561 23607 30619 23613
rect 31938 23604 31944 23656
rect 31996 23644 32002 23656
rect 32306 23644 32312 23656
rect 31996 23616 32312 23644
rect 31996 23604 32002 23616
rect 32306 23604 32312 23616
rect 32364 23644 32370 23656
rect 32416 23644 32444 23675
rect 33042 23672 33048 23684
rect 33100 23672 33106 23724
rect 32364 23616 32444 23644
rect 32364 23604 32370 23616
rect 27525 23579 27583 23585
rect 27525 23545 27537 23579
rect 27571 23545 27583 23579
rect 27525 23539 27583 23545
rect 29822 23536 29828 23588
rect 29880 23576 29886 23588
rect 30101 23579 30159 23585
rect 30101 23576 30113 23579
rect 29880 23548 30113 23576
rect 29880 23536 29886 23548
rect 30101 23545 30113 23548
rect 30147 23545 30159 23579
rect 30101 23539 30159 23545
rect 30653 23579 30711 23585
rect 30653 23545 30665 23579
rect 30699 23576 30711 23579
rect 31570 23576 31576 23588
rect 30699 23548 31576 23576
rect 30699 23545 30711 23548
rect 30653 23539 30711 23545
rect 31570 23536 31576 23548
rect 31628 23536 31634 23588
rect 33244 23576 33272 23820
rect 33594 23740 33600 23792
rect 33652 23780 33658 23792
rect 33689 23783 33747 23789
rect 33689 23780 33701 23783
rect 33652 23752 33701 23780
rect 33652 23740 33658 23752
rect 33689 23749 33701 23752
rect 33735 23749 33747 23783
rect 33689 23743 33747 23749
rect 33318 23672 33324 23724
rect 33376 23712 33382 23724
rect 33965 23715 34023 23721
rect 33965 23712 33977 23715
rect 33376 23684 33977 23712
rect 33376 23672 33382 23684
rect 33965 23681 33977 23684
rect 34011 23681 34023 23715
rect 33965 23675 34023 23681
rect 33781 23647 33839 23653
rect 33781 23613 33793 23647
rect 33827 23613 33839 23647
rect 34072 23644 34100 23820
rect 34149 23817 34161 23851
rect 34195 23817 34207 23851
rect 35342 23848 35348 23860
rect 35303 23820 35348 23848
rect 34149 23811 34207 23817
rect 34164 23780 34192 23811
rect 35342 23808 35348 23820
rect 35400 23808 35406 23860
rect 40770 23848 40776 23860
rect 40731 23820 40776 23848
rect 40770 23808 40776 23820
rect 40828 23808 40834 23860
rect 40862 23808 40868 23860
rect 40920 23848 40926 23860
rect 41417 23851 41475 23857
rect 41417 23848 41429 23851
rect 40920 23820 41429 23848
rect 40920 23808 40926 23820
rect 41417 23817 41429 23820
rect 41463 23848 41475 23851
rect 42334 23848 42340 23860
rect 41463 23820 42340 23848
rect 41463 23817 41475 23820
rect 41417 23811 41475 23817
rect 42334 23808 42340 23820
rect 42392 23808 42398 23860
rect 42518 23848 42524 23860
rect 42479 23820 42524 23848
rect 42518 23808 42524 23820
rect 42576 23808 42582 23860
rect 40880 23780 40908 23808
rect 44174 23780 44180 23792
rect 34164 23752 39160 23780
rect 35342 23672 35348 23724
rect 35400 23712 35406 23724
rect 35437 23715 35495 23721
rect 35437 23712 35449 23715
rect 35400 23684 35449 23712
rect 35400 23672 35406 23684
rect 35437 23681 35449 23684
rect 35483 23681 35495 23715
rect 35437 23675 35495 23681
rect 35802 23672 35808 23724
rect 35860 23712 35866 23724
rect 36173 23715 36231 23721
rect 36173 23712 36185 23715
rect 35860 23684 36185 23712
rect 35860 23672 35866 23684
rect 36173 23681 36185 23684
rect 36219 23681 36231 23715
rect 37642 23712 37648 23724
rect 37603 23684 37648 23712
rect 36173 23675 36231 23681
rect 37642 23672 37648 23684
rect 37700 23672 37706 23724
rect 39132 23721 39160 23752
rect 39224 23752 40908 23780
rect 44135 23752 44180 23780
rect 39117 23715 39175 23721
rect 39117 23681 39129 23715
rect 39163 23681 39175 23715
rect 39117 23675 39175 23681
rect 36081 23647 36139 23653
rect 36081 23644 36093 23647
rect 34072 23616 36093 23644
rect 33781 23607 33839 23613
rect 36081 23613 36093 23616
rect 36127 23613 36139 23647
rect 37553 23647 37611 23653
rect 37553 23644 37565 23647
rect 36081 23607 36139 23613
rect 36556 23616 37565 23644
rect 32876 23548 33272 23576
rect 16482 23508 16488 23520
rect 15580 23480 16488 23508
rect 16482 23468 16488 23480
rect 16540 23468 16546 23520
rect 23477 23511 23535 23517
rect 23477 23477 23489 23511
rect 23523 23508 23535 23511
rect 23658 23508 23664 23520
rect 23523 23480 23664 23508
rect 23523 23477 23535 23480
rect 23477 23471 23535 23477
rect 23658 23468 23664 23480
rect 23716 23468 23722 23520
rect 28258 23508 28264 23520
rect 28219 23480 28264 23508
rect 28258 23468 28264 23480
rect 28316 23468 28322 23520
rect 29089 23511 29147 23517
rect 29089 23477 29101 23511
rect 29135 23508 29147 23511
rect 29914 23508 29920 23520
rect 29135 23480 29920 23508
rect 29135 23477 29147 23480
rect 29089 23471 29147 23477
rect 29914 23468 29920 23480
rect 29972 23468 29978 23520
rect 30742 23468 30748 23520
rect 30800 23508 30806 23520
rect 32876 23508 32904 23548
rect 30800 23480 32904 23508
rect 32953 23511 33011 23517
rect 30800 23468 30806 23480
rect 32953 23477 32965 23511
rect 32999 23508 33011 23511
rect 33226 23508 33232 23520
rect 32999 23480 33232 23508
rect 32999 23477 33011 23480
rect 32953 23471 33011 23477
rect 33226 23468 33232 23480
rect 33284 23468 33290 23520
rect 33686 23508 33692 23520
rect 33647 23480 33692 23508
rect 33686 23468 33692 23480
rect 33744 23468 33750 23520
rect 33796 23508 33824 23607
rect 36556 23585 36584 23616
rect 37553 23613 37565 23616
rect 37599 23613 37611 23647
rect 38654 23644 38660 23656
rect 38615 23616 38660 23644
rect 37553 23607 37611 23613
rect 38654 23604 38660 23616
rect 38712 23604 38718 23656
rect 39025 23647 39083 23653
rect 39025 23613 39037 23647
rect 39071 23644 39083 23647
rect 39224 23644 39252 23752
rect 44174 23740 44180 23752
rect 44232 23740 44238 23792
rect 44634 23740 44640 23792
rect 44692 23740 44698 23792
rect 47578 23740 47584 23792
rect 47636 23740 47642 23792
rect 39301 23715 39359 23721
rect 39301 23681 39313 23715
rect 39347 23712 39359 23715
rect 40037 23715 40095 23721
rect 40037 23712 40049 23715
rect 39347 23684 40049 23712
rect 39347 23681 39359 23684
rect 39301 23675 39359 23681
rect 40037 23681 40049 23684
rect 40083 23681 40095 23715
rect 41230 23712 41236 23724
rect 41191 23684 41236 23712
rect 40037 23675 40095 23681
rect 41230 23672 41236 23684
rect 41288 23672 41294 23724
rect 42613 23715 42671 23721
rect 42613 23681 42625 23715
rect 42659 23681 42671 23715
rect 43254 23712 43260 23724
rect 43215 23684 43260 23712
rect 42613 23675 42671 23681
rect 39758 23644 39764 23656
rect 39071 23616 39252 23644
rect 39719 23616 39764 23644
rect 39071 23613 39083 23616
rect 39025 23607 39083 23613
rect 39758 23604 39764 23616
rect 39816 23604 39822 23656
rect 42628 23644 42656 23675
rect 43254 23672 43260 23684
rect 43312 23672 43318 23724
rect 43622 23672 43628 23724
rect 43680 23712 43686 23724
rect 43901 23715 43959 23721
rect 43901 23712 43913 23715
rect 43680 23684 43913 23712
rect 43680 23672 43686 23684
rect 43901 23681 43913 23684
rect 43947 23681 43959 23715
rect 47596 23712 47624 23740
rect 47857 23715 47915 23721
rect 47857 23712 47869 23715
rect 47596 23684 47869 23712
rect 43901 23675 43959 23681
rect 47857 23681 47869 23684
rect 47903 23681 47915 23715
rect 48682 23712 48688 23724
rect 48643 23684 48688 23712
rect 47857 23675 47915 23681
rect 48682 23672 48688 23684
rect 48740 23712 48746 23724
rect 57698 23712 57704 23724
rect 48740 23684 57704 23712
rect 48740 23672 48746 23684
rect 57698 23672 57704 23684
rect 57756 23672 57762 23724
rect 42794 23644 42800 23656
rect 42628 23616 42800 23644
rect 42794 23604 42800 23616
rect 42852 23644 42858 23656
rect 44266 23644 44272 23656
rect 42852 23616 44272 23644
rect 42852 23604 42858 23616
rect 44266 23604 44272 23616
rect 44324 23604 44330 23656
rect 46014 23604 46020 23656
rect 46072 23644 46078 23656
rect 46109 23647 46167 23653
rect 46109 23644 46121 23647
rect 46072 23616 46121 23644
rect 46072 23604 46078 23616
rect 46109 23613 46121 23616
rect 46155 23613 46167 23647
rect 46109 23607 46167 23613
rect 46842 23604 46848 23656
rect 46900 23644 46906 23656
rect 47581 23647 47639 23653
rect 47581 23644 47593 23647
rect 46900 23616 47593 23644
rect 46900 23604 46906 23616
rect 47581 23613 47593 23616
rect 47627 23613 47639 23647
rect 47581 23607 47639 23613
rect 36541 23579 36599 23585
rect 36541 23545 36553 23579
rect 36587 23545 36599 23579
rect 36541 23539 36599 23545
rect 45649 23579 45707 23585
rect 45649 23545 45661 23579
rect 45695 23576 45707 23579
rect 46477 23579 46535 23585
rect 46477 23576 46489 23579
rect 45695 23548 46489 23576
rect 45695 23545 45707 23548
rect 45649 23539 45707 23545
rect 46477 23545 46489 23548
rect 46523 23576 46535 23579
rect 46934 23576 46940 23588
rect 46523 23548 46940 23576
rect 46523 23545 46535 23548
rect 46477 23539 46535 23545
rect 46934 23536 46940 23548
rect 46992 23536 46998 23588
rect 37369 23511 37427 23517
rect 37369 23508 37381 23511
rect 33796 23480 37381 23508
rect 37369 23477 37381 23480
rect 37415 23477 37427 23511
rect 37369 23471 37427 23477
rect 43441 23511 43499 23517
rect 43441 23477 43453 23511
rect 43487 23508 43499 23511
rect 44542 23508 44548 23520
rect 43487 23480 44548 23508
rect 43487 23477 43499 23480
rect 43441 23471 43499 23477
rect 44542 23468 44548 23480
rect 44600 23468 44606 23520
rect 46569 23511 46627 23517
rect 46569 23477 46581 23511
rect 46615 23508 46627 23511
rect 47394 23508 47400 23520
rect 46615 23480 47400 23508
rect 46615 23477 46627 23480
rect 46569 23471 46627 23477
rect 47394 23468 47400 23480
rect 47452 23468 47458 23520
rect 1104 23418 68816 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 65654 23418
rect 65706 23366 65718 23418
rect 65770 23366 65782 23418
rect 65834 23366 65846 23418
rect 65898 23366 65910 23418
rect 65962 23366 68816 23418
rect 1104 23344 68816 23366
rect 8294 23304 8300 23316
rect 8255 23276 8300 23304
rect 8294 23264 8300 23276
rect 8352 23264 8358 23316
rect 11146 23304 11152 23316
rect 11107 23276 11152 23304
rect 11146 23264 11152 23276
rect 11204 23264 11210 23316
rect 13998 23264 14004 23316
rect 14056 23304 14062 23316
rect 14093 23307 14151 23313
rect 14093 23304 14105 23307
rect 14056 23276 14105 23304
rect 14056 23264 14062 23276
rect 14093 23273 14105 23276
rect 14139 23273 14151 23307
rect 16758 23304 16764 23316
rect 16671 23276 16764 23304
rect 14093 23267 14151 23273
rect 16758 23264 16764 23276
rect 16816 23304 16822 23316
rect 19242 23304 19248 23316
rect 16816 23276 18184 23304
rect 19203 23276 19248 23304
rect 16816 23264 16822 23276
rect 5997 23239 6055 23245
rect 5997 23205 6009 23239
rect 6043 23236 6055 23239
rect 11422 23236 11428 23248
rect 6043 23208 11428 23236
rect 6043 23205 6055 23208
rect 5997 23199 6055 23205
rect 11422 23196 11428 23208
rect 11480 23196 11486 23248
rect 11514 23196 11520 23248
rect 11572 23236 11578 23248
rect 11572 23208 12434 23236
rect 11572 23196 11578 23208
rect 11698 23168 11704 23180
rect 11659 23140 11704 23168
rect 11698 23128 11704 23140
rect 11756 23128 11762 23180
rect 12406 23168 12434 23208
rect 17678 23196 17684 23248
rect 17736 23236 17742 23248
rect 17865 23239 17923 23245
rect 17865 23236 17877 23239
rect 17736 23208 17877 23236
rect 17736 23196 17742 23208
rect 17865 23205 17877 23208
rect 17911 23205 17923 23239
rect 18156 23236 18184 23276
rect 19242 23264 19248 23276
rect 19300 23264 19306 23316
rect 20254 23264 20260 23316
rect 20312 23304 20318 23316
rect 20441 23307 20499 23313
rect 20441 23304 20453 23307
rect 20312 23276 20453 23304
rect 20312 23264 20318 23276
rect 20441 23273 20453 23276
rect 20487 23273 20499 23307
rect 28166 23304 28172 23316
rect 20441 23267 20499 23273
rect 20548 23276 28172 23304
rect 20548 23236 20576 23276
rect 28166 23264 28172 23276
rect 28224 23264 28230 23316
rect 28905 23307 28963 23313
rect 28905 23273 28917 23307
rect 28951 23304 28963 23307
rect 29270 23304 29276 23316
rect 28951 23276 29276 23304
rect 28951 23273 28963 23276
rect 28905 23267 28963 23273
rect 29270 23264 29276 23276
rect 29328 23264 29334 23316
rect 34885 23307 34943 23313
rect 34885 23273 34897 23307
rect 34931 23304 34943 23307
rect 35434 23304 35440 23316
rect 34931 23276 35440 23304
rect 34931 23273 34943 23276
rect 34885 23267 34943 23273
rect 35434 23264 35440 23276
rect 35492 23264 35498 23316
rect 37826 23264 37832 23316
rect 37884 23304 37890 23316
rect 38102 23304 38108 23316
rect 37884 23276 38108 23304
rect 37884 23264 37890 23276
rect 38102 23264 38108 23276
rect 38160 23264 38166 23316
rect 38654 23304 38660 23316
rect 38580 23276 38660 23304
rect 18156 23208 20576 23236
rect 23201 23239 23259 23245
rect 17865 23199 17923 23205
rect 23201 23205 23213 23239
rect 23247 23236 23259 23239
rect 23382 23236 23388 23248
rect 23247 23208 23388 23236
rect 23247 23205 23259 23208
rect 23201 23199 23259 23205
rect 23382 23196 23388 23208
rect 23440 23236 23446 23248
rect 23753 23239 23811 23245
rect 23753 23236 23765 23239
rect 23440 23208 23765 23236
rect 23440 23196 23446 23208
rect 23753 23205 23765 23208
rect 23799 23205 23811 23239
rect 23753 23199 23811 23205
rect 26513 23239 26571 23245
rect 26513 23205 26525 23239
rect 26559 23236 26571 23239
rect 30834 23236 30840 23248
rect 26559 23208 30840 23236
rect 26559 23205 26571 23208
rect 26513 23199 26571 23205
rect 30834 23196 30840 23208
rect 30892 23196 30898 23248
rect 33318 23236 33324 23248
rect 33279 23208 33324 23236
rect 33318 23196 33324 23208
rect 33376 23196 33382 23248
rect 35069 23239 35127 23245
rect 35069 23205 35081 23239
rect 35115 23236 35127 23239
rect 38580 23236 38608 23276
rect 38654 23264 38660 23276
rect 38712 23264 38718 23316
rect 41230 23304 41236 23316
rect 41191 23276 41236 23304
rect 41230 23264 41236 23276
rect 41288 23264 41294 23316
rect 43254 23264 43260 23316
rect 43312 23304 43318 23316
rect 43901 23307 43959 23313
rect 43901 23304 43913 23307
rect 43312 23276 43913 23304
rect 43312 23264 43318 23276
rect 43901 23273 43913 23276
rect 43947 23273 43959 23307
rect 45646 23304 45652 23316
rect 43901 23267 43959 23273
rect 44008 23276 45652 23304
rect 40037 23239 40095 23245
rect 40037 23236 40049 23239
rect 35115 23208 40049 23236
rect 35115 23205 35127 23208
rect 35069 23199 35127 23205
rect 40037 23205 40049 23208
rect 40083 23205 40095 23239
rect 41049 23239 41107 23245
rect 41049 23236 41061 23239
rect 40037 23199 40095 23205
rect 40144 23208 41061 23236
rect 13081 23171 13139 23177
rect 13081 23168 13093 23171
rect 12406 23140 13093 23168
rect 13081 23137 13093 23140
rect 13127 23137 13139 23171
rect 14090 23168 14096 23180
rect 13081 23131 13139 23137
rect 13832 23140 14096 23168
rect 5350 23100 5356 23112
rect 5311 23072 5356 23100
rect 5350 23060 5356 23072
rect 5408 23060 5414 23112
rect 5534 23109 5540 23112
rect 5501 23103 5540 23109
rect 5501 23069 5513 23103
rect 5501 23063 5540 23069
rect 5534 23060 5540 23063
rect 5592 23060 5598 23112
rect 5718 23100 5724 23112
rect 5679 23072 5724 23100
rect 5718 23060 5724 23072
rect 5776 23060 5782 23112
rect 5810 23060 5816 23112
rect 5868 23109 5874 23112
rect 5868 23100 5876 23109
rect 12345 23103 12403 23109
rect 5868 23072 5913 23100
rect 5868 23063 5876 23072
rect 12345 23069 12357 23103
rect 12391 23100 12403 23103
rect 13832 23100 13860 23140
rect 14090 23128 14096 23140
rect 14148 23128 14154 23180
rect 14458 23128 14464 23180
rect 14516 23168 14522 23180
rect 14645 23171 14703 23177
rect 14645 23168 14657 23171
rect 14516 23140 14657 23168
rect 14516 23128 14522 23140
rect 14645 23137 14657 23140
rect 14691 23137 14703 23171
rect 14645 23131 14703 23137
rect 19518 23128 19524 23180
rect 19576 23168 19582 23180
rect 19613 23171 19671 23177
rect 19613 23168 19625 23171
rect 19576 23140 19625 23168
rect 19576 23128 19582 23140
rect 19613 23137 19625 23140
rect 19659 23168 19671 23171
rect 20162 23168 20168 23180
rect 19659 23140 20168 23168
rect 19659 23137 19671 23140
rect 19613 23131 19671 23137
rect 20162 23128 20168 23140
rect 20220 23128 20226 23180
rect 21453 23171 21511 23177
rect 21453 23137 21465 23171
rect 21499 23168 21511 23171
rect 22094 23168 22100 23180
rect 21499 23140 22100 23168
rect 21499 23137 21511 23140
rect 21453 23131 21511 23137
rect 22094 23128 22100 23140
rect 22152 23128 22158 23180
rect 30374 23128 30380 23180
rect 30432 23168 30438 23180
rect 31389 23171 31447 23177
rect 31389 23168 31401 23171
rect 30432 23140 31401 23168
rect 30432 23128 30438 23140
rect 31389 23137 31401 23140
rect 31435 23137 31447 23171
rect 31389 23131 31447 23137
rect 31570 23128 31576 23180
rect 31628 23168 31634 23180
rect 32861 23171 32919 23177
rect 32861 23168 32873 23171
rect 31628 23140 32873 23168
rect 31628 23128 31634 23140
rect 32861 23137 32873 23140
rect 32907 23137 32919 23171
rect 33873 23171 33931 23177
rect 33873 23168 33885 23171
rect 32861 23131 32919 23137
rect 32968 23140 33885 23168
rect 12391 23072 13860 23100
rect 12391 23069 12403 23072
rect 12345 23063 12403 23069
rect 5868 23060 5874 23063
rect 13906 23060 13912 23112
rect 13964 23100 13970 23112
rect 15654 23109 15660 23112
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 13964 23072 15393 23100
rect 13964 23060 13970 23072
rect 15381 23069 15393 23072
rect 15427 23069 15439 23103
rect 15648 23100 15660 23109
rect 15615 23072 15660 23100
rect 15381 23063 15439 23069
rect 15648 23063 15660 23072
rect 15654 23060 15660 23063
rect 15712 23060 15718 23112
rect 17770 23060 17776 23112
rect 17828 23100 17834 23112
rect 17865 23103 17923 23109
rect 17865 23100 17877 23103
rect 17828 23072 17877 23100
rect 17828 23060 17834 23072
rect 17865 23069 17877 23072
rect 17911 23069 17923 23103
rect 17865 23063 17923 23069
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23100 18107 23103
rect 18322 23100 18328 23112
rect 18095 23072 18328 23100
rect 18095 23069 18107 23072
rect 18049 23063 18107 23069
rect 18322 23060 18328 23072
rect 18380 23060 18386 23112
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 19392 23072 19441 23100
rect 19392 23060 19398 23072
rect 19429 23069 19441 23072
rect 19475 23069 19487 23103
rect 20806 23100 20812 23112
rect 19429 23063 19487 23069
rect 20272 23072 20812 23100
rect 5629 23035 5687 23041
rect 5629 23001 5641 23035
rect 5675 23032 5687 23035
rect 6362 23032 6368 23044
rect 5675 23004 6368 23032
rect 5675 23001 5687 23004
rect 5629 22995 5687 23001
rect 6362 22992 6368 23004
rect 6420 22992 6426 23044
rect 11517 23035 11575 23041
rect 11517 23001 11529 23035
rect 11563 23032 11575 23035
rect 12894 23032 12900 23044
rect 11563 23004 12900 23032
rect 11563 23001 11575 23004
rect 11517 22995 11575 23001
rect 12894 22992 12900 23004
rect 12952 22992 12958 23044
rect 13814 22992 13820 23044
rect 13872 23032 13878 23044
rect 14461 23035 14519 23041
rect 14461 23032 14473 23035
rect 13872 23004 14473 23032
rect 13872 22992 13878 23004
rect 14461 23001 14473 23004
rect 14507 23001 14519 23035
rect 14461 22995 14519 23001
rect 11609 22967 11667 22973
rect 11609 22933 11621 22967
rect 11655 22964 11667 22967
rect 12434 22964 12440 22976
rect 11655 22936 12440 22964
rect 11655 22933 11667 22936
rect 11609 22927 11667 22933
rect 12434 22924 12440 22936
rect 12492 22964 12498 22976
rect 13722 22964 13728 22976
rect 12492 22936 13728 22964
rect 12492 22924 12498 22936
rect 13722 22924 13728 22936
rect 13780 22924 13786 22976
rect 14550 22964 14556 22976
rect 14511 22936 14556 22964
rect 14550 22924 14556 22936
rect 14608 22924 14614 22976
rect 19444 22964 19472 23063
rect 20272 23041 20300 23072
rect 20806 23060 20812 23072
rect 20864 23060 20870 23112
rect 22830 23060 22836 23112
rect 22888 23060 22894 23112
rect 26418 23100 26424 23112
rect 26379 23072 26424 23100
rect 26418 23060 26424 23072
rect 26476 23060 26482 23112
rect 26602 23100 26608 23112
rect 26563 23072 26608 23100
rect 26602 23060 26608 23072
rect 26660 23060 26666 23112
rect 27706 23100 27712 23112
rect 27667 23072 27712 23100
rect 27706 23060 27712 23072
rect 27764 23060 27770 23112
rect 27893 23103 27951 23109
rect 27893 23069 27905 23103
rect 27939 23100 27951 23103
rect 28350 23100 28356 23112
rect 27939 23072 28356 23100
rect 27939 23069 27951 23072
rect 27893 23063 27951 23069
rect 28350 23060 28356 23072
rect 28408 23060 28414 23112
rect 29546 23100 29552 23112
rect 29507 23072 29552 23100
rect 29546 23060 29552 23072
rect 29604 23060 29610 23112
rect 29730 23109 29736 23112
rect 29697 23103 29736 23109
rect 29697 23069 29709 23103
rect 29697 23063 29736 23069
rect 29730 23060 29736 23063
rect 29788 23060 29794 23112
rect 29914 23100 29920 23112
rect 29875 23072 29920 23100
rect 29914 23060 29920 23072
rect 29972 23060 29978 23112
rect 30098 23109 30104 23112
rect 30055 23103 30104 23109
rect 30055 23069 30067 23103
rect 30101 23069 30104 23103
rect 30055 23063 30104 23069
rect 30098 23060 30104 23063
rect 30156 23060 30162 23112
rect 31478 23100 31484 23112
rect 31439 23072 31484 23100
rect 31478 23060 31484 23072
rect 31536 23060 31542 23112
rect 32766 23060 32772 23112
rect 32824 23100 32830 23112
rect 32968 23109 32996 23140
rect 33873 23137 33885 23140
rect 33919 23168 33931 23171
rect 37826 23168 37832 23180
rect 33919 23140 37832 23168
rect 33919 23137 33931 23140
rect 33873 23131 33931 23137
rect 37826 23128 37832 23140
rect 37884 23128 37890 23180
rect 38562 23128 38568 23180
rect 38620 23168 38626 23180
rect 38657 23171 38715 23177
rect 38657 23168 38669 23171
rect 38620 23140 38669 23168
rect 38620 23128 38626 23140
rect 38657 23137 38669 23140
rect 38703 23137 38715 23171
rect 38657 23131 38715 23137
rect 39022 23128 39028 23180
rect 39080 23168 39086 23180
rect 40144 23168 40172 23208
rect 41049 23205 41061 23208
rect 41095 23236 41107 23239
rect 42242 23236 42248 23248
rect 41095 23208 42248 23236
rect 41095 23205 41107 23208
rect 41049 23199 41107 23205
rect 39080 23140 40172 23168
rect 40313 23171 40371 23177
rect 39080 23128 39086 23140
rect 40313 23137 40325 23171
rect 40359 23168 40371 23171
rect 40862 23168 40868 23180
rect 40359 23140 40868 23168
rect 40359 23137 40371 23140
rect 40313 23131 40371 23137
rect 40862 23128 40868 23140
rect 40920 23128 40926 23180
rect 42076 23177 42104 23208
rect 42242 23196 42248 23208
rect 42300 23196 42306 23248
rect 42794 23236 42800 23248
rect 42755 23208 42800 23236
rect 42794 23196 42800 23208
rect 42852 23196 42858 23248
rect 43714 23196 43720 23248
rect 43772 23236 43778 23248
rect 44008 23245 44036 23276
rect 45646 23264 45652 23276
rect 45704 23264 45710 23316
rect 43993 23239 44051 23245
rect 43993 23236 44005 23239
rect 43772 23208 44005 23236
rect 43772 23196 43778 23208
rect 43993 23205 44005 23208
rect 44039 23205 44051 23239
rect 43993 23199 44051 23205
rect 46014 23196 46020 23248
rect 46072 23236 46078 23248
rect 46569 23239 46627 23245
rect 46569 23236 46581 23239
rect 46072 23208 46581 23236
rect 46072 23196 46078 23208
rect 46569 23205 46581 23208
rect 46615 23205 46627 23239
rect 46569 23199 46627 23205
rect 42061 23171 42119 23177
rect 42061 23137 42073 23171
rect 42107 23137 42119 23171
rect 42061 23131 42119 23137
rect 44361 23171 44419 23177
rect 44361 23137 44373 23171
rect 44407 23168 44419 23171
rect 45278 23168 45284 23180
rect 44407 23140 45284 23168
rect 44407 23137 44419 23140
rect 44361 23131 44419 23137
rect 45278 23128 45284 23140
rect 45336 23128 45342 23180
rect 46934 23168 46940 23180
rect 46895 23140 46940 23168
rect 46934 23128 46940 23140
rect 46992 23128 46998 23180
rect 32953 23103 33011 23109
rect 32953 23100 32965 23103
rect 32824 23072 32965 23100
rect 32824 23060 32830 23072
rect 32953 23069 32965 23072
rect 32999 23069 33011 23103
rect 32953 23063 33011 23069
rect 34514 23060 34520 23112
rect 34572 23100 34578 23112
rect 34701 23103 34759 23109
rect 34701 23100 34713 23103
rect 34572 23072 34713 23100
rect 34572 23060 34578 23072
rect 34701 23069 34713 23072
rect 34747 23069 34759 23103
rect 34701 23063 34759 23069
rect 34885 23103 34943 23109
rect 34885 23069 34897 23103
rect 34931 23100 34943 23103
rect 35526 23100 35532 23112
rect 34931 23072 35532 23100
rect 34931 23069 34943 23072
rect 34885 23063 34943 23069
rect 35526 23060 35532 23072
rect 35584 23060 35590 23112
rect 41874 23100 41880 23112
rect 41386 23072 41880 23100
rect 20530 23041 20536 23044
rect 20257 23035 20315 23041
rect 20257 23001 20269 23035
rect 20303 23001 20315 23035
rect 20257 22995 20315 23001
rect 20473 23035 20536 23041
rect 20473 23001 20485 23035
rect 20519 23001 20536 23035
rect 20473 22995 20536 23001
rect 20530 22992 20536 22995
rect 20588 22992 20594 23044
rect 20898 22992 20904 23044
rect 20956 23032 20962 23044
rect 21729 23035 21787 23041
rect 21729 23032 21741 23035
rect 20956 23004 21741 23032
rect 20956 22992 20962 23004
rect 21729 23001 21741 23004
rect 21775 23001 21787 23035
rect 23474 23032 23480 23044
rect 21729 22995 21787 23001
rect 23124 23004 23480 23032
rect 20622 22964 20628 22976
rect 19444 22936 20628 22964
rect 20622 22924 20628 22936
rect 20680 22924 20686 22976
rect 21910 22924 21916 22976
rect 21968 22964 21974 22976
rect 23124 22964 23152 23004
rect 23474 22992 23480 23004
rect 23532 22992 23538 23044
rect 26234 22992 26240 23044
rect 26292 23032 26298 23044
rect 26620 23032 26648 23060
rect 29822 23032 29828 23044
rect 26292 23004 26648 23032
rect 27356 23004 29684 23032
rect 29783 23004 29828 23032
rect 26292 22992 26298 23004
rect 27356 22976 27384 23004
rect 21968 22936 23152 22964
rect 21968 22924 21974 22936
rect 24670 22924 24676 22976
rect 24728 22964 24734 22976
rect 27157 22967 27215 22973
rect 27157 22964 27169 22967
rect 24728 22936 27169 22964
rect 24728 22924 24734 22936
rect 27157 22933 27169 22936
rect 27203 22964 27215 22967
rect 27338 22964 27344 22976
rect 27203 22936 27344 22964
rect 27203 22933 27215 22936
rect 27157 22927 27215 22933
rect 27338 22924 27344 22936
rect 27396 22924 27402 22976
rect 27798 22964 27804 22976
rect 27759 22936 27804 22964
rect 27798 22924 27804 22936
rect 27856 22924 27862 22976
rect 29656 22964 29684 23004
rect 29822 22992 29828 23004
rect 29880 22992 29886 23044
rect 31202 23032 31208 23044
rect 30024 23004 31208 23032
rect 30024 22964 30052 23004
rect 31202 22992 31208 23004
rect 31260 22992 31266 23044
rect 37921 23035 37979 23041
rect 37921 23001 37933 23035
rect 37967 23001 37979 23035
rect 40770 23032 40776 23044
rect 40731 23004 40776 23032
rect 37921 22995 37979 23001
rect 30190 22964 30196 22976
rect 29656 22936 30052 22964
rect 30151 22936 30196 22964
rect 30190 22924 30196 22936
rect 30248 22924 30254 22976
rect 31849 22967 31907 22973
rect 31849 22933 31861 22967
rect 31895 22964 31907 22967
rect 32398 22964 32404 22976
rect 31895 22936 32404 22964
rect 31895 22933 31907 22936
rect 31849 22927 31907 22933
rect 32398 22924 32404 22936
rect 32456 22924 32462 22976
rect 35526 22924 35532 22976
rect 35584 22964 35590 22976
rect 35710 22964 35716 22976
rect 35584 22936 35716 22964
rect 35584 22924 35590 22936
rect 35710 22924 35716 22936
rect 35768 22924 35774 22976
rect 37461 22967 37519 22973
rect 37461 22933 37473 22967
rect 37507 22964 37519 22967
rect 37550 22964 37556 22976
rect 37507 22936 37556 22964
rect 37507 22933 37519 22936
rect 37461 22927 37519 22933
rect 37550 22924 37556 22936
rect 37608 22964 37614 22976
rect 37936 22964 37964 22995
rect 40770 22992 40776 23004
rect 40828 23032 40834 23044
rect 41386 23032 41414 23072
rect 41874 23060 41880 23072
rect 41932 23060 41938 23112
rect 44542 23060 44548 23112
rect 44600 23100 44606 23112
rect 45741 23103 45799 23109
rect 45741 23100 45753 23103
rect 44600 23072 45753 23100
rect 44600 23060 44606 23072
rect 45741 23069 45753 23072
rect 45787 23069 45799 23103
rect 45741 23063 45799 23069
rect 45830 23060 45836 23112
rect 45888 23100 45894 23112
rect 46017 23103 46075 23109
rect 46017 23100 46029 23103
rect 45888 23072 46029 23100
rect 45888 23060 45894 23072
rect 46017 23069 46029 23072
rect 46063 23069 46075 23103
rect 47394 23100 47400 23112
rect 47355 23072 47400 23100
rect 46017 23063 46075 23069
rect 47394 23060 47400 23072
rect 47452 23060 47458 23112
rect 42610 23032 42616 23044
rect 40828 23004 41414 23032
rect 42571 23004 42616 23032
rect 40828 22992 40834 23004
rect 42610 22992 42616 23004
rect 42668 23032 42674 23044
rect 43257 23035 43315 23041
rect 43257 23032 43269 23035
rect 42668 23004 43269 23032
rect 42668 22992 42674 23004
rect 43257 23001 43269 23004
rect 43303 23001 43315 23035
rect 43257 22995 43315 23001
rect 39850 22964 39856 22976
rect 37608 22936 37964 22964
rect 39811 22936 39856 22964
rect 37608 22924 37614 22936
rect 39850 22924 39856 22936
rect 39908 22924 39914 22976
rect 39942 22924 39948 22976
rect 40000 22964 40006 22976
rect 41693 22967 41751 22973
rect 41693 22964 41705 22967
rect 40000 22936 41705 22964
rect 40000 22924 40006 22936
rect 41693 22933 41705 22936
rect 41739 22933 41751 22967
rect 41693 22927 41751 22933
rect 44174 22924 44180 22976
rect 44232 22964 44238 22976
rect 45005 22967 45063 22973
rect 45005 22964 45017 22967
rect 44232 22936 45017 22964
rect 44232 22924 44238 22936
rect 45005 22933 45017 22936
rect 45051 22933 45063 22967
rect 45005 22927 45063 22933
rect 46106 22924 46112 22976
rect 46164 22964 46170 22976
rect 46477 22967 46535 22973
rect 46477 22964 46489 22967
rect 46164 22936 46489 22964
rect 46164 22924 46170 22936
rect 46477 22933 46489 22936
rect 46523 22933 46535 22967
rect 47578 22964 47584 22976
rect 47539 22936 47584 22964
rect 46477 22927 46535 22933
rect 47578 22924 47584 22936
rect 47636 22924 47642 22976
rect 1104 22874 68816 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 68816 22874
rect 1104 22800 68816 22822
rect 5534 22760 5540 22772
rect 5495 22732 5540 22760
rect 5534 22720 5540 22732
rect 5592 22720 5598 22772
rect 6362 22760 6368 22772
rect 6323 22732 6368 22760
rect 6362 22720 6368 22732
rect 6420 22720 6426 22772
rect 10413 22763 10471 22769
rect 10413 22729 10425 22763
rect 10459 22760 10471 22763
rect 11054 22760 11060 22772
rect 10459 22732 11060 22760
rect 10459 22729 10471 22732
rect 10413 22723 10471 22729
rect 11054 22720 11060 22732
rect 11112 22720 11118 22772
rect 12437 22763 12495 22769
rect 12437 22729 12449 22763
rect 12483 22760 12495 22763
rect 12526 22760 12532 22772
rect 12483 22732 12532 22760
rect 12483 22729 12495 22732
rect 12437 22723 12495 22729
rect 12526 22720 12532 22732
rect 12584 22720 12590 22772
rect 14642 22760 14648 22772
rect 12636 22732 14648 22760
rect 5169 22695 5227 22701
rect 5169 22692 5181 22695
rect 4724 22664 5181 22692
rect 4341 22627 4399 22633
rect 4341 22593 4353 22627
rect 4387 22593 4399 22627
rect 4341 22587 4399 22593
rect 4249 22559 4307 22565
rect 4249 22525 4261 22559
rect 4295 22525 4307 22559
rect 4249 22519 4307 22525
rect 4264 22420 4292 22519
rect 4356 22488 4384 22587
rect 4724 22565 4752 22664
rect 5169 22661 5181 22664
rect 5215 22692 5227 22695
rect 5215 22664 6592 22692
rect 5215 22661 5227 22664
rect 5169 22655 5227 22661
rect 5350 22624 5356 22636
rect 5263 22596 5356 22624
rect 5350 22584 5356 22596
rect 5408 22624 5414 22636
rect 6564 22633 6592 22664
rect 6365 22627 6423 22633
rect 6365 22624 6377 22627
rect 5408 22596 6377 22624
rect 5408 22584 5414 22596
rect 6365 22593 6377 22596
rect 6411 22593 6423 22627
rect 6365 22587 6423 22593
rect 6549 22627 6607 22633
rect 6549 22593 6561 22627
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 11977 22627 12035 22633
rect 11977 22593 11989 22627
rect 12023 22624 12035 22627
rect 12434 22624 12440 22636
rect 12023 22596 12440 22624
rect 12023 22593 12035 22596
rect 11977 22587 12035 22593
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 12636 22633 12664 22732
rect 14642 22720 14648 22732
rect 14700 22720 14706 22772
rect 16758 22720 16764 22772
rect 16816 22760 16822 22772
rect 17126 22760 17132 22772
rect 16816 22732 17132 22760
rect 16816 22720 16822 22732
rect 17126 22720 17132 22732
rect 17184 22720 17190 22772
rect 17218 22720 17224 22772
rect 17276 22760 17282 22772
rect 17773 22763 17831 22769
rect 17773 22760 17785 22763
rect 17276 22732 17785 22760
rect 17276 22720 17282 22732
rect 17773 22729 17785 22732
rect 17819 22729 17831 22763
rect 17773 22723 17831 22729
rect 18414 22720 18420 22772
rect 18472 22760 18478 22772
rect 19518 22760 19524 22772
rect 18472 22732 19524 22760
rect 18472 22720 18478 22732
rect 19518 22720 19524 22732
rect 19576 22720 19582 22772
rect 23382 22720 23388 22772
rect 23440 22760 23446 22772
rect 23753 22763 23811 22769
rect 23753 22760 23765 22763
rect 23440 22732 23765 22760
rect 23440 22720 23446 22732
rect 23753 22729 23765 22732
rect 23799 22729 23811 22763
rect 23753 22723 23811 22729
rect 25777 22763 25835 22769
rect 25777 22729 25789 22763
rect 25823 22760 25835 22763
rect 25866 22760 25872 22772
rect 25823 22732 25872 22760
rect 25823 22729 25835 22732
rect 25777 22723 25835 22729
rect 25866 22720 25872 22732
rect 25924 22760 25930 22772
rect 26786 22760 26792 22772
rect 25924 22732 26792 22760
rect 25924 22720 25930 22732
rect 26786 22720 26792 22732
rect 26844 22720 26850 22772
rect 26973 22763 27031 22769
rect 26973 22729 26985 22763
rect 27019 22729 27031 22763
rect 27338 22760 27344 22772
rect 27299 22732 27344 22760
rect 26973 22723 27031 22729
rect 13078 22692 13084 22704
rect 13039 22664 13084 22692
rect 13078 22652 13084 22664
rect 13136 22652 13142 22704
rect 14550 22652 14556 22704
rect 14608 22692 14614 22704
rect 15013 22695 15071 22701
rect 15013 22692 15025 22695
rect 14608 22664 15025 22692
rect 14608 22652 14614 22664
rect 15013 22661 15025 22664
rect 15059 22692 15071 22695
rect 16117 22695 16175 22701
rect 16117 22692 16129 22695
rect 15059 22664 16129 22692
rect 15059 22661 15071 22664
rect 15013 22655 15071 22661
rect 16117 22661 16129 22664
rect 16163 22692 16175 22695
rect 17037 22695 17095 22701
rect 17037 22692 17049 22695
rect 16163 22664 17049 22692
rect 16163 22661 16175 22664
rect 16117 22655 16175 22661
rect 17037 22661 17049 22664
rect 17083 22692 17095 22695
rect 18598 22692 18604 22704
rect 17083 22664 18604 22692
rect 17083 22661 17095 22664
rect 17037 22655 17095 22661
rect 18598 22652 18604 22664
rect 18656 22652 18662 22704
rect 20254 22652 20260 22704
rect 20312 22692 20318 22704
rect 20625 22695 20683 22701
rect 20625 22692 20637 22695
rect 20312 22664 20637 22692
rect 20312 22652 20318 22664
rect 20625 22661 20637 22664
rect 20671 22661 20683 22695
rect 20625 22655 20683 22661
rect 12621 22627 12679 22633
rect 12621 22593 12633 22627
rect 12667 22593 12679 22627
rect 12621 22587 12679 22593
rect 12713 22627 12771 22633
rect 12713 22593 12725 22627
rect 12759 22624 12771 22627
rect 12894 22624 12900 22636
rect 12759 22596 12900 22624
rect 12759 22593 12771 22596
rect 12713 22587 12771 22593
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 13817 22627 13875 22633
rect 13817 22593 13829 22627
rect 13863 22624 13875 22627
rect 14182 22624 14188 22636
rect 13863 22596 14188 22624
rect 13863 22593 13875 22596
rect 13817 22587 13875 22593
rect 14182 22584 14188 22596
rect 14240 22584 14246 22636
rect 17681 22627 17739 22633
rect 17681 22593 17693 22627
rect 17727 22593 17739 22627
rect 17954 22624 17960 22636
rect 17915 22596 17960 22624
rect 17681 22587 17739 22593
rect 4709 22559 4767 22565
rect 4709 22525 4721 22559
rect 4755 22525 4767 22559
rect 4709 22519 4767 22525
rect 12989 22559 13047 22565
rect 12989 22525 13001 22559
rect 13035 22525 13047 22559
rect 17696 22556 17724 22587
rect 17954 22584 17960 22596
rect 18012 22584 18018 22636
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22624 18475 22627
rect 18690 22624 18696 22636
rect 18463 22596 18696 22624
rect 18463 22593 18475 22596
rect 18417 22587 18475 22593
rect 18690 22584 18696 22596
rect 18748 22584 18754 22636
rect 19613 22627 19671 22633
rect 19613 22593 19625 22627
rect 19659 22624 19671 22627
rect 20162 22624 20168 22636
rect 19659 22596 20168 22624
rect 19659 22593 19671 22596
rect 19613 22587 19671 22593
rect 20162 22584 20168 22596
rect 20220 22584 20226 22636
rect 20530 22624 20536 22636
rect 20491 22596 20536 22624
rect 20530 22584 20536 22596
rect 20588 22584 20594 22636
rect 20806 22624 20812 22636
rect 20767 22596 20812 22624
rect 20806 22584 20812 22596
rect 20864 22584 20870 22636
rect 21542 22584 21548 22636
rect 21600 22624 21606 22636
rect 22629 22627 22687 22633
rect 22629 22624 22641 22627
rect 21600 22596 22641 22624
rect 21600 22584 21606 22596
rect 22629 22593 22641 22596
rect 22675 22593 22687 22627
rect 22629 22587 22687 22593
rect 24581 22627 24639 22633
rect 24581 22593 24593 22627
rect 24627 22624 24639 22627
rect 26421 22627 26479 22633
rect 24627 22596 25176 22624
rect 24627 22593 24639 22596
rect 24581 22587 24639 22593
rect 18046 22556 18052 22568
rect 17696 22528 18052 22556
rect 12989 22519 13047 22525
rect 5902 22488 5908 22500
rect 4356 22460 5908 22488
rect 5902 22448 5908 22460
rect 5960 22448 5966 22500
rect 7926 22420 7932 22432
rect 4264 22392 7932 22420
rect 7926 22380 7932 22392
rect 7984 22380 7990 22432
rect 13004 22420 13032 22519
rect 18046 22516 18052 22528
rect 18104 22516 18110 22568
rect 22094 22516 22100 22568
rect 22152 22556 22158 22568
rect 22278 22556 22284 22568
rect 22152 22528 22284 22556
rect 22152 22516 22158 22528
rect 22278 22516 22284 22528
rect 22336 22556 22342 22568
rect 22373 22559 22431 22565
rect 22373 22556 22385 22559
rect 22336 22528 22385 22556
rect 22336 22516 22342 22528
rect 22373 22525 22385 22528
rect 22419 22525 22431 22559
rect 22373 22519 22431 22525
rect 25148 22500 25176 22596
rect 26421 22593 26433 22627
rect 26467 22624 26479 22627
rect 26988 22624 27016 22723
rect 27338 22720 27344 22732
rect 27396 22720 27402 22772
rect 27430 22720 27436 22772
rect 27488 22760 27494 22772
rect 30009 22763 30067 22769
rect 27488 22732 27660 22760
rect 27488 22720 27494 22732
rect 26467 22596 27016 22624
rect 27264 22664 27476 22692
rect 26467 22593 26479 22596
rect 26421 22587 26479 22593
rect 26786 22516 26792 22568
rect 26844 22556 26850 22568
rect 27264 22556 27292 22664
rect 27448 22624 27476 22664
rect 27448 22596 27568 22624
rect 27540 22565 27568 22596
rect 26844 22528 27292 22556
rect 27525 22559 27583 22565
rect 26844 22516 26850 22528
rect 27525 22525 27537 22559
rect 27571 22525 27583 22559
rect 27525 22519 27583 22525
rect 13998 22488 14004 22500
rect 13959 22460 14004 22488
rect 13998 22448 14004 22460
rect 14056 22448 14062 22500
rect 17770 22448 17776 22500
rect 17828 22488 17834 22500
rect 17957 22491 18015 22497
rect 17957 22488 17969 22491
rect 17828 22460 17969 22488
rect 17828 22448 17834 22460
rect 17957 22457 17969 22460
rect 18003 22457 18015 22491
rect 18874 22488 18880 22500
rect 17957 22451 18015 22457
rect 18340 22460 18880 22488
rect 18340 22420 18368 22460
rect 18874 22448 18880 22460
rect 18932 22448 18938 22500
rect 23474 22448 23480 22500
rect 23532 22488 23538 22500
rect 24397 22491 24455 22497
rect 24397 22488 24409 22491
rect 23532 22460 24409 22488
rect 23532 22448 23538 22460
rect 24397 22457 24409 22460
rect 24443 22457 24455 22491
rect 25130 22488 25136 22500
rect 25091 22460 25136 22488
rect 24397 22451 24455 22457
rect 25130 22448 25136 22460
rect 25188 22448 25194 22500
rect 27632 22488 27660 22732
rect 30009 22729 30021 22763
rect 30055 22760 30067 22763
rect 30282 22760 30288 22772
rect 30055 22732 30288 22760
rect 30055 22729 30067 22732
rect 30009 22723 30067 22729
rect 30282 22720 30288 22732
rect 30340 22720 30346 22772
rect 31573 22763 31631 22769
rect 31573 22729 31585 22763
rect 31619 22760 31631 22763
rect 31938 22760 31944 22772
rect 31619 22732 31944 22760
rect 31619 22729 31631 22732
rect 31573 22723 31631 22729
rect 31938 22720 31944 22732
rect 31996 22720 32002 22772
rect 32125 22763 32183 22769
rect 32125 22729 32137 22763
rect 32171 22760 32183 22763
rect 32214 22760 32220 22772
rect 32171 22732 32220 22760
rect 32171 22729 32183 22732
rect 32125 22723 32183 22729
rect 32214 22720 32220 22732
rect 32272 22720 32278 22772
rect 33597 22763 33655 22769
rect 33597 22729 33609 22763
rect 33643 22729 33655 22763
rect 35434 22760 35440 22772
rect 35395 22732 35440 22760
rect 33597 22723 33655 22729
rect 27798 22652 27804 22704
rect 27856 22692 27862 22704
rect 33137 22695 33195 22701
rect 33137 22692 33149 22695
rect 27856 22664 33149 22692
rect 27856 22652 27862 22664
rect 33137 22661 33149 22664
rect 33183 22661 33195 22695
rect 33612 22692 33640 22723
rect 35434 22720 35440 22732
rect 35492 22720 35498 22772
rect 45649 22763 45707 22769
rect 36004 22732 41414 22760
rect 36004 22692 36032 22732
rect 33612 22664 36032 22692
rect 36081 22695 36139 22701
rect 33137 22655 33195 22661
rect 36081 22661 36093 22695
rect 36127 22692 36139 22695
rect 40770 22692 40776 22704
rect 36127 22664 40776 22692
rect 36127 22661 36139 22664
rect 36081 22655 36139 22661
rect 40770 22652 40776 22664
rect 40828 22652 40834 22704
rect 41386 22692 41414 22732
rect 45649 22729 45661 22763
rect 45695 22760 45707 22763
rect 46014 22760 46020 22772
rect 45695 22732 46020 22760
rect 45695 22729 45707 22732
rect 45649 22723 45707 22729
rect 46014 22720 46020 22732
rect 46072 22720 46078 22772
rect 43714 22692 43720 22704
rect 41386 22664 43720 22692
rect 43714 22652 43720 22664
rect 43772 22652 43778 22704
rect 44174 22692 44180 22704
rect 44135 22664 44180 22692
rect 44174 22652 44180 22664
rect 44232 22652 44238 22704
rect 45462 22692 45468 22704
rect 45402 22664 45468 22692
rect 45462 22652 45468 22664
rect 45520 22652 45526 22704
rect 29914 22624 29920 22636
rect 29875 22596 29920 22624
rect 29914 22584 29920 22596
rect 29972 22584 29978 22636
rect 30098 22584 30104 22636
rect 30156 22624 30162 22636
rect 30193 22627 30251 22633
rect 30193 22624 30205 22627
rect 30156 22596 30205 22624
rect 30156 22584 30162 22596
rect 30193 22593 30205 22596
rect 30239 22593 30251 22627
rect 30193 22587 30251 22593
rect 31754 22584 31760 22636
rect 31812 22624 31818 22636
rect 32585 22627 32643 22633
rect 32585 22624 32597 22627
rect 31812 22596 32597 22624
rect 31812 22584 31818 22596
rect 32585 22593 32597 22596
rect 32631 22593 32643 22627
rect 33410 22624 33416 22636
rect 33371 22596 33416 22624
rect 32585 22587 32643 22593
rect 33410 22584 33416 22596
rect 33468 22584 33474 22636
rect 35621 22627 35679 22633
rect 35621 22624 35633 22627
rect 34900 22596 35633 22624
rect 29932 22556 29960 22584
rect 30282 22556 30288 22568
rect 29932 22528 30288 22556
rect 30282 22516 30288 22528
rect 30340 22516 30346 22568
rect 31113 22559 31171 22565
rect 31113 22525 31125 22559
rect 31159 22556 31171 22559
rect 33226 22556 33232 22568
rect 31159 22528 31754 22556
rect 33187 22528 33232 22556
rect 31159 22525 31171 22528
rect 31113 22519 31171 22525
rect 31128 22488 31156 22519
rect 31478 22488 31484 22500
rect 27632 22460 31156 22488
rect 31439 22460 31484 22488
rect 31478 22448 31484 22460
rect 31536 22448 31542 22500
rect 31726 22488 31754 22528
rect 33226 22516 33232 22528
rect 33284 22516 33290 22568
rect 32217 22491 32275 22497
rect 32217 22488 32229 22491
rect 31726 22460 32229 22488
rect 32217 22457 32229 22460
rect 32263 22457 32275 22491
rect 34698 22488 34704 22500
rect 32217 22451 32275 22457
rect 33428 22460 34704 22488
rect 18506 22420 18512 22432
rect 13004 22392 18368 22420
rect 18467 22392 18512 22420
rect 18506 22380 18512 22392
rect 18564 22380 18570 22432
rect 20809 22423 20867 22429
rect 20809 22389 20821 22423
rect 20855 22420 20867 22423
rect 21082 22420 21088 22432
rect 20855 22392 21088 22420
rect 20855 22389 20867 22392
rect 20809 22383 20867 22389
rect 21082 22380 21088 22392
rect 21140 22380 21146 22432
rect 26237 22423 26295 22429
rect 26237 22389 26249 22423
rect 26283 22420 26295 22423
rect 26326 22420 26332 22432
rect 26283 22392 26332 22420
rect 26283 22389 26295 22392
rect 26237 22383 26295 22389
rect 26326 22380 26332 22392
rect 26384 22380 26390 22432
rect 30377 22423 30435 22429
rect 30377 22389 30389 22423
rect 30423 22420 30435 22423
rect 32122 22420 32128 22432
rect 30423 22392 32128 22420
rect 30423 22389 30435 22392
rect 30377 22383 30435 22389
rect 32122 22380 32128 22392
rect 32180 22380 32186 22432
rect 33428 22429 33456 22460
rect 34698 22448 34704 22460
rect 34756 22448 34762 22500
rect 33413 22423 33471 22429
rect 33413 22389 33425 22423
rect 33459 22389 33471 22423
rect 33413 22383 33471 22389
rect 34790 22380 34796 22432
rect 34848 22420 34854 22432
rect 34900 22429 34928 22596
rect 35621 22593 35633 22596
rect 35667 22593 35679 22627
rect 35621 22587 35679 22593
rect 35805 22627 35863 22633
rect 35805 22593 35817 22627
rect 35851 22624 35863 22627
rect 39022 22624 39028 22636
rect 35851 22596 39028 22624
rect 35851 22593 35863 22596
rect 35805 22587 35863 22593
rect 39022 22584 39028 22596
rect 39080 22584 39086 22636
rect 39117 22627 39175 22633
rect 39117 22593 39129 22627
rect 39163 22624 39175 22627
rect 39942 22624 39948 22636
rect 39163 22596 39948 22624
rect 39163 22593 39175 22596
rect 39117 22587 39175 22593
rect 39942 22584 39948 22596
rect 40000 22584 40006 22636
rect 40034 22584 40040 22636
rect 40092 22624 40098 22636
rect 40497 22627 40555 22633
rect 40497 22624 40509 22627
rect 40092 22596 40509 22624
rect 40092 22584 40098 22596
rect 40497 22593 40509 22596
rect 40543 22593 40555 22627
rect 40497 22587 40555 22593
rect 43622 22584 43628 22636
rect 43680 22624 43686 22636
rect 43901 22627 43959 22633
rect 43901 22624 43913 22627
rect 43680 22596 43913 22624
rect 43680 22584 43686 22596
rect 43901 22593 43913 22596
rect 43947 22593 43959 22627
rect 46106 22624 46112 22636
rect 46067 22596 46112 22624
rect 43901 22587 43959 22593
rect 46106 22584 46112 22596
rect 46164 22584 46170 22636
rect 46293 22627 46351 22633
rect 46293 22593 46305 22627
rect 46339 22624 46351 22627
rect 47578 22624 47584 22636
rect 46339 22596 47584 22624
rect 46339 22593 46351 22596
rect 46293 22587 46351 22593
rect 39758 22516 39764 22568
rect 39816 22556 39822 22568
rect 40221 22559 40279 22565
rect 40221 22556 40233 22559
rect 39816 22528 40233 22556
rect 39816 22516 39822 22528
rect 40221 22525 40233 22528
rect 40267 22525 40279 22559
rect 40221 22519 40279 22525
rect 45370 22516 45376 22568
rect 45428 22556 45434 22568
rect 46308 22556 46336 22587
rect 47578 22584 47584 22596
rect 47636 22584 47642 22636
rect 45428 22528 46336 22556
rect 45428 22516 45434 22528
rect 39301 22491 39359 22497
rect 39301 22457 39313 22491
rect 39347 22488 39359 22491
rect 39776 22488 39804 22516
rect 39347 22460 39804 22488
rect 39347 22457 39359 22460
rect 39301 22451 39359 22457
rect 34885 22423 34943 22429
rect 34885 22420 34897 22423
rect 34848 22392 34897 22420
rect 34848 22380 34854 22392
rect 34885 22389 34897 22392
rect 34931 22389 34943 22423
rect 35802 22420 35808 22432
rect 35763 22392 35808 22420
rect 34885 22383 34943 22389
rect 35802 22380 35808 22392
rect 35860 22380 35866 22432
rect 41230 22420 41236 22432
rect 41191 22392 41236 22420
rect 41230 22380 41236 22392
rect 41288 22380 41294 22432
rect 46014 22380 46020 22432
rect 46072 22420 46078 22432
rect 46109 22423 46167 22429
rect 46109 22420 46121 22423
rect 46072 22392 46121 22420
rect 46072 22380 46078 22392
rect 46109 22389 46121 22392
rect 46155 22389 46167 22423
rect 46109 22383 46167 22389
rect 1104 22330 68816 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 65654 22330
rect 65706 22278 65718 22330
rect 65770 22278 65782 22330
rect 65834 22278 65846 22330
rect 65898 22278 65910 22330
rect 65962 22278 68816 22330
rect 1104 22256 68816 22278
rect 4341 22219 4399 22225
rect 4341 22185 4353 22219
rect 4387 22216 4399 22219
rect 5350 22216 5356 22228
rect 4387 22188 5356 22216
rect 4387 22185 4399 22188
rect 4341 22179 4399 22185
rect 5350 22176 5356 22188
rect 5408 22176 5414 22228
rect 10686 22176 10692 22228
rect 10744 22216 10750 22228
rect 10781 22219 10839 22225
rect 10781 22216 10793 22219
rect 10744 22188 10793 22216
rect 10744 22176 10750 22188
rect 10781 22185 10793 22188
rect 10827 22216 10839 22219
rect 11054 22216 11060 22228
rect 10827 22188 11060 22216
rect 10827 22185 10839 22188
rect 10781 22179 10839 22185
rect 11054 22176 11060 22188
rect 11112 22176 11118 22228
rect 17218 22176 17224 22228
rect 17276 22216 17282 22228
rect 17957 22219 18015 22225
rect 17957 22216 17969 22219
rect 17276 22188 17969 22216
rect 17276 22176 17282 22188
rect 17957 22185 17969 22188
rect 18003 22185 18015 22219
rect 20898 22216 20904 22228
rect 20859 22188 20904 22216
rect 17957 22179 18015 22185
rect 20898 22176 20904 22188
rect 20956 22176 20962 22228
rect 21542 22216 21548 22228
rect 21503 22188 21548 22216
rect 21542 22176 21548 22188
rect 21600 22176 21606 22228
rect 24302 22176 24308 22228
rect 24360 22216 24366 22228
rect 25225 22219 25283 22225
rect 25225 22216 25237 22219
rect 24360 22188 25237 22216
rect 24360 22176 24366 22188
rect 25225 22185 25237 22188
rect 25271 22216 25283 22219
rect 27430 22216 27436 22228
rect 25271 22188 27292 22216
rect 27391 22188 27436 22216
rect 25271 22185 25283 22188
rect 25225 22179 25283 22185
rect 13998 22108 14004 22160
rect 14056 22148 14062 22160
rect 15378 22148 15384 22160
rect 14056 22120 15384 22148
rect 14056 22108 14062 22120
rect 15378 22108 15384 22120
rect 15436 22108 15442 22160
rect 16482 22148 16488 22160
rect 16132 22120 16488 22148
rect 5721 22083 5779 22089
rect 5721 22049 5733 22083
rect 5767 22080 5779 22083
rect 6638 22080 6644 22092
rect 5767 22052 6644 22080
rect 5767 22049 5779 22052
rect 5721 22043 5779 22049
rect 6638 22040 6644 22052
rect 6696 22080 6702 22092
rect 11514 22080 11520 22092
rect 6696 22052 11520 22080
rect 6696 22040 6702 22052
rect 11514 22040 11520 22052
rect 11572 22040 11578 22092
rect 11606 22040 11612 22092
rect 11664 22080 11670 22092
rect 13814 22080 13820 22092
rect 11664 22052 13820 22080
rect 11664 22040 11670 22052
rect 13814 22040 13820 22052
rect 13872 22040 13878 22092
rect 16132 22089 16160 22120
rect 16482 22108 16488 22120
rect 16540 22108 16546 22160
rect 16758 22108 16764 22160
rect 16816 22148 16822 22160
rect 20714 22148 20720 22160
rect 16816 22120 20720 22148
rect 16816 22108 16822 22120
rect 20714 22108 20720 22120
rect 20772 22108 20778 22160
rect 27264 22148 27292 22188
rect 27430 22176 27436 22188
rect 27488 22176 27494 22228
rect 32493 22219 32551 22225
rect 32493 22185 32505 22219
rect 32539 22216 32551 22219
rect 33686 22216 33692 22228
rect 32539 22188 33692 22216
rect 32539 22185 32551 22188
rect 32493 22179 32551 22185
rect 33686 22176 33692 22188
rect 33744 22176 33750 22228
rect 34698 22216 34704 22228
rect 34659 22188 34704 22216
rect 34698 22176 34704 22188
rect 34756 22176 34762 22228
rect 34882 22216 34888 22228
rect 34843 22188 34888 22216
rect 34882 22176 34888 22188
rect 34940 22176 34946 22228
rect 40034 22216 40040 22228
rect 39995 22188 40040 22216
rect 40034 22176 40040 22188
rect 40092 22176 40098 22228
rect 40852 22219 40910 22225
rect 40852 22185 40864 22219
rect 40898 22216 40910 22219
rect 41230 22216 41236 22228
rect 40898 22188 41236 22216
rect 40898 22185 40910 22188
rect 40852 22179 40910 22185
rect 41230 22176 41236 22188
rect 41288 22176 41294 22228
rect 41874 22176 41880 22228
rect 41932 22216 41938 22228
rect 42337 22219 42395 22225
rect 42337 22216 42349 22219
rect 41932 22188 42349 22216
rect 41932 22176 41938 22188
rect 42337 22185 42349 22188
rect 42383 22185 42395 22219
rect 42337 22179 42395 22185
rect 36265 22151 36323 22157
rect 27264 22120 30972 22148
rect 16117 22083 16175 22089
rect 16117 22049 16129 22083
rect 16163 22080 16175 22083
rect 17954 22080 17960 22092
rect 16163 22052 16197 22080
rect 17788 22052 17960 22080
rect 16163 22049 16175 22052
rect 16117 22043 16175 22049
rect 5810 21972 5816 22024
rect 5868 22012 5874 22024
rect 6365 22015 6423 22021
rect 6365 22012 6377 22015
rect 5868 21984 6377 22012
rect 5868 21972 5874 21984
rect 6365 21981 6377 21984
rect 6411 21981 6423 22015
rect 10042 22012 10048 22024
rect 10003 21984 10048 22012
rect 6365 21975 6423 21981
rect 10042 21972 10048 21984
rect 10100 21972 10106 22024
rect 10226 21972 10232 22024
rect 10284 22012 10290 22024
rect 10686 22012 10692 22024
rect 10284 21984 10692 22012
rect 10284 21972 10290 21984
rect 10686 21972 10692 21984
rect 10744 21972 10750 22024
rect 12526 22012 12532 22024
rect 12487 21984 12532 22012
rect 12526 21972 12532 21984
rect 12584 21972 12590 22024
rect 12713 22015 12771 22021
rect 12713 21981 12725 22015
rect 12759 22012 12771 22015
rect 16850 22012 16856 22024
rect 12759 21984 16856 22012
rect 12759 21981 12771 21984
rect 12713 21975 12771 21981
rect 16850 21972 16856 21984
rect 16908 21972 16914 22024
rect 5476 21947 5534 21953
rect 5476 21913 5488 21947
rect 5522 21944 5534 21947
rect 5522 21916 6224 21944
rect 5522 21913 5534 21916
rect 5476 21907 5534 21913
rect 6196 21885 6224 21916
rect 8202 21904 8208 21956
rect 8260 21944 8266 21956
rect 12621 21947 12679 21953
rect 12621 21944 12633 21947
rect 8260 21916 12633 21944
rect 8260 21904 8266 21916
rect 12621 21913 12633 21916
rect 12667 21913 12679 21947
rect 12621 21907 12679 21913
rect 16301 21947 16359 21953
rect 16301 21913 16313 21947
rect 16347 21944 16359 21947
rect 16942 21944 16948 21956
rect 16347 21916 16948 21944
rect 16347 21913 16359 21916
rect 16301 21907 16359 21913
rect 16942 21904 16948 21916
rect 17000 21904 17006 21956
rect 17788 21953 17816 22052
rect 17954 22040 17960 22052
rect 18012 22040 18018 22092
rect 18046 22040 18052 22092
rect 18104 22040 18110 22092
rect 19889 22083 19947 22089
rect 19889 22049 19901 22083
rect 19935 22080 19947 22083
rect 19935 22052 22232 22080
rect 19935 22049 19947 22052
rect 19889 22043 19947 22049
rect 17773 21947 17831 21953
rect 17773 21913 17785 21947
rect 17819 21913 17831 21947
rect 17773 21907 17831 21913
rect 17973 21947 18031 21953
rect 17973 21913 17985 21947
rect 18019 21944 18031 21947
rect 18064 21944 18092 22040
rect 20622 21972 20628 22024
rect 20680 22012 20686 22024
rect 20717 22015 20775 22021
rect 20717 22012 20729 22015
rect 20680 21984 20729 22012
rect 20680 21972 20686 21984
rect 20717 21981 20729 21984
rect 20763 21981 20775 22015
rect 20717 21975 20775 21981
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 22012 20959 22015
rect 21082 22012 21088 22024
rect 20947 21984 21088 22012
rect 20947 21981 20959 21984
rect 20901 21975 20959 21981
rect 21082 21972 21088 21984
rect 21140 21972 21146 22024
rect 21266 21972 21272 22024
rect 21324 22012 21330 22024
rect 21361 22015 21419 22021
rect 21361 22012 21373 22015
rect 21324 21984 21373 22012
rect 21324 21972 21330 21984
rect 21361 21981 21373 21984
rect 21407 21981 21419 22015
rect 21361 21975 21419 21981
rect 21450 21972 21456 22024
rect 21508 22012 21514 22024
rect 22005 22015 22063 22021
rect 22005 22012 22017 22015
rect 21508 21984 22017 22012
rect 21508 21972 21514 21984
rect 22005 21981 22017 21984
rect 22051 21981 22063 22015
rect 22204 22012 22232 22052
rect 22278 22040 22284 22092
rect 22336 22080 22342 22092
rect 24394 22080 24400 22092
rect 22336 22052 24400 22080
rect 22336 22040 22342 22052
rect 24394 22040 24400 22052
rect 24452 22080 24458 22092
rect 26053 22083 26111 22089
rect 26053 22080 26065 22083
rect 24452 22052 26065 22080
rect 24452 22040 24458 22052
rect 26053 22049 26065 22052
rect 26099 22049 26111 22083
rect 26053 22043 26111 22049
rect 29362 22040 29368 22092
rect 29420 22080 29426 22092
rect 29549 22083 29607 22089
rect 29549 22080 29561 22083
rect 29420 22052 29561 22080
rect 29420 22040 29426 22052
rect 29549 22049 29561 22052
rect 29595 22049 29607 22083
rect 29914 22080 29920 22092
rect 29875 22052 29920 22080
rect 29549 22043 29607 22049
rect 29914 22040 29920 22052
rect 29972 22040 29978 22092
rect 30009 22083 30067 22089
rect 30009 22049 30021 22083
rect 30055 22080 30067 22083
rect 30190 22080 30196 22092
rect 30055 22052 30196 22080
rect 30055 22049 30067 22052
rect 30009 22043 30067 22049
rect 30190 22040 30196 22052
rect 30248 22040 30254 22092
rect 30944 22089 30972 22120
rect 36265 22117 36277 22151
rect 36311 22148 36323 22151
rect 36817 22151 36875 22157
rect 36817 22148 36829 22151
rect 36311 22120 36829 22148
rect 36311 22117 36323 22120
rect 36265 22111 36323 22117
rect 36817 22117 36829 22120
rect 36863 22117 36875 22151
rect 36817 22111 36875 22117
rect 40420 22120 40724 22148
rect 30929 22083 30987 22089
rect 30929 22049 30941 22083
rect 30975 22080 30987 22083
rect 31478 22080 31484 22092
rect 30975 22052 31484 22080
rect 30975 22049 30987 22052
rect 30929 22043 30987 22049
rect 31478 22040 31484 22052
rect 31536 22080 31542 22092
rect 36280 22080 36308 22111
rect 31536 22052 36308 22080
rect 36357 22083 36415 22089
rect 31536 22040 31542 22052
rect 36357 22049 36369 22083
rect 36403 22049 36415 22083
rect 36357 22043 36415 22049
rect 22830 22012 22836 22024
rect 22204 21984 22324 22012
rect 22791 21984 22836 22012
rect 22005 21975 22063 21981
rect 19705 21947 19763 21953
rect 19705 21944 19717 21947
rect 18019 21916 18092 21944
rect 18616 21916 19717 21944
rect 18019 21913 18031 21916
rect 17973 21907 18031 21913
rect 18616 21888 18644 21916
rect 19705 21913 19717 21916
rect 19751 21913 19763 21947
rect 22186 21944 22192 21956
rect 22147 21916 22192 21944
rect 19705 21907 19763 21913
rect 22186 21904 22192 21916
rect 22244 21904 22250 21956
rect 22296 21944 22324 21984
rect 22830 21972 22836 21984
rect 22888 21972 22894 22024
rect 22925 22015 22983 22021
rect 22925 21981 22937 22015
rect 22971 22012 22983 22015
rect 23474 22012 23480 22024
rect 22971 21984 23480 22012
rect 22971 21981 22983 21984
rect 22925 21975 22983 21981
rect 23474 21972 23480 21984
rect 23532 21972 23538 22024
rect 24486 21972 24492 22024
rect 24544 22012 24550 22024
rect 26326 22021 26332 22024
rect 25133 22015 25191 22021
rect 25133 22012 25145 22015
rect 24544 21984 25145 22012
rect 24544 21972 24550 21984
rect 25133 21981 25145 21984
rect 25179 21981 25191 22015
rect 25133 21975 25191 21981
rect 26320 21975 26332 22021
rect 26384 22012 26390 22024
rect 26384 21984 26420 22012
rect 26326 21972 26332 21975
rect 26384 21972 26390 21984
rect 29638 21972 29644 22024
rect 29696 22012 29702 22024
rect 29733 22015 29791 22021
rect 29733 22012 29745 22015
rect 29696 21984 29745 22012
rect 29696 21972 29702 21984
rect 29733 21981 29745 21984
rect 29779 21981 29791 22015
rect 29733 21975 29791 21981
rect 29822 21972 29828 22024
rect 29880 22012 29886 22024
rect 31938 22012 31944 22024
rect 29880 21984 29925 22012
rect 31899 21984 31944 22012
rect 29880 21972 29886 21984
rect 31938 21972 31944 21984
rect 31996 21972 32002 22024
rect 32033 22015 32091 22021
rect 32033 21981 32045 22015
rect 32079 21981 32091 22015
rect 32214 22012 32220 22024
rect 32175 21984 32220 22012
rect 32033 21975 32091 21981
rect 24670 21944 24676 21956
rect 22296 21916 24676 21944
rect 24670 21904 24676 21916
rect 24728 21904 24734 21956
rect 25498 21904 25504 21956
rect 25556 21944 25562 21956
rect 31481 21947 31539 21953
rect 25556 21916 26556 21944
rect 25556 21904 25562 21916
rect 6181 21879 6239 21885
rect 6181 21845 6193 21879
rect 6227 21845 6239 21879
rect 6181 21839 6239 21845
rect 9766 21836 9772 21888
rect 9824 21876 9830 21888
rect 10137 21879 10195 21885
rect 10137 21876 10149 21879
rect 9824 21848 10149 21876
rect 9824 21836 9830 21848
rect 10137 21845 10149 21848
rect 10183 21845 10195 21879
rect 14182 21876 14188 21888
rect 14143 21848 14188 21876
rect 10137 21839 10195 21845
rect 14182 21836 14188 21848
rect 14240 21836 14246 21888
rect 15102 21836 15108 21888
rect 15160 21876 15166 21888
rect 15565 21879 15623 21885
rect 15565 21876 15577 21879
rect 15160 21848 15577 21876
rect 15160 21836 15166 21848
rect 15565 21845 15577 21848
rect 15611 21876 15623 21879
rect 16393 21879 16451 21885
rect 16393 21876 16405 21879
rect 15611 21848 16405 21876
rect 15611 21845 15623 21848
rect 15565 21839 15623 21845
rect 16393 21845 16405 21848
rect 16439 21845 16451 21879
rect 16758 21876 16764 21888
rect 16719 21848 16764 21876
rect 16393 21839 16451 21845
rect 16758 21836 16764 21848
rect 16816 21836 16822 21888
rect 18141 21879 18199 21885
rect 18141 21845 18153 21879
rect 18187 21876 18199 21879
rect 18322 21876 18328 21888
rect 18187 21848 18328 21876
rect 18187 21845 18199 21848
rect 18141 21839 18199 21845
rect 18322 21836 18328 21848
rect 18380 21836 18386 21888
rect 18598 21876 18604 21888
rect 18559 21848 18604 21876
rect 18598 21836 18604 21848
rect 18656 21836 18662 21888
rect 24302 21836 24308 21888
rect 24360 21876 24366 21888
rect 24581 21879 24639 21885
rect 24581 21876 24593 21879
rect 24360 21848 24593 21876
rect 24360 21836 24366 21848
rect 24581 21845 24593 21848
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 25593 21879 25651 21885
rect 25593 21845 25605 21879
rect 25639 21876 25651 21879
rect 26418 21876 26424 21888
rect 25639 21848 26424 21876
rect 25639 21845 25651 21848
rect 25593 21839 25651 21845
rect 26418 21836 26424 21848
rect 26476 21836 26482 21888
rect 26528 21876 26556 21916
rect 31481 21913 31493 21947
rect 31527 21944 31539 21947
rect 31846 21944 31852 21956
rect 31527 21916 31852 21944
rect 31527 21913 31539 21916
rect 31481 21907 31539 21913
rect 31846 21904 31852 21916
rect 31904 21904 31910 21956
rect 32048 21944 32076 21975
rect 32214 21972 32220 21984
rect 32272 21972 32278 22024
rect 32309 22015 32367 22021
rect 32309 21981 32321 22015
rect 32355 22012 32367 22015
rect 32398 22012 32404 22024
rect 32355 21984 32404 22012
rect 32355 21981 32367 21984
rect 32309 21975 32367 21981
rect 32398 21972 32404 21984
rect 32456 21972 32462 22024
rect 34790 21972 34796 22024
rect 34848 22012 34854 22024
rect 34885 22015 34943 22021
rect 34885 22012 34897 22015
rect 34848 21984 34897 22012
rect 34848 21972 34854 21984
rect 34885 21981 34897 21984
rect 34931 21981 34943 22015
rect 34885 21975 34943 21981
rect 35253 22015 35311 22021
rect 35253 21981 35265 22015
rect 35299 22012 35311 22015
rect 36372 22012 36400 22043
rect 36722 22012 36728 22024
rect 35299 21984 36308 22012
rect 36372 21984 36728 22012
rect 35299 21981 35311 21984
rect 35253 21975 35311 21981
rect 32122 21944 32128 21956
rect 32048 21916 32128 21944
rect 32122 21904 32128 21916
rect 32180 21904 32186 21956
rect 34057 21879 34115 21885
rect 34057 21876 34069 21879
rect 26528 21848 34069 21876
rect 34057 21845 34069 21848
rect 34103 21876 34115 21879
rect 34900 21876 34928 21975
rect 35434 21904 35440 21956
rect 35492 21944 35498 21956
rect 35897 21947 35955 21953
rect 35897 21944 35909 21947
rect 35492 21916 35909 21944
rect 35492 21904 35498 21916
rect 35897 21913 35909 21916
rect 35943 21913 35955 21947
rect 36280 21944 36308 21984
rect 36722 21972 36728 21984
rect 36780 22012 36786 22024
rect 37553 22015 37611 22021
rect 37553 22012 37565 22015
rect 36780 21984 37565 22012
rect 36780 21972 36786 21984
rect 37553 21981 37565 21984
rect 37599 21981 37611 22015
rect 37826 22012 37832 22024
rect 37787 21984 37832 22012
rect 37553 21975 37611 21981
rect 37826 21972 37832 21984
rect 37884 22012 37890 22024
rect 38286 22012 38292 22024
rect 37884 21984 38292 22012
rect 37884 21972 37890 21984
rect 38286 21972 38292 21984
rect 38344 21972 38350 22024
rect 39850 22012 39856 22024
rect 39811 21984 39856 22012
rect 39850 21972 39856 21984
rect 39908 21972 39914 22024
rect 40420 21944 40448 22120
rect 40494 22040 40500 22092
rect 40552 22080 40558 22092
rect 40589 22083 40647 22089
rect 40589 22080 40601 22083
rect 40552 22052 40601 22080
rect 40552 22040 40558 22052
rect 40589 22049 40601 22052
rect 40635 22049 40647 22083
rect 40696 22080 40724 22120
rect 46106 22080 46112 22092
rect 40696 22052 46112 22080
rect 40589 22043 40647 22049
rect 46106 22040 46112 22052
rect 46164 22040 46170 22092
rect 36280 21916 40448 21944
rect 35897 21907 35955 21913
rect 41874 21904 41880 21956
rect 41932 21904 41938 21956
rect 37366 21876 37372 21888
rect 34103 21848 34928 21876
rect 37327 21848 37372 21876
rect 34103 21845 34115 21848
rect 34057 21839 34115 21845
rect 37366 21836 37372 21848
rect 37424 21836 37430 21888
rect 37734 21876 37740 21888
rect 37695 21848 37740 21876
rect 37734 21836 37740 21848
rect 37792 21836 37798 21888
rect 1104 21786 68816 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 68816 21786
rect 1104 21712 68816 21734
rect 5350 21632 5356 21684
rect 5408 21672 5414 21684
rect 5445 21675 5503 21681
rect 5445 21672 5457 21675
rect 5408 21644 5457 21672
rect 5408 21632 5414 21644
rect 5445 21641 5457 21644
rect 5491 21641 5503 21675
rect 5810 21672 5816 21684
rect 5771 21644 5816 21672
rect 5445 21635 5503 21641
rect 5810 21632 5816 21644
rect 5868 21632 5874 21684
rect 5902 21632 5908 21684
rect 5960 21672 5966 21684
rect 8021 21675 8079 21681
rect 8021 21672 8033 21675
rect 5960 21644 8033 21672
rect 5960 21632 5966 21644
rect 8021 21641 8033 21644
rect 8067 21641 8079 21675
rect 8021 21635 8079 21641
rect 10965 21675 11023 21681
rect 10965 21641 10977 21675
rect 11011 21641 11023 21675
rect 20254 21672 20260 21684
rect 10965 21635 11023 21641
rect 17236 21644 20260 21672
rect 8036 21604 8064 21635
rect 10980 21604 11008 21635
rect 17236 21616 17264 21644
rect 20254 21632 20260 21644
rect 20312 21632 20318 21684
rect 20806 21632 20812 21684
rect 20864 21672 20870 21684
rect 20901 21675 20959 21681
rect 20901 21672 20913 21675
rect 20864 21644 20913 21672
rect 20864 21632 20870 21644
rect 20901 21641 20913 21644
rect 20947 21641 20959 21675
rect 21266 21672 21272 21684
rect 21227 21644 21272 21672
rect 20901 21635 20959 21641
rect 21266 21632 21272 21644
rect 21324 21632 21330 21684
rect 21818 21632 21824 21684
rect 21876 21672 21882 21684
rect 23658 21672 23664 21684
rect 21876 21644 23664 21672
rect 21876 21632 21882 21644
rect 23658 21632 23664 21644
rect 23716 21632 23722 21684
rect 24581 21675 24639 21681
rect 24581 21641 24593 21675
rect 24627 21672 24639 21675
rect 26234 21672 26240 21684
rect 24627 21644 26240 21672
rect 24627 21641 24639 21644
rect 24581 21635 24639 21641
rect 26234 21632 26240 21644
rect 26292 21632 26298 21684
rect 26421 21675 26479 21681
rect 26421 21641 26433 21675
rect 26467 21672 26479 21675
rect 27154 21672 27160 21684
rect 26467 21644 27160 21672
rect 26467 21641 26479 21644
rect 26421 21635 26479 21641
rect 27154 21632 27160 21644
rect 27212 21632 27218 21684
rect 29914 21672 29920 21684
rect 29748 21644 29920 21672
rect 11762 21607 11820 21613
rect 11762 21604 11774 21607
rect 8036 21576 10916 21604
rect 10980 21576 11774 21604
rect 7098 21536 7104 21548
rect 7059 21508 7104 21536
rect 7098 21496 7104 21508
rect 7156 21496 7162 21548
rect 7926 21536 7932 21548
rect 7887 21508 7932 21536
rect 7926 21496 7932 21508
rect 7984 21496 7990 21548
rect 8202 21536 8208 21548
rect 8163 21508 8208 21536
rect 8202 21496 8208 21508
rect 8260 21496 8266 21548
rect 9140 21545 9168 21576
rect 9125 21539 9183 21545
rect 9125 21505 9137 21539
rect 9171 21505 9183 21539
rect 10042 21536 10048 21548
rect 9955 21508 10048 21536
rect 9125 21499 9183 21505
rect 10042 21496 10048 21508
rect 10100 21496 10106 21548
rect 10226 21536 10232 21548
rect 10187 21508 10232 21536
rect 10226 21496 10232 21508
rect 10284 21496 10290 21548
rect 10778 21536 10784 21548
rect 10739 21508 10784 21536
rect 10778 21496 10784 21508
rect 10836 21496 10842 21548
rect 10888 21536 10916 21576
rect 11762 21573 11774 21576
rect 11808 21573 11820 21607
rect 17218 21604 17224 21616
rect 11762 21567 11820 21573
rect 14200 21576 17224 21604
rect 11514 21536 11520 21548
rect 10888 21508 11376 21536
rect 11475 21508 11520 21536
rect 5261 21471 5319 21477
rect 5261 21437 5273 21471
rect 5307 21437 5319 21471
rect 5261 21431 5319 21437
rect 5353 21471 5411 21477
rect 5353 21437 5365 21471
rect 5399 21468 5411 21471
rect 6365 21471 6423 21477
rect 6365 21468 6377 21471
rect 5399 21440 6377 21468
rect 5399 21437 5411 21440
rect 5353 21431 5411 21437
rect 6365 21437 6377 21440
rect 6411 21468 6423 21471
rect 7006 21468 7012 21480
rect 6411 21440 7012 21468
rect 6411 21437 6423 21440
rect 6365 21431 6423 21437
rect 5276 21400 5304 21431
rect 7006 21428 7012 21440
rect 7064 21428 7070 21480
rect 7193 21471 7251 21477
rect 7193 21437 7205 21471
rect 7239 21468 7251 21471
rect 8938 21468 8944 21480
rect 7239 21440 8944 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 8938 21428 8944 21440
rect 8996 21428 9002 21480
rect 10060 21468 10088 21496
rect 11054 21468 11060 21480
rect 10060 21440 11060 21468
rect 11054 21428 11060 21440
rect 11112 21428 11118 21480
rect 11348 21468 11376 21508
rect 11514 21496 11520 21508
rect 11572 21496 11578 21548
rect 14200 21545 14228 21576
rect 17218 21564 17224 21576
rect 17276 21564 17282 21616
rect 17862 21604 17868 21616
rect 17512 21576 17868 21604
rect 13357 21539 13415 21545
rect 13357 21536 13369 21539
rect 11624 21508 13369 21536
rect 11624 21468 11652 21508
rect 13357 21505 13369 21508
rect 13403 21505 13415 21539
rect 13357 21499 13415 21505
rect 14185 21539 14243 21545
rect 14185 21505 14197 21539
rect 14231 21505 14243 21539
rect 14185 21499 14243 21505
rect 15105 21539 15163 21545
rect 15105 21505 15117 21539
rect 15151 21536 15163 21539
rect 15286 21536 15292 21548
rect 15151 21508 15292 21536
rect 15151 21505 15163 21508
rect 15105 21499 15163 21505
rect 15286 21496 15292 21508
rect 15344 21496 15350 21548
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21536 16727 21539
rect 16758 21536 16764 21548
rect 16715 21508 16764 21536
rect 16715 21505 16727 21508
rect 16669 21499 16727 21505
rect 16758 21496 16764 21508
rect 16816 21496 16822 21548
rect 17512 21545 17540 21576
rect 17862 21564 17868 21576
rect 17920 21564 17926 21616
rect 18506 21564 18512 21616
rect 18564 21564 18570 21616
rect 21082 21604 21088 21616
rect 20824 21576 21088 21604
rect 17497 21539 17555 21545
rect 17497 21505 17509 21539
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 20346 21496 20352 21548
rect 20404 21536 20410 21548
rect 20824 21536 20852 21576
rect 21082 21564 21088 21576
rect 21140 21564 21146 21616
rect 21174 21564 21180 21616
rect 21232 21564 21238 21616
rect 21358 21564 21364 21616
rect 21416 21604 21422 21616
rect 22741 21607 22799 21613
rect 22741 21604 22753 21607
rect 21416 21576 22753 21604
rect 21416 21564 21422 21576
rect 22741 21573 22753 21576
rect 22787 21604 22799 21607
rect 22787 21576 25544 21604
rect 22787 21573 22799 21576
rect 22741 21567 22799 21573
rect 20990 21536 20996 21548
rect 20404 21508 20852 21536
rect 20903 21508 20996 21536
rect 20404 21496 20410 21508
rect 11348 21440 11652 21468
rect 12526 21428 12532 21480
rect 12584 21468 12590 21480
rect 13909 21471 13967 21477
rect 13909 21468 13921 21471
rect 12584 21440 13921 21468
rect 12584 21428 12590 21440
rect 5442 21400 5448 21412
rect 5276 21372 5448 21400
rect 5442 21360 5448 21372
rect 5500 21400 5506 21412
rect 7558 21400 7564 21412
rect 5500 21372 7564 21400
rect 5500 21360 5506 21372
rect 7558 21360 7564 21372
rect 7616 21360 7622 21412
rect 9309 21403 9367 21409
rect 9309 21369 9321 21403
rect 9355 21400 9367 21403
rect 9490 21400 9496 21412
rect 9355 21372 9496 21400
rect 9355 21369 9367 21372
rect 9309 21363 9367 21369
rect 9490 21360 9496 21372
rect 9548 21360 9554 21412
rect 12912 21409 12940 21440
rect 13909 21437 13921 21440
rect 13955 21437 13967 21471
rect 17770 21468 17776 21480
rect 17731 21440 17776 21468
rect 13909 21431 13967 21437
rect 17770 21428 17776 21440
rect 17828 21428 17834 21480
rect 20732 21477 20760 21508
rect 20717 21471 20775 21477
rect 20717 21437 20729 21471
rect 20763 21437 20775 21471
rect 20717 21431 20775 21437
rect 20809 21471 20867 21477
rect 20809 21437 20821 21471
rect 20855 21468 20867 21471
rect 20916 21468 20944 21508
rect 20990 21496 20996 21508
rect 21048 21536 21054 21548
rect 21192 21536 21220 21564
rect 22922 21536 22928 21548
rect 21048 21508 21220 21536
rect 22835 21508 22928 21536
rect 21048 21496 21054 21508
rect 22922 21496 22928 21508
rect 22980 21536 22986 21548
rect 24121 21539 24179 21545
rect 24121 21536 24133 21539
rect 22980 21508 24133 21536
rect 22980 21496 22986 21508
rect 24121 21505 24133 21508
rect 24167 21505 24179 21539
rect 25516 21536 25544 21576
rect 25516 21508 25912 21536
rect 24121 21499 24179 21505
rect 20855 21440 20944 21468
rect 20855 21437 20867 21440
rect 20809 21431 20867 21437
rect 21174 21428 21180 21480
rect 21232 21468 21238 21480
rect 25498 21468 25504 21480
rect 21232 21440 25504 21468
rect 21232 21428 21238 21440
rect 25498 21428 25504 21440
rect 25556 21428 25562 21480
rect 25774 21468 25780 21480
rect 25735 21440 25780 21468
rect 25774 21428 25780 21440
rect 25832 21428 25838 21480
rect 25884 21468 25912 21508
rect 26050 21496 26056 21548
rect 26108 21536 26114 21548
rect 26145 21539 26203 21545
rect 26145 21536 26157 21539
rect 26108 21508 26157 21536
rect 26108 21496 26114 21508
rect 26145 21505 26157 21508
rect 26191 21505 26203 21539
rect 26145 21499 26203 21505
rect 26237 21539 26295 21545
rect 26237 21505 26249 21539
rect 26283 21536 26295 21539
rect 26694 21536 26700 21548
rect 26283 21508 26700 21536
rect 26283 21505 26295 21508
rect 26237 21499 26295 21505
rect 26694 21496 26700 21508
rect 26752 21536 26758 21548
rect 27154 21536 27160 21548
rect 26752 21508 27160 21536
rect 26752 21496 26758 21508
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 27798 21496 27804 21548
rect 27856 21536 27862 21548
rect 28813 21539 28871 21545
rect 28813 21536 28825 21539
rect 27856 21508 28825 21536
rect 27856 21496 27862 21508
rect 28813 21505 28825 21508
rect 28859 21505 28871 21539
rect 29638 21536 29644 21548
rect 29599 21508 29644 21536
rect 28813 21499 28871 21505
rect 29638 21496 29644 21508
rect 29696 21496 29702 21548
rect 29748 21545 29776 21644
rect 29914 21632 29920 21644
rect 29972 21632 29978 21684
rect 30101 21675 30159 21681
rect 30101 21641 30113 21675
rect 30147 21672 30159 21675
rect 30282 21672 30288 21684
rect 30147 21644 30288 21672
rect 30147 21641 30159 21644
rect 30101 21635 30159 21641
rect 30282 21632 30288 21644
rect 30340 21632 30346 21684
rect 30374 21632 30380 21684
rect 30432 21672 30438 21684
rect 30432 21644 46888 21672
rect 30432 21632 30438 21644
rect 29822 21564 29828 21616
rect 29880 21604 29886 21616
rect 34701 21607 34759 21613
rect 29880 21576 30604 21604
rect 29880 21564 29886 21576
rect 29733 21539 29791 21545
rect 29733 21505 29745 21539
rect 29779 21505 29791 21539
rect 29914 21536 29920 21548
rect 29875 21508 29920 21536
rect 29733 21499 29791 21505
rect 29748 21468 29776 21499
rect 29914 21496 29920 21508
rect 29972 21496 29978 21548
rect 30576 21545 30604 21576
rect 34701 21573 34713 21607
rect 34747 21604 34759 21607
rect 35526 21604 35532 21616
rect 34747 21576 35532 21604
rect 34747 21573 34759 21576
rect 34701 21567 34759 21573
rect 35526 21564 35532 21576
rect 35584 21564 35590 21616
rect 45830 21564 45836 21616
rect 45888 21564 45894 21616
rect 30561 21539 30619 21545
rect 30561 21505 30573 21539
rect 30607 21505 30619 21539
rect 30742 21536 30748 21548
rect 30703 21508 30748 21536
rect 30561 21499 30619 21505
rect 30742 21496 30748 21508
rect 30800 21496 30806 21548
rect 32306 21536 32312 21548
rect 32267 21508 32312 21536
rect 32306 21496 32312 21508
rect 32364 21496 32370 21548
rect 32398 21496 32404 21548
rect 32456 21536 32462 21548
rect 32456 21508 32501 21536
rect 32456 21496 32462 21508
rect 35710 21496 35716 21548
rect 35768 21536 35774 21548
rect 36541 21539 36599 21545
rect 36541 21536 36553 21539
rect 35768 21508 36553 21536
rect 35768 21496 35774 21508
rect 36541 21505 36553 21508
rect 36587 21505 36599 21539
rect 36722 21536 36728 21548
rect 36683 21508 36728 21536
rect 36541 21499 36599 21505
rect 36722 21496 36728 21508
rect 36780 21496 36786 21548
rect 37277 21539 37335 21545
rect 37277 21505 37289 21539
rect 37323 21536 37335 21539
rect 38013 21539 38071 21545
rect 38013 21536 38025 21539
rect 37323 21508 38025 21536
rect 37323 21505 37335 21508
rect 37277 21499 37335 21505
rect 38013 21505 38025 21508
rect 38059 21536 38071 21539
rect 38102 21536 38108 21548
rect 38059 21508 38108 21536
rect 38059 21505 38071 21508
rect 38013 21499 38071 21505
rect 38102 21496 38108 21508
rect 38160 21496 38166 21548
rect 44266 21536 44272 21548
rect 44227 21508 44272 21536
rect 44266 21496 44272 21508
rect 44324 21496 44330 21548
rect 45741 21539 45799 21545
rect 45741 21505 45753 21539
rect 45787 21536 45799 21539
rect 45848 21536 45876 21564
rect 46860 21548 46888 21644
rect 46014 21536 46020 21548
rect 45787 21508 45876 21536
rect 45975 21508 46020 21536
rect 45787 21505 45799 21508
rect 45741 21499 45799 21505
rect 46014 21496 46020 21508
rect 46072 21496 46078 21548
rect 46842 21536 46848 21548
rect 46803 21508 46848 21536
rect 46842 21496 46848 21508
rect 46900 21496 46906 21548
rect 30760 21468 30788 21496
rect 32674 21468 32680 21480
rect 25884 21440 28580 21468
rect 29748 21440 30788 21468
rect 32635 21440 32680 21468
rect 12897 21403 12955 21409
rect 12897 21369 12909 21403
rect 12943 21369 12955 21403
rect 28442 21400 28448 21412
rect 12897 21363 12955 21369
rect 18800 21372 28448 21400
rect 7374 21332 7380 21344
rect 7335 21304 7380 21332
rect 7374 21292 7380 21304
rect 7432 21292 7438 21344
rect 8386 21332 8392 21344
rect 8347 21304 8392 21332
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 9398 21292 9404 21344
rect 9456 21332 9462 21344
rect 10137 21335 10195 21341
rect 10137 21332 10149 21335
rect 9456 21304 10149 21332
rect 9456 21292 9462 21304
rect 10137 21301 10149 21304
rect 10183 21301 10195 21335
rect 10137 21295 10195 21301
rect 14734 21292 14740 21344
rect 14792 21332 14798 21344
rect 14921 21335 14979 21341
rect 14921 21332 14933 21335
rect 14792 21304 14933 21332
rect 14792 21292 14798 21304
rect 14921 21301 14933 21304
rect 14967 21301 14979 21335
rect 16850 21332 16856 21344
rect 16811 21304 16856 21332
rect 14921 21295 14979 21301
rect 16850 21292 16856 21304
rect 16908 21292 16914 21344
rect 16942 21292 16948 21344
rect 17000 21332 17006 21344
rect 18800 21332 18828 21372
rect 28442 21360 28448 21372
rect 28500 21360 28506 21412
rect 28552 21400 28580 21440
rect 32674 21428 32680 21440
rect 32732 21428 32738 21480
rect 32766 21428 32772 21480
rect 32824 21468 32830 21480
rect 35250 21468 35256 21480
rect 32824 21440 32869 21468
rect 35211 21440 35256 21468
rect 32824 21428 32830 21440
rect 35250 21428 35256 21440
rect 35308 21428 35314 21480
rect 35434 21468 35440 21480
rect 35395 21440 35440 21468
rect 35434 21428 35440 21440
rect 35492 21428 35498 21480
rect 37366 21428 37372 21480
rect 37424 21468 37430 21480
rect 37921 21471 37979 21477
rect 37921 21468 37933 21471
rect 37424 21440 37933 21468
rect 37424 21428 37430 21440
rect 37921 21437 37933 21440
rect 37967 21437 37979 21471
rect 37921 21431 37979 21437
rect 43806 21428 43812 21480
rect 43864 21468 43870 21480
rect 44085 21471 44143 21477
rect 44085 21468 44097 21471
rect 43864 21440 44097 21468
rect 43864 21428 43870 21440
rect 44085 21437 44097 21440
rect 44131 21437 44143 21471
rect 44085 21431 44143 21437
rect 31846 21400 31852 21412
rect 28552 21372 31852 21400
rect 31846 21360 31852 21372
rect 31904 21360 31910 21412
rect 31938 21360 31944 21412
rect 31996 21400 32002 21412
rect 32125 21403 32183 21409
rect 32125 21400 32137 21403
rect 31996 21372 32137 21400
rect 31996 21360 32002 21372
rect 32125 21369 32137 21372
rect 32171 21369 32183 21403
rect 32125 21363 32183 21369
rect 32858 21360 32864 21412
rect 32916 21400 32922 21412
rect 33321 21403 33379 21409
rect 33321 21400 33333 21403
rect 32916 21372 33333 21400
rect 32916 21360 32922 21372
rect 33321 21369 33333 21372
rect 33367 21400 33379 21403
rect 37550 21400 37556 21412
rect 33367 21372 37556 21400
rect 33367 21369 33379 21372
rect 33321 21363 33379 21369
rect 37550 21360 37556 21372
rect 37608 21360 37614 21412
rect 17000 21304 18828 21332
rect 17000 21292 17006 21304
rect 18966 21292 18972 21344
rect 19024 21332 19030 21344
rect 19245 21335 19303 21341
rect 19245 21332 19257 21335
rect 19024 21304 19257 21332
rect 19024 21292 19030 21304
rect 19245 21301 19257 21304
rect 19291 21301 19303 21335
rect 19245 21295 19303 21301
rect 19889 21335 19947 21341
rect 19889 21301 19901 21335
rect 19935 21332 19947 21335
rect 20162 21332 20168 21344
rect 19935 21304 20168 21332
rect 19935 21301 19947 21304
rect 19889 21295 19947 21301
rect 20162 21292 20168 21304
rect 20220 21292 20226 21344
rect 20898 21292 20904 21344
rect 20956 21332 20962 21344
rect 21818 21332 21824 21344
rect 20956 21304 21824 21332
rect 20956 21292 20962 21304
rect 21818 21292 21824 21304
rect 21876 21292 21882 21344
rect 24397 21335 24455 21341
rect 24397 21301 24409 21335
rect 24443 21332 24455 21335
rect 24486 21332 24492 21344
rect 24443 21304 24492 21332
rect 24443 21301 24455 21304
rect 24397 21295 24455 21301
rect 24486 21292 24492 21304
rect 24544 21292 24550 21344
rect 24762 21292 24768 21344
rect 24820 21332 24826 21344
rect 25041 21335 25099 21341
rect 25041 21332 25053 21335
rect 24820 21304 25053 21332
rect 24820 21292 24826 21304
rect 25041 21301 25053 21304
rect 25087 21301 25099 21335
rect 27798 21332 27804 21344
rect 27759 21304 27804 21332
rect 25041 21295 25099 21301
rect 27798 21292 27804 21304
rect 27856 21292 27862 21344
rect 28353 21335 28411 21341
rect 28353 21301 28365 21335
rect 28399 21332 28411 21335
rect 28534 21332 28540 21344
rect 28399 21304 28540 21332
rect 28399 21301 28411 21304
rect 28353 21295 28411 21301
rect 28534 21292 28540 21304
rect 28592 21292 28598 21344
rect 30466 21292 30472 21344
rect 30524 21332 30530 21344
rect 30653 21335 30711 21341
rect 30653 21332 30665 21335
rect 30524 21304 30665 21332
rect 30524 21292 30530 21304
rect 30653 21301 30665 21304
rect 30699 21301 30711 21335
rect 30653 21295 30711 21301
rect 34606 21292 34612 21344
rect 34664 21332 34670 21344
rect 34882 21332 34888 21344
rect 34664 21304 34888 21332
rect 34664 21292 34670 21304
rect 34882 21292 34888 21304
rect 34940 21292 34946 21344
rect 35897 21335 35955 21341
rect 35897 21301 35909 21335
rect 35943 21332 35955 21335
rect 36262 21332 36268 21344
rect 35943 21304 36268 21332
rect 35943 21301 35955 21304
rect 35897 21295 35955 21301
rect 36262 21292 36268 21304
rect 36320 21292 36326 21344
rect 36725 21335 36783 21341
rect 36725 21301 36737 21335
rect 36771 21332 36783 21335
rect 37734 21332 37740 21344
rect 36771 21304 37740 21332
rect 36771 21301 36783 21304
rect 36725 21295 36783 21301
rect 37734 21292 37740 21304
rect 37792 21292 37798 21344
rect 38289 21335 38347 21341
rect 38289 21301 38301 21335
rect 38335 21332 38347 21335
rect 39850 21332 39856 21344
rect 38335 21304 39856 21332
rect 38335 21301 38347 21304
rect 38289 21295 38347 21301
rect 39850 21292 39856 21304
rect 39908 21292 39914 21344
rect 42334 21292 42340 21344
rect 42392 21332 42398 21344
rect 43898 21332 43904 21344
rect 42392 21304 43904 21332
rect 42392 21292 42398 21304
rect 43898 21292 43904 21304
rect 43956 21292 43962 21344
rect 44453 21335 44511 21341
rect 44453 21301 44465 21335
rect 44499 21332 44511 21335
rect 45002 21332 45008 21344
rect 44499 21304 45008 21332
rect 44499 21301 44511 21304
rect 44453 21295 44511 21301
rect 45002 21292 45008 21304
rect 45060 21292 45066 21344
rect 1104 21242 68816 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 65654 21242
rect 65706 21190 65718 21242
rect 65770 21190 65782 21242
rect 65834 21190 65846 21242
rect 65898 21190 65910 21242
rect 65962 21190 68816 21242
rect 1104 21168 68816 21190
rect 8938 21088 8944 21140
rect 8996 21128 9002 21140
rect 10505 21131 10563 21137
rect 10505 21128 10517 21131
rect 8996 21100 10517 21128
rect 8996 21088 9002 21100
rect 10505 21097 10517 21100
rect 10551 21097 10563 21131
rect 10505 21091 10563 21097
rect 10778 21088 10784 21140
rect 10836 21128 10842 21140
rect 11425 21131 11483 21137
rect 11425 21128 11437 21131
rect 10836 21100 11437 21128
rect 10836 21088 10842 21100
rect 11425 21097 11437 21100
rect 11471 21097 11483 21131
rect 11425 21091 11483 21097
rect 11698 21088 11704 21140
rect 11756 21128 11762 21140
rect 11756 21100 12112 21128
rect 11756 21088 11762 21100
rect 7006 21020 7012 21072
rect 7064 21060 7070 21072
rect 7064 21032 11928 21060
rect 7064 21020 7070 21032
rect 6549 20995 6607 21001
rect 6549 20961 6561 20995
rect 6595 20992 6607 20995
rect 6638 20992 6644 21004
rect 6595 20964 6644 20992
rect 6595 20961 6607 20964
rect 6549 20955 6607 20961
rect 6638 20952 6644 20964
rect 6696 20952 6702 21004
rect 6914 20952 6920 21004
rect 6972 20992 6978 21004
rect 7469 20995 7527 21001
rect 7469 20992 7481 20995
rect 6972 20964 7481 20992
rect 6972 20952 6978 20964
rect 7469 20961 7481 20964
rect 7515 20961 7527 20995
rect 7469 20955 7527 20961
rect 6270 20856 6276 20868
rect 6328 20865 6334 20868
rect 6240 20828 6276 20856
rect 6270 20816 6276 20828
rect 6328 20819 6340 20865
rect 7098 20856 7104 20868
rect 6564 20828 7104 20856
rect 6328 20816 6334 20819
rect 5169 20791 5227 20797
rect 5169 20757 5181 20791
rect 5215 20788 5227 20791
rect 6564 20788 6592 20828
rect 7098 20816 7104 20828
rect 7156 20856 7162 20868
rect 7377 20859 7435 20865
rect 7377 20856 7389 20859
rect 7156 20828 7389 20856
rect 7156 20816 7162 20828
rect 7377 20825 7389 20828
rect 7423 20825 7435 20859
rect 7484 20856 7512 20955
rect 7558 20952 7564 21004
rect 7616 20992 7622 21004
rect 7616 20964 7661 20992
rect 7616 20952 7622 20964
rect 8294 20952 8300 21004
rect 8352 20992 8358 21004
rect 10873 20995 10931 21001
rect 8352 20964 9628 20992
rect 8352 20952 8358 20964
rect 8202 20884 8208 20936
rect 8260 20924 8266 20936
rect 9263 20927 9321 20933
rect 9263 20924 9275 20927
rect 8260 20896 9275 20924
rect 8260 20884 8266 20896
rect 9263 20893 9275 20896
rect 9309 20893 9321 20927
rect 9263 20887 9321 20893
rect 9398 20884 9404 20936
rect 9456 20924 9462 20936
rect 9600 20933 9628 20964
rect 10873 20961 10885 20995
rect 10919 20992 10931 20995
rect 11054 20992 11060 21004
rect 10919 20964 11060 20992
rect 10919 20961 10931 20964
rect 10873 20955 10931 20961
rect 11054 20952 11060 20964
rect 11112 20952 11118 21004
rect 11900 21001 11928 21032
rect 12084 21001 12112 21100
rect 14274 21088 14280 21140
rect 14332 21128 14338 21140
rect 16577 21131 16635 21137
rect 14332 21100 16528 21128
rect 14332 21088 14338 21100
rect 11885 20995 11943 21001
rect 11885 20992 11897 20995
rect 11716 20964 11897 20992
rect 9600 20927 9679 20933
rect 9456 20896 9501 20924
rect 9600 20896 9633 20927
rect 9456 20884 9462 20896
rect 9621 20893 9633 20896
rect 9667 20893 9679 20927
rect 9621 20887 9679 20893
rect 9766 20884 9772 20936
rect 9824 20924 9830 20936
rect 10781 20927 10839 20933
rect 9824 20896 9869 20924
rect 9824 20884 9830 20896
rect 10781 20893 10793 20927
rect 10827 20924 10839 20927
rect 11238 20924 11244 20936
rect 10827 20896 11244 20924
rect 10827 20893 10839 20896
rect 10781 20887 10839 20893
rect 11238 20884 11244 20896
rect 11296 20884 11302 20936
rect 9490 20856 9496 20868
rect 7484 20828 9352 20856
rect 9451 20828 9496 20856
rect 7377 20819 7435 20825
rect 7006 20788 7012 20800
rect 5215 20760 6592 20788
rect 6967 20760 7012 20788
rect 5215 20757 5227 20760
rect 5169 20751 5227 20757
rect 7006 20748 7012 20760
rect 7064 20748 7070 20800
rect 9125 20791 9183 20797
rect 9125 20757 9137 20791
rect 9171 20788 9183 20791
rect 9214 20788 9220 20800
rect 9171 20760 9220 20788
rect 9171 20757 9183 20760
rect 9125 20751 9183 20757
rect 9214 20748 9220 20760
rect 9272 20748 9278 20800
rect 9324 20788 9352 20828
rect 9490 20816 9496 20828
rect 9548 20816 9554 20868
rect 11606 20788 11612 20800
rect 9324 20760 11612 20788
rect 11606 20748 11612 20760
rect 11664 20748 11670 20800
rect 11716 20788 11744 20964
rect 11885 20961 11897 20964
rect 11931 20961 11943 20995
rect 11885 20955 11943 20961
rect 12069 20995 12127 21001
rect 12069 20961 12081 20995
rect 12115 20992 12127 20995
rect 12250 20992 12256 21004
rect 12115 20964 12256 20992
rect 12115 20961 12127 20964
rect 12069 20955 12127 20961
rect 12250 20952 12256 20964
rect 12308 20952 12314 21004
rect 13906 20952 13912 21004
rect 13964 20992 13970 21004
rect 14458 20992 14464 21004
rect 13964 20964 14464 20992
rect 13964 20952 13970 20964
rect 14458 20952 14464 20964
rect 14516 20952 14522 21004
rect 11793 20927 11851 20933
rect 11793 20893 11805 20927
rect 11839 20924 11851 20927
rect 12526 20924 12532 20936
rect 11839 20896 12532 20924
rect 11839 20893 11851 20896
rect 11793 20887 11851 20893
rect 12526 20884 12532 20896
rect 12584 20884 12590 20936
rect 14734 20933 14740 20936
rect 14728 20924 14740 20933
rect 14695 20896 14740 20924
rect 14728 20887 14740 20896
rect 14734 20884 14740 20887
rect 14792 20884 14798 20936
rect 15010 20884 15016 20936
rect 15068 20924 15074 20936
rect 15068 20896 16436 20924
rect 15068 20884 15074 20896
rect 13538 20816 13544 20868
rect 13596 20856 13602 20868
rect 16022 20856 16028 20868
rect 13596 20828 16028 20856
rect 13596 20816 13602 20828
rect 16022 20816 16028 20828
rect 16080 20816 16086 20868
rect 12713 20791 12771 20797
rect 12713 20788 12725 20791
rect 11716 20760 12725 20788
rect 12713 20757 12725 20760
rect 12759 20788 12771 20791
rect 14182 20788 14188 20800
rect 12759 20760 14188 20788
rect 12759 20757 12771 20760
rect 12713 20751 12771 20757
rect 14182 20748 14188 20760
rect 14240 20748 14246 20800
rect 15838 20788 15844 20800
rect 15799 20760 15844 20788
rect 15838 20748 15844 20760
rect 15896 20748 15902 20800
rect 16408 20788 16436 20896
rect 16500 20856 16528 21100
rect 16577 21097 16589 21131
rect 16623 21128 16635 21131
rect 16942 21128 16948 21140
rect 16623 21100 16948 21128
rect 16623 21097 16635 21100
rect 16577 21091 16635 21097
rect 16942 21088 16948 21100
rect 17000 21088 17006 21140
rect 17954 21088 17960 21140
rect 18012 21128 18018 21140
rect 18417 21131 18475 21137
rect 18417 21128 18429 21131
rect 18012 21100 18429 21128
rect 18012 21088 18018 21100
rect 18417 21097 18429 21100
rect 18463 21097 18475 21131
rect 18417 21091 18475 21097
rect 20162 21088 20168 21140
rect 20220 21128 20226 21140
rect 21174 21128 21180 21140
rect 20220 21100 21180 21128
rect 20220 21088 20226 21100
rect 21174 21088 21180 21100
rect 21232 21088 21238 21140
rect 23566 21128 23572 21140
rect 23479 21100 23572 21128
rect 23566 21088 23572 21100
rect 23624 21128 23630 21140
rect 24486 21128 24492 21140
rect 23624 21100 24492 21128
rect 23624 21088 23630 21100
rect 24486 21088 24492 21100
rect 24544 21088 24550 21140
rect 25590 21088 25596 21140
rect 25648 21128 25654 21140
rect 25685 21131 25743 21137
rect 25685 21128 25697 21131
rect 25648 21100 25697 21128
rect 25648 21088 25654 21100
rect 25685 21097 25697 21100
rect 25731 21097 25743 21131
rect 28442 21128 28448 21140
rect 28403 21100 28448 21128
rect 25685 21091 25743 21097
rect 28442 21088 28448 21100
rect 28500 21088 28506 21140
rect 29914 21128 29920 21140
rect 28736 21100 29920 21128
rect 25038 21060 25044 21072
rect 24999 21032 25044 21060
rect 25038 21020 25044 21032
rect 25096 21020 25102 21072
rect 27893 21063 27951 21069
rect 27893 21029 27905 21063
rect 27939 21060 27951 21063
rect 28736 21060 28764 21100
rect 29914 21088 29920 21100
rect 29972 21088 29978 21140
rect 30742 21088 30748 21140
rect 30800 21128 30806 21140
rect 30837 21131 30895 21137
rect 30837 21128 30849 21131
rect 30800 21100 30849 21128
rect 30800 21088 30806 21100
rect 30837 21097 30849 21100
rect 30883 21097 30895 21131
rect 30837 21091 30895 21097
rect 32125 21131 32183 21137
rect 32125 21097 32137 21131
rect 32171 21128 32183 21131
rect 32674 21128 32680 21140
rect 32171 21100 32680 21128
rect 32171 21097 32183 21100
rect 32125 21091 32183 21097
rect 32674 21088 32680 21100
rect 32732 21088 32738 21140
rect 35710 21128 35716 21140
rect 35671 21100 35716 21128
rect 35710 21088 35716 21100
rect 35768 21088 35774 21140
rect 39945 21131 40003 21137
rect 39945 21097 39957 21131
rect 39991 21128 40003 21131
rect 40126 21128 40132 21140
rect 39991 21100 40132 21128
rect 39991 21097 40003 21100
rect 39945 21091 40003 21097
rect 40126 21088 40132 21100
rect 40184 21088 40190 21140
rect 41785 21131 41843 21137
rect 41785 21097 41797 21131
rect 41831 21128 41843 21131
rect 41874 21128 41880 21140
rect 41831 21100 41880 21128
rect 41831 21097 41843 21100
rect 41785 21091 41843 21097
rect 41874 21088 41880 21100
rect 41932 21088 41938 21140
rect 46106 21128 46112 21140
rect 42720 21100 46112 21128
rect 27939 21032 28764 21060
rect 28813 21063 28871 21069
rect 27939 21029 27951 21032
rect 27893 21023 27951 21029
rect 28813 21029 28825 21063
rect 28859 21060 28871 21063
rect 29825 21063 29883 21069
rect 29825 21060 29837 21063
rect 28859 21032 29837 21060
rect 28859 21029 28871 21032
rect 28813 21023 28871 21029
rect 29825 21029 29837 21032
rect 29871 21029 29883 21063
rect 29825 21023 29883 21029
rect 18874 20952 18880 21004
rect 18932 20992 18938 21004
rect 19245 20995 19303 21001
rect 19245 20992 19257 20995
rect 18932 20964 19257 20992
rect 18932 20952 18938 20964
rect 19245 20961 19257 20964
rect 19291 20961 19303 20995
rect 19245 20955 19303 20961
rect 19426 20952 19432 21004
rect 19484 20992 19490 21004
rect 19521 20995 19579 21001
rect 19521 20992 19533 20995
rect 19484 20964 19533 20992
rect 19484 20952 19490 20964
rect 19521 20961 19533 20964
rect 19567 20961 19579 20995
rect 19521 20955 19579 20961
rect 20533 20995 20591 21001
rect 20533 20961 20545 20995
rect 20579 20992 20591 20995
rect 20898 20992 20904 21004
rect 20579 20964 20904 20992
rect 20579 20961 20591 20964
rect 20533 20955 20591 20961
rect 20898 20952 20904 20964
rect 20956 20952 20962 21004
rect 28828 20992 28856 21023
rect 31846 21020 31852 21072
rect 31904 21060 31910 21072
rect 31904 21032 34836 21060
rect 31904 21020 31910 21032
rect 27632 20964 28856 20992
rect 16850 20884 16856 20936
rect 16908 20924 16914 20936
rect 17690 20927 17748 20933
rect 17690 20924 17702 20927
rect 16908 20896 17702 20924
rect 16908 20884 16914 20896
rect 17690 20893 17702 20896
rect 17736 20893 17748 20927
rect 17690 20887 17748 20893
rect 17862 20884 17868 20936
rect 17920 20924 17926 20936
rect 17957 20927 18015 20933
rect 17957 20924 17969 20927
rect 17920 20896 17969 20924
rect 17920 20884 17926 20896
rect 17957 20893 17969 20896
rect 18003 20893 18015 20927
rect 17957 20887 18015 20893
rect 18601 20927 18659 20933
rect 18601 20893 18613 20927
rect 18647 20893 18659 20927
rect 20806 20924 20812 20936
rect 20767 20896 20812 20924
rect 18601 20887 18659 20893
rect 18046 20856 18052 20868
rect 16500 20828 18052 20856
rect 18046 20816 18052 20828
rect 18104 20856 18110 20868
rect 18616 20856 18644 20887
rect 20806 20884 20812 20896
rect 20864 20884 20870 20936
rect 22189 20927 22247 20933
rect 22189 20893 22201 20927
rect 22235 20924 22247 20927
rect 22278 20924 22284 20936
rect 22235 20896 22284 20924
rect 22235 20893 22247 20896
rect 22189 20887 22247 20893
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 25774 20884 25780 20936
rect 25832 20924 25838 20936
rect 25869 20927 25927 20933
rect 25869 20924 25881 20927
rect 25832 20896 25881 20924
rect 25832 20884 25838 20896
rect 25869 20893 25881 20896
rect 25915 20893 25927 20927
rect 25869 20887 25927 20893
rect 25958 20884 25964 20936
rect 26016 20924 26022 20936
rect 27632 20933 27660 20964
rect 29546 20952 29552 21004
rect 29604 20992 29610 21004
rect 30009 20995 30067 21001
rect 30009 20992 30021 20995
rect 29604 20964 30021 20992
rect 29604 20952 29610 20964
rect 30009 20961 30021 20964
rect 30055 20992 30067 20995
rect 32490 20992 32496 21004
rect 30055 20964 30696 20992
rect 30055 20961 30067 20964
rect 30009 20955 30067 20961
rect 27617 20927 27675 20933
rect 26016 20896 26061 20924
rect 26016 20884 26022 20896
rect 27617 20893 27629 20927
rect 27663 20893 27675 20927
rect 27617 20887 27675 20893
rect 28353 20927 28411 20933
rect 28353 20893 28365 20927
rect 28399 20924 28411 20927
rect 28442 20924 28448 20936
rect 28399 20896 28448 20924
rect 28399 20893 28411 20896
rect 28353 20887 28411 20893
rect 28442 20884 28448 20896
rect 28500 20924 28506 20936
rect 28500 20896 29684 20924
rect 28500 20884 28506 20896
rect 21358 20856 21364 20868
rect 18104 20828 21364 20856
rect 18104 20816 18110 20828
rect 21358 20816 21364 20828
rect 21416 20816 21422 20868
rect 22462 20865 22468 20868
rect 22456 20819 22468 20865
rect 22520 20856 22526 20868
rect 24762 20856 24768 20868
rect 22520 20828 22556 20856
rect 24723 20828 24768 20856
rect 22462 20816 22468 20819
rect 22520 20816 22526 20828
rect 24762 20816 24768 20828
rect 24820 20816 24826 20868
rect 25685 20859 25743 20865
rect 25685 20856 25697 20859
rect 25240 20828 25697 20856
rect 18782 20788 18788 20800
rect 16408 20760 18788 20788
rect 18782 20748 18788 20760
rect 18840 20748 18846 20800
rect 18966 20748 18972 20800
rect 19024 20788 19030 20800
rect 22922 20788 22928 20800
rect 19024 20760 22928 20788
rect 19024 20748 19030 20760
rect 22922 20748 22928 20760
rect 22980 20748 22986 20800
rect 25240 20797 25268 20828
rect 25685 20825 25697 20828
rect 25731 20825 25743 20859
rect 25685 20819 25743 20825
rect 27893 20859 27951 20865
rect 27893 20825 27905 20859
rect 27939 20856 27951 20859
rect 28534 20856 28540 20868
rect 27939 20828 28540 20856
rect 27939 20825 27951 20828
rect 27893 20819 27951 20825
rect 28534 20816 28540 20828
rect 28592 20856 28598 20868
rect 29549 20859 29607 20865
rect 29549 20856 29561 20859
rect 28592 20828 29561 20856
rect 28592 20816 28598 20828
rect 29549 20825 29561 20828
rect 29595 20825 29607 20859
rect 29549 20819 29607 20825
rect 25225 20791 25283 20797
rect 25225 20757 25237 20791
rect 25271 20757 25283 20791
rect 26418 20788 26424 20800
rect 26379 20760 26424 20788
rect 25225 20751 25283 20757
rect 26418 20748 26424 20760
rect 26476 20748 26482 20800
rect 27709 20791 27767 20797
rect 27709 20757 27721 20791
rect 27755 20788 27767 20791
rect 29362 20788 29368 20800
rect 27755 20760 29368 20788
rect 27755 20757 27767 20760
rect 27709 20751 27767 20757
rect 29362 20748 29368 20760
rect 29420 20748 29426 20800
rect 29656 20788 29684 20896
rect 30098 20884 30104 20936
rect 30156 20924 30162 20936
rect 30668 20933 30696 20964
rect 32048 20964 32496 20992
rect 32048 20933 32076 20964
rect 32490 20952 32496 20964
rect 32548 20952 32554 21004
rect 33502 20992 33508 21004
rect 33463 20964 33508 20992
rect 33502 20952 33508 20964
rect 33560 20952 33566 21004
rect 34808 21001 34836 21032
rect 35434 21020 35440 21072
rect 35492 21060 35498 21072
rect 35621 21063 35679 21069
rect 35621 21060 35633 21063
rect 35492 21032 35633 21060
rect 35492 21020 35498 21032
rect 35621 21029 35633 21032
rect 35667 21060 35679 21063
rect 36173 21063 36231 21069
rect 36173 21060 36185 21063
rect 35667 21032 36185 21060
rect 35667 21029 35679 21032
rect 35621 21023 35679 21029
rect 36173 21029 36185 21032
rect 36219 21029 36231 21063
rect 36173 21023 36231 21029
rect 40313 21063 40371 21069
rect 40313 21029 40325 21063
rect 40359 21060 40371 21063
rect 42426 21060 42432 21072
rect 40359 21032 42432 21060
rect 40359 21029 40371 21032
rect 40313 21023 40371 21029
rect 42426 21020 42432 21032
rect 42484 21020 42490 21072
rect 34793 20995 34851 21001
rect 34793 20961 34805 20995
rect 34839 20992 34851 20995
rect 35253 20995 35311 21001
rect 35253 20992 35265 20995
rect 34839 20964 35265 20992
rect 34839 20961 34851 20964
rect 34793 20955 34851 20961
rect 35253 20961 35265 20964
rect 35299 20961 35311 20995
rect 35253 20955 35311 20961
rect 37826 20952 37832 21004
rect 37884 20992 37890 21004
rect 38289 20995 38347 21001
rect 38289 20992 38301 20995
rect 37884 20964 38301 20992
rect 37884 20952 37890 20964
rect 38289 20961 38301 20964
rect 38335 20961 38347 20995
rect 39942 20992 39948 21004
rect 39903 20964 39948 20992
rect 38289 20955 38347 20961
rect 39942 20952 39948 20964
rect 40000 20952 40006 21004
rect 42610 20952 42616 21004
rect 42668 20992 42674 21004
rect 42720 20992 42748 21100
rect 46106 21088 46112 21100
rect 46164 21088 46170 21140
rect 42668 20964 42748 20992
rect 42668 20952 42674 20964
rect 30469 20927 30527 20933
rect 30469 20924 30481 20927
rect 30156 20896 30481 20924
rect 30156 20884 30162 20896
rect 30469 20893 30481 20896
rect 30515 20893 30527 20927
rect 30469 20887 30527 20893
rect 30653 20927 30711 20933
rect 30653 20893 30665 20927
rect 30699 20893 30711 20927
rect 30653 20887 30711 20893
rect 32033 20927 32091 20933
rect 32033 20893 32045 20927
rect 32079 20893 32091 20927
rect 32214 20924 32220 20936
rect 32175 20896 32220 20924
rect 32033 20887 32091 20893
rect 32214 20884 32220 20896
rect 32272 20884 32278 20936
rect 32677 20927 32735 20933
rect 32677 20893 32689 20927
rect 32723 20924 32735 20927
rect 32858 20924 32864 20936
rect 32723 20896 32864 20924
rect 32723 20893 32735 20896
rect 32677 20887 32735 20893
rect 30282 20816 30288 20868
rect 30340 20856 30346 20868
rect 32692 20856 32720 20887
rect 32858 20884 32864 20896
rect 32916 20884 32922 20936
rect 37553 20927 37611 20933
rect 37553 20893 37565 20927
rect 37599 20893 37611 20927
rect 37553 20887 37611 20893
rect 37274 20856 37280 20868
rect 37332 20865 37338 20868
rect 30340 20828 32720 20856
rect 37244 20828 37280 20856
rect 30340 20816 30346 20828
rect 37274 20816 37280 20828
rect 37332 20819 37344 20865
rect 37568 20856 37596 20887
rect 37734 20884 37740 20936
rect 37792 20924 37798 20936
rect 38381 20927 38439 20933
rect 38381 20924 38393 20927
rect 37792 20896 38393 20924
rect 37792 20884 37798 20896
rect 38381 20893 38393 20896
rect 38427 20924 38439 20927
rect 39850 20924 39856 20936
rect 38427 20896 39436 20924
rect 39811 20896 39856 20924
rect 38427 20893 38439 20896
rect 38381 20887 38439 20893
rect 39298 20856 39304 20868
rect 37568 20828 39304 20856
rect 37332 20816 37338 20819
rect 39298 20816 39304 20828
rect 39356 20816 39362 20868
rect 39408 20856 39436 20896
rect 39850 20884 39856 20896
rect 39908 20884 39914 20936
rect 40126 20924 40132 20936
rect 40087 20896 40132 20924
rect 40126 20884 40132 20896
rect 40184 20884 40190 20936
rect 41877 20927 41935 20933
rect 41877 20893 41889 20927
rect 41923 20924 41935 20927
rect 42334 20924 42340 20936
rect 41923 20896 42340 20924
rect 41923 20893 41935 20896
rect 41877 20887 41935 20893
rect 42334 20884 42340 20896
rect 42392 20884 42398 20936
rect 42720 20933 42748 20964
rect 42521 20927 42579 20933
rect 42521 20893 42533 20927
rect 42567 20893 42579 20927
rect 42521 20887 42579 20893
rect 42705 20927 42763 20933
rect 42705 20893 42717 20927
rect 42751 20893 42763 20927
rect 42705 20887 42763 20893
rect 41230 20856 41236 20868
rect 39408 20828 41236 20856
rect 41230 20816 41236 20828
rect 41288 20816 41294 20868
rect 35618 20788 35624 20800
rect 29656 20760 35624 20788
rect 35618 20748 35624 20760
rect 35676 20748 35682 20800
rect 38010 20788 38016 20800
rect 37971 20760 38016 20788
rect 38010 20748 38016 20760
rect 38068 20748 38074 20800
rect 40957 20791 41015 20797
rect 40957 20757 40969 20791
rect 41003 20788 41015 20791
rect 41598 20788 41604 20800
rect 41003 20760 41604 20788
rect 41003 20757 41015 20760
rect 40957 20751 41015 20757
rect 41598 20748 41604 20760
rect 41656 20748 41662 20800
rect 42536 20788 42564 20887
rect 42794 20884 42800 20936
rect 42852 20924 42858 20936
rect 43165 20927 43223 20933
rect 43165 20924 43177 20927
rect 42852 20896 43177 20924
rect 42852 20884 42858 20896
rect 43165 20893 43177 20896
rect 43211 20893 43223 20927
rect 43165 20887 43223 20893
rect 43441 20927 43499 20933
rect 43441 20893 43453 20927
rect 43487 20893 43499 20927
rect 45002 20924 45008 20936
rect 44963 20896 45008 20924
rect 43441 20887 43499 20893
rect 42613 20859 42671 20865
rect 42613 20825 42625 20859
rect 42659 20856 42671 20859
rect 43456 20856 43484 20887
rect 45002 20884 45008 20896
rect 45060 20884 45066 20936
rect 45646 20924 45652 20936
rect 45607 20896 45652 20924
rect 45646 20884 45652 20896
rect 45704 20884 45710 20936
rect 42659 20828 43484 20856
rect 44008 20828 45232 20856
rect 42659 20825 42671 20828
rect 42613 20819 42671 20825
rect 42702 20788 42708 20800
rect 42536 20760 42708 20788
rect 42702 20748 42708 20760
rect 42760 20748 42766 20800
rect 42794 20748 42800 20800
rect 42852 20788 42858 20800
rect 44008 20788 44036 20828
rect 45204 20800 45232 20828
rect 44174 20788 44180 20800
rect 42852 20760 44036 20788
rect 44135 20760 44180 20788
rect 42852 20748 42858 20760
rect 44174 20748 44180 20760
rect 44232 20748 44238 20800
rect 45186 20788 45192 20800
rect 45099 20760 45192 20788
rect 45186 20748 45192 20760
rect 45244 20748 45250 20800
rect 45833 20791 45891 20797
rect 45833 20757 45845 20791
rect 45879 20788 45891 20791
rect 46106 20788 46112 20800
rect 45879 20760 46112 20788
rect 45879 20757 45891 20760
rect 45833 20751 45891 20757
rect 46106 20748 46112 20760
rect 46164 20748 46170 20800
rect 1104 20698 68816 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 68816 20698
rect 1104 20624 68816 20646
rect 6270 20544 6276 20596
rect 6328 20584 6334 20596
rect 6365 20587 6423 20593
rect 6365 20584 6377 20587
rect 6328 20556 6377 20584
rect 6328 20544 6334 20556
rect 6365 20553 6377 20556
rect 6411 20553 6423 20587
rect 6365 20547 6423 20553
rect 9122 20544 9128 20596
rect 9180 20584 9186 20596
rect 9401 20587 9459 20593
rect 9401 20584 9413 20587
rect 9180 20556 9413 20584
rect 9180 20544 9186 20556
rect 9401 20553 9413 20556
rect 9447 20553 9459 20587
rect 9401 20547 9459 20553
rect 11238 20544 11244 20596
rect 11296 20584 11302 20596
rect 11517 20587 11575 20593
rect 11517 20584 11529 20587
rect 11296 20556 11529 20584
rect 11296 20544 11302 20556
rect 11517 20553 11529 20556
rect 11563 20553 11575 20587
rect 11517 20547 11575 20553
rect 11532 20516 11560 20547
rect 11606 20544 11612 20596
rect 11664 20584 11670 20596
rect 12342 20584 12348 20596
rect 11664 20556 12348 20584
rect 11664 20544 11670 20556
rect 12342 20544 12348 20556
rect 12400 20584 12406 20596
rect 13998 20584 14004 20596
rect 12400 20556 14004 20584
rect 12400 20544 12406 20556
rect 13998 20544 14004 20556
rect 14056 20544 14062 20596
rect 16942 20584 16948 20596
rect 14108 20556 15332 20584
rect 14108 20516 14136 20556
rect 11532 20488 14136 20516
rect 14182 20476 14188 20528
rect 14240 20516 14246 20528
rect 14369 20519 14427 20525
rect 14369 20516 14381 20519
rect 14240 20488 14381 20516
rect 14240 20476 14246 20488
rect 14369 20485 14381 20488
rect 14415 20516 14427 20519
rect 15194 20516 15200 20528
rect 14415 20488 15200 20516
rect 14415 20485 14427 20488
rect 14369 20479 14427 20485
rect 15194 20476 15200 20488
rect 15252 20476 15258 20528
rect 15304 20516 15332 20556
rect 15580 20556 16948 20584
rect 15580 20516 15608 20556
rect 16942 20544 16948 20556
rect 17000 20544 17006 20596
rect 17126 20584 17132 20596
rect 17087 20556 17132 20584
rect 17126 20544 17132 20556
rect 17184 20544 17190 20596
rect 18782 20544 18788 20596
rect 18840 20584 18846 20596
rect 18840 20556 20484 20584
rect 18840 20544 18846 20556
rect 15304 20488 15608 20516
rect 15657 20519 15715 20525
rect 15657 20485 15669 20519
rect 15703 20516 15715 20519
rect 15838 20516 15844 20528
rect 15703 20488 15844 20516
rect 15703 20485 15715 20488
rect 15657 20479 15715 20485
rect 15838 20476 15844 20488
rect 15896 20516 15902 20528
rect 18049 20519 18107 20525
rect 15896 20488 18000 20516
rect 15896 20476 15902 20488
rect 6549 20451 6607 20457
rect 6549 20417 6561 20451
rect 6595 20448 6607 20451
rect 7006 20448 7012 20460
rect 6595 20420 7012 20448
rect 6595 20417 6607 20420
rect 6549 20411 6607 20417
rect 7006 20408 7012 20420
rect 7064 20408 7070 20460
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20448 7527 20451
rect 8386 20448 8392 20460
rect 7515 20420 8392 20448
rect 7515 20417 7527 20420
rect 7469 20411 7527 20417
rect 8386 20408 8392 20420
rect 8444 20408 8450 20460
rect 8941 20451 8999 20457
rect 8941 20417 8953 20451
rect 8987 20417 8999 20451
rect 8941 20411 8999 20417
rect 7374 20380 7380 20392
rect 7335 20352 7380 20380
rect 7374 20340 7380 20352
rect 7432 20340 7438 20392
rect 8202 20340 8208 20392
rect 8260 20380 8266 20392
rect 8956 20380 8984 20411
rect 9030 20408 9036 20460
rect 9088 20448 9094 20460
rect 9214 20448 9220 20460
rect 9088 20420 9133 20448
rect 9175 20420 9220 20448
rect 9088 20408 9094 20420
rect 9214 20408 9220 20420
rect 9272 20408 9278 20460
rect 10318 20448 10324 20460
rect 10279 20420 10324 20448
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 10965 20451 11023 20457
rect 10965 20417 10977 20451
rect 11011 20448 11023 20451
rect 11974 20448 11980 20460
rect 11011 20420 11980 20448
rect 11011 20417 11023 20420
rect 10965 20411 11023 20417
rect 11974 20408 11980 20420
rect 12032 20408 12038 20460
rect 14461 20451 14519 20457
rect 14461 20417 14473 20451
rect 14507 20448 14519 20451
rect 15470 20448 15476 20460
rect 14507 20420 15476 20448
rect 14507 20417 14519 20420
rect 14461 20411 14519 20417
rect 15470 20408 15476 20420
rect 15528 20408 15534 20460
rect 17972 20457 18000 20488
rect 18049 20485 18061 20519
rect 18095 20516 18107 20519
rect 18693 20519 18751 20525
rect 18693 20516 18705 20519
rect 18095 20488 18705 20516
rect 18095 20485 18107 20488
rect 18049 20479 18107 20485
rect 18693 20485 18705 20488
rect 18739 20516 18751 20519
rect 18739 20488 19104 20516
rect 18739 20485 18751 20488
rect 18693 20479 18751 20485
rect 17037 20451 17095 20457
rect 15672 20420 15884 20448
rect 8260 20352 8984 20380
rect 8260 20340 8266 20352
rect 9306 20340 9312 20392
rect 9364 20380 9370 20392
rect 9861 20383 9919 20389
rect 9861 20380 9873 20383
rect 9364 20352 9873 20380
rect 9364 20340 9370 20352
rect 9861 20349 9873 20352
rect 9907 20349 9919 20383
rect 10336 20380 10364 20408
rect 12069 20383 12127 20389
rect 12069 20380 12081 20383
rect 10336 20352 12081 20380
rect 9861 20343 9919 20349
rect 12069 20349 12081 20352
rect 12115 20380 12127 20383
rect 12158 20380 12164 20392
rect 12115 20352 12164 20380
rect 12115 20349 12127 20352
rect 12069 20343 12127 20349
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20380 14335 20383
rect 15672 20380 15700 20420
rect 15856 20392 15884 20420
rect 17037 20417 17049 20451
rect 17083 20448 17095 20451
rect 17957 20451 18015 20457
rect 17083 20420 17816 20448
rect 17083 20417 17095 20420
rect 17037 20411 17095 20417
rect 14323 20352 15700 20380
rect 15749 20383 15807 20389
rect 14323 20349 14335 20352
rect 14277 20343 14335 20349
rect 15749 20349 15761 20383
rect 15795 20349 15807 20383
rect 15749 20343 15807 20349
rect 7837 20315 7895 20321
rect 7837 20281 7849 20315
rect 7883 20312 7895 20315
rect 9214 20312 9220 20324
rect 7883 20284 9220 20312
rect 7883 20281 7895 20284
rect 7837 20275 7895 20281
rect 9214 20272 9220 20284
rect 9272 20272 9278 20324
rect 15286 20312 15292 20324
rect 15247 20284 15292 20312
rect 15286 20272 15292 20284
rect 15344 20272 15350 20324
rect 15764 20312 15792 20343
rect 15838 20340 15844 20392
rect 15896 20380 15902 20392
rect 17221 20383 17279 20389
rect 17221 20380 17233 20383
rect 15896 20352 17233 20380
rect 15896 20340 15902 20352
rect 17221 20349 17233 20352
rect 17267 20349 17279 20383
rect 17788 20380 17816 20420
rect 17957 20417 17969 20451
rect 18003 20417 18015 20451
rect 17957 20411 18015 20417
rect 18601 20451 18659 20457
rect 18601 20417 18613 20451
rect 18647 20448 18659 20451
rect 18874 20448 18880 20460
rect 18647 20420 18880 20448
rect 18647 20417 18659 20420
rect 18601 20411 18659 20417
rect 18874 20408 18880 20420
rect 18932 20408 18938 20460
rect 18969 20451 19027 20457
rect 18969 20417 18981 20451
rect 19015 20417 19027 20451
rect 19076 20448 19104 20488
rect 19426 20476 19432 20528
rect 19484 20516 19490 20528
rect 20456 20525 20484 20556
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 21177 20587 21235 20593
rect 21177 20584 21189 20587
rect 20772 20556 21189 20584
rect 20772 20544 20778 20556
rect 21177 20553 21189 20556
rect 21223 20584 21235 20587
rect 22649 20587 22707 20593
rect 22649 20584 22661 20587
rect 21223 20556 22661 20584
rect 21223 20553 21235 20556
rect 21177 20547 21235 20553
rect 22649 20553 22661 20556
rect 22695 20553 22707 20587
rect 22649 20547 22707 20553
rect 22741 20587 22799 20593
rect 22741 20553 22753 20587
rect 22787 20584 22799 20587
rect 23566 20584 23572 20596
rect 22787 20556 23572 20584
rect 22787 20553 22799 20556
rect 22741 20547 22799 20553
rect 23566 20544 23572 20556
rect 23624 20544 23630 20596
rect 25774 20544 25780 20596
rect 25832 20584 25838 20596
rect 25961 20587 26019 20593
rect 25961 20584 25973 20587
rect 25832 20556 25973 20584
rect 25832 20544 25838 20556
rect 25961 20553 25973 20556
rect 26007 20553 26019 20587
rect 28258 20584 28264 20596
rect 28219 20556 28264 20584
rect 25961 20547 26019 20553
rect 28258 20544 28264 20556
rect 28316 20544 28322 20596
rect 29362 20584 29368 20596
rect 29323 20556 29368 20584
rect 29362 20544 29368 20556
rect 29420 20544 29426 20596
rect 30009 20587 30067 20593
rect 30009 20553 30021 20587
rect 30055 20584 30067 20587
rect 31294 20584 31300 20596
rect 30055 20556 31300 20584
rect 30055 20553 30067 20556
rect 30009 20547 30067 20553
rect 31294 20544 31300 20556
rect 31352 20544 31358 20596
rect 32766 20544 32772 20596
rect 32824 20584 32830 20596
rect 32861 20587 32919 20593
rect 32861 20584 32873 20587
rect 32824 20556 32873 20584
rect 32824 20544 32830 20556
rect 32861 20553 32873 20556
rect 32907 20553 32919 20587
rect 32861 20547 32919 20553
rect 33965 20587 34023 20593
rect 33965 20553 33977 20587
rect 34011 20553 34023 20587
rect 33965 20547 34023 20553
rect 36449 20587 36507 20593
rect 36449 20553 36461 20587
rect 36495 20584 36507 20587
rect 37274 20584 37280 20596
rect 36495 20556 37280 20584
rect 36495 20553 36507 20556
rect 36449 20547 36507 20553
rect 20441 20519 20499 20525
rect 19484 20488 19932 20516
rect 19484 20476 19490 20488
rect 19904 20457 19932 20488
rect 20441 20485 20453 20519
rect 20487 20516 20499 20519
rect 20990 20516 20996 20528
rect 20487 20488 20996 20516
rect 20487 20485 20499 20488
rect 20441 20479 20499 20485
rect 20990 20476 20996 20488
rect 21048 20476 21054 20528
rect 22094 20476 22100 20528
rect 22152 20516 22158 20528
rect 26418 20516 26424 20528
rect 22152 20488 26424 20516
rect 22152 20476 22158 20488
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 19076 20420 19717 20448
rect 18969 20411 19027 20417
rect 19705 20417 19717 20420
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 19889 20451 19947 20457
rect 19889 20417 19901 20451
rect 19935 20417 19947 20451
rect 24581 20451 24639 20457
rect 24581 20448 24593 20451
rect 19889 20411 19947 20417
rect 24044 20420 24593 20448
rect 18506 20380 18512 20392
rect 17788 20352 18512 20380
rect 17221 20343 17279 20349
rect 18506 20340 18512 20352
rect 18564 20380 18570 20392
rect 18984 20380 19012 20411
rect 18564 20352 19012 20380
rect 19061 20383 19119 20389
rect 18564 20340 18570 20352
rect 19061 20349 19073 20383
rect 19107 20380 19119 20383
rect 19150 20380 19156 20392
rect 19107 20352 19156 20380
rect 19107 20349 19119 20352
rect 19061 20343 19119 20349
rect 19150 20340 19156 20352
rect 19208 20340 19214 20392
rect 22186 20340 22192 20392
rect 22244 20380 22250 20392
rect 22830 20380 22836 20392
rect 22244 20352 22836 20380
rect 22244 20340 22250 20352
rect 22830 20340 22836 20352
rect 22888 20340 22894 20392
rect 16758 20312 16764 20324
rect 15764 20284 16764 20312
rect 16758 20272 16764 20284
rect 16816 20312 16822 20324
rect 18138 20312 18144 20324
rect 16816 20284 18144 20312
rect 16816 20272 16822 20284
rect 18138 20272 18144 20284
rect 18196 20272 18202 20324
rect 19886 20312 19892 20324
rect 19076 20284 19892 20312
rect 5534 20244 5540 20256
rect 5495 20216 5540 20244
rect 5534 20204 5540 20216
rect 5592 20204 5598 20256
rect 10229 20247 10287 20253
rect 10229 20213 10241 20247
rect 10275 20244 10287 20247
rect 10594 20244 10600 20256
rect 10275 20216 10600 20244
rect 10275 20213 10287 20216
rect 10229 20207 10287 20213
rect 10594 20204 10600 20216
rect 10652 20204 10658 20256
rect 10778 20244 10784 20256
rect 10739 20216 10784 20244
rect 10778 20204 10784 20216
rect 10836 20204 10842 20256
rect 14826 20244 14832 20256
rect 14787 20216 14832 20244
rect 14826 20204 14832 20216
rect 14884 20204 14890 20256
rect 16114 20204 16120 20256
rect 16172 20244 16178 20256
rect 16669 20247 16727 20253
rect 16669 20244 16681 20247
rect 16172 20216 16681 20244
rect 16172 20204 16178 20216
rect 16669 20213 16681 20216
rect 16715 20213 16727 20247
rect 16669 20207 16727 20213
rect 16942 20204 16948 20256
rect 17000 20244 17006 20256
rect 19076 20244 19104 20284
rect 19886 20272 19892 20284
rect 19944 20312 19950 20324
rect 20898 20312 20904 20324
rect 19944 20284 20904 20312
rect 19944 20272 19950 20284
rect 20898 20272 20904 20284
rect 20956 20272 20962 20324
rect 19242 20244 19248 20256
rect 17000 20216 19104 20244
rect 19203 20216 19248 20244
rect 17000 20204 17006 20216
rect 19242 20204 19248 20216
rect 19300 20204 19306 20256
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 19705 20247 19763 20253
rect 19705 20244 19717 20247
rect 19392 20216 19717 20244
rect 19392 20204 19398 20216
rect 19705 20213 19717 20216
rect 19751 20213 19763 20247
rect 22278 20244 22284 20256
rect 22239 20216 22284 20244
rect 19705 20207 19763 20213
rect 22278 20204 22284 20216
rect 22336 20204 22342 20256
rect 23382 20204 23388 20256
rect 23440 20244 23446 20256
rect 24044 20253 24072 20420
rect 24581 20417 24593 20420
rect 24627 20448 24639 20451
rect 24762 20448 24768 20460
rect 24627 20420 24768 20448
rect 24627 20417 24639 20420
rect 24581 20411 24639 20417
rect 24762 20408 24768 20420
rect 24820 20408 24826 20460
rect 25516 20457 25544 20488
rect 26418 20476 26424 20488
rect 26476 20476 26482 20528
rect 32214 20476 32220 20528
rect 32272 20516 32278 20528
rect 32677 20519 32735 20525
rect 32677 20516 32689 20519
rect 32272 20488 32689 20516
rect 32272 20476 32278 20488
rect 32677 20485 32689 20488
rect 32723 20516 32735 20519
rect 33594 20516 33600 20528
rect 32723 20488 33600 20516
rect 32723 20485 32735 20488
rect 32677 20479 32735 20485
rect 33594 20476 33600 20488
rect 33652 20476 33658 20528
rect 33980 20516 34008 20547
rect 37274 20544 37280 20556
rect 37332 20544 37338 20596
rect 40126 20544 40132 20596
rect 40184 20584 40190 20596
rect 40589 20587 40647 20593
rect 40589 20584 40601 20587
rect 40184 20556 40601 20584
rect 40184 20544 40190 20556
rect 40589 20553 40601 20556
rect 40635 20553 40647 20587
rect 41230 20584 41236 20596
rect 41191 20556 41236 20584
rect 40589 20547 40647 20553
rect 41230 20544 41236 20556
rect 41288 20544 41294 20596
rect 41325 20587 41383 20593
rect 41325 20553 41337 20587
rect 41371 20584 41383 20587
rect 42521 20587 42579 20593
rect 41371 20556 41736 20584
rect 41371 20553 41383 20556
rect 41325 20547 41383 20553
rect 34670 20519 34728 20525
rect 34670 20516 34682 20519
rect 33980 20488 34682 20516
rect 34670 20485 34682 20488
rect 34716 20485 34728 20519
rect 34670 20479 34728 20485
rect 37550 20476 37556 20528
rect 37608 20516 37614 20528
rect 37645 20519 37703 20525
rect 37645 20516 37657 20519
rect 37608 20488 37657 20516
rect 37608 20476 37614 20488
rect 37645 20485 37657 20488
rect 37691 20516 37703 20519
rect 38105 20519 38163 20525
rect 38105 20516 38117 20519
rect 37691 20488 38117 20516
rect 37691 20485 37703 20488
rect 37645 20479 37703 20485
rect 38105 20485 38117 20488
rect 38151 20485 38163 20519
rect 38105 20479 38163 20485
rect 25501 20451 25559 20457
rect 25501 20417 25513 20451
rect 25547 20417 25559 20451
rect 25501 20411 25559 20417
rect 27893 20451 27951 20457
rect 27893 20417 27905 20451
rect 27939 20448 27951 20451
rect 29638 20448 29644 20460
rect 27939 20420 29644 20448
rect 27939 20417 27951 20420
rect 27893 20411 27951 20417
rect 29638 20408 29644 20420
rect 29696 20408 29702 20460
rect 29733 20451 29791 20457
rect 29733 20417 29745 20451
rect 29779 20448 29791 20451
rect 30098 20448 30104 20460
rect 29779 20420 30104 20448
rect 29779 20417 29791 20420
rect 29733 20411 29791 20417
rect 30098 20408 30104 20420
rect 30156 20408 30162 20460
rect 32490 20448 32496 20460
rect 32451 20420 32496 20448
rect 32490 20408 32496 20420
rect 32548 20408 32554 20460
rect 33778 20448 33784 20460
rect 33739 20420 33784 20448
rect 33778 20408 33784 20420
rect 33836 20408 33842 20460
rect 36262 20448 36268 20460
rect 36223 20420 36268 20448
rect 36262 20408 36268 20420
rect 36320 20408 36326 20460
rect 40034 20448 40040 20460
rect 39995 20420 40040 20448
rect 40034 20408 40040 20420
rect 40092 20408 40098 20460
rect 40129 20451 40187 20457
rect 40129 20417 40141 20451
rect 40175 20417 40187 20451
rect 40310 20448 40316 20460
rect 40271 20420 40316 20448
rect 40129 20411 40187 20417
rect 25041 20383 25099 20389
rect 25041 20349 25053 20383
rect 25087 20380 25099 20383
rect 25958 20380 25964 20392
rect 25087 20352 25964 20380
rect 25087 20349 25099 20352
rect 25041 20343 25099 20349
rect 25958 20340 25964 20352
rect 26016 20340 26022 20392
rect 27338 20340 27344 20392
rect 27396 20380 27402 20392
rect 27801 20383 27859 20389
rect 27801 20380 27813 20383
rect 27396 20352 27813 20380
rect 27396 20340 27402 20352
rect 27801 20349 27813 20352
rect 27847 20349 27859 20383
rect 29822 20380 29828 20392
rect 29783 20352 29828 20380
rect 27801 20343 27859 20349
rect 29822 20340 29828 20352
rect 29880 20340 29886 20392
rect 33502 20340 33508 20392
rect 33560 20380 33566 20392
rect 34425 20383 34483 20389
rect 34425 20380 34437 20383
rect 33560 20352 34437 20380
rect 33560 20340 33566 20352
rect 34425 20349 34437 20352
rect 34471 20349 34483 20383
rect 34425 20343 34483 20349
rect 38933 20383 38991 20389
rect 38933 20349 38945 20383
rect 38979 20380 38991 20383
rect 39298 20380 39304 20392
rect 38979 20352 39304 20380
rect 38979 20349 38991 20352
rect 38933 20343 38991 20349
rect 39298 20340 39304 20352
rect 39356 20340 39362 20392
rect 40144 20312 40172 20411
rect 40310 20408 40316 20420
rect 40368 20408 40374 20460
rect 40402 20408 40408 20460
rect 40460 20448 40466 20460
rect 40460 20420 40505 20448
rect 40460 20408 40466 20420
rect 41708 20380 41736 20556
rect 42521 20553 42533 20587
rect 42567 20584 42579 20587
rect 42610 20584 42616 20596
rect 42567 20556 42616 20584
rect 42567 20553 42579 20556
rect 42521 20547 42579 20553
rect 42610 20544 42616 20556
rect 42668 20544 42674 20596
rect 41785 20519 41843 20525
rect 41785 20485 41797 20519
rect 41831 20516 41843 20519
rect 43806 20516 43812 20528
rect 41831 20488 43812 20516
rect 41831 20485 41843 20488
rect 41785 20479 41843 20485
rect 43806 20476 43812 20488
rect 43864 20476 43870 20528
rect 43901 20519 43959 20525
rect 43901 20485 43913 20519
rect 43947 20516 43959 20519
rect 44174 20516 44180 20528
rect 43947 20488 44180 20516
rect 43947 20485 43959 20488
rect 43901 20479 43959 20485
rect 44174 20476 44180 20488
rect 44232 20476 44238 20528
rect 42426 20448 42432 20460
rect 42387 20420 42432 20448
rect 42426 20408 42432 20420
rect 42484 20408 42490 20460
rect 42702 20448 42708 20460
rect 42663 20420 42708 20448
rect 42702 20408 42708 20420
rect 42760 20408 42766 20460
rect 45002 20408 45008 20460
rect 45060 20408 45066 20460
rect 45186 20408 45192 20460
rect 45244 20448 45250 20460
rect 45833 20451 45891 20457
rect 45833 20448 45845 20451
rect 45244 20420 45845 20448
rect 45244 20408 45250 20420
rect 45833 20417 45845 20420
rect 45879 20417 45891 20451
rect 46106 20448 46112 20460
rect 46067 20420 46112 20448
rect 45833 20411 45891 20417
rect 46106 20408 46112 20420
rect 46164 20408 46170 20460
rect 41708 20352 43300 20380
rect 40144 20284 41552 20312
rect 24029 20247 24087 20253
rect 24029 20244 24041 20247
rect 23440 20216 24041 20244
rect 23440 20204 23446 20216
rect 24029 20213 24041 20216
rect 24075 20213 24087 20247
rect 24029 20207 24087 20213
rect 24765 20247 24823 20253
rect 24765 20213 24777 20247
rect 24811 20244 24823 20247
rect 24946 20244 24952 20256
rect 24811 20216 24952 20244
rect 24811 20213 24823 20216
rect 24765 20207 24823 20213
rect 24946 20204 24952 20216
rect 25004 20204 25010 20256
rect 25774 20244 25780 20256
rect 25735 20216 25780 20244
rect 25774 20204 25780 20216
rect 25832 20204 25838 20256
rect 27798 20204 27804 20256
rect 27856 20244 27862 20256
rect 28442 20244 28448 20256
rect 27856 20216 28448 20244
rect 27856 20204 27862 20216
rect 28442 20204 28448 20216
rect 28500 20244 28506 20256
rect 28721 20247 28779 20253
rect 28721 20244 28733 20247
rect 28500 20216 28733 20244
rect 28500 20204 28506 20216
rect 28721 20213 28733 20216
rect 28767 20213 28779 20247
rect 35802 20244 35808 20256
rect 35763 20216 35808 20244
rect 28721 20207 28779 20213
rect 35802 20204 35808 20216
rect 35860 20204 35866 20256
rect 41049 20247 41107 20253
rect 41049 20213 41061 20247
rect 41095 20244 41107 20247
rect 41414 20244 41420 20256
rect 41095 20216 41420 20244
rect 41095 20213 41107 20216
rect 41049 20207 41107 20213
rect 41414 20204 41420 20216
rect 41472 20204 41478 20256
rect 41524 20244 41552 20284
rect 41598 20272 41604 20324
rect 41656 20312 41662 20324
rect 41785 20315 41843 20321
rect 41785 20312 41797 20315
rect 41656 20284 41797 20312
rect 41656 20272 41662 20284
rect 41785 20281 41797 20284
rect 41831 20281 41843 20315
rect 43272 20312 43300 20352
rect 43346 20340 43352 20392
rect 43404 20380 43410 20392
rect 43625 20383 43683 20389
rect 43625 20380 43637 20383
rect 43404 20352 43637 20380
rect 43404 20340 43410 20352
rect 43625 20349 43637 20352
rect 43671 20349 43683 20383
rect 44266 20380 44272 20392
rect 43625 20343 43683 20349
rect 43732 20352 44272 20380
rect 43732 20312 43760 20352
rect 44266 20340 44272 20352
rect 44324 20380 44330 20392
rect 44910 20380 44916 20392
rect 44324 20352 44916 20380
rect 44324 20340 44330 20352
rect 44910 20340 44916 20352
rect 44968 20380 44974 20392
rect 45373 20383 45431 20389
rect 45373 20380 45385 20383
rect 44968 20352 45385 20380
rect 44968 20340 44974 20352
rect 45373 20349 45385 20352
rect 45419 20349 45431 20383
rect 45373 20343 45431 20349
rect 41785 20275 41843 20281
rect 41892 20284 43208 20312
rect 43272 20284 43760 20312
rect 41892 20244 41920 20284
rect 41524 20216 41920 20244
rect 42889 20247 42947 20253
rect 42889 20213 42901 20247
rect 42935 20244 42947 20247
rect 43070 20244 43076 20256
rect 42935 20216 43076 20244
rect 42935 20213 42947 20216
rect 42889 20207 42947 20213
rect 43070 20204 43076 20216
rect 43128 20204 43134 20256
rect 43180 20244 43208 20284
rect 45186 20244 45192 20256
rect 43180 20216 45192 20244
rect 45186 20204 45192 20216
rect 45244 20204 45250 20256
rect 46845 20247 46903 20253
rect 46845 20213 46857 20247
rect 46891 20244 46903 20247
rect 55122 20244 55128 20256
rect 46891 20216 55128 20244
rect 46891 20213 46903 20216
rect 46845 20207 46903 20213
rect 55122 20204 55128 20216
rect 55180 20244 55186 20256
rect 60550 20244 60556 20256
rect 55180 20216 60556 20244
rect 55180 20204 55186 20216
rect 60550 20204 60556 20216
rect 60608 20204 60614 20256
rect 1104 20154 68816 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 65654 20154
rect 65706 20102 65718 20154
rect 65770 20102 65782 20154
rect 65834 20102 65846 20154
rect 65898 20102 65910 20154
rect 65962 20102 68816 20154
rect 1104 20080 68816 20102
rect 6181 20043 6239 20049
rect 6181 20040 6193 20043
rect 5736 20012 6193 20040
rect 5736 19916 5764 20012
rect 6181 20009 6193 20012
rect 6227 20009 6239 20043
rect 6181 20003 6239 20009
rect 7653 20043 7711 20049
rect 7653 20009 7665 20043
rect 7699 20040 7711 20043
rect 7926 20040 7932 20052
rect 7699 20012 7932 20040
rect 7699 20009 7711 20012
rect 7653 20003 7711 20009
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 11974 20040 11980 20052
rect 11935 20012 11980 20040
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 12158 20000 12164 20052
rect 12216 20040 12222 20052
rect 22186 20040 22192 20052
rect 12216 20012 22192 20040
rect 12216 20000 12222 20012
rect 22186 20000 22192 20012
rect 22244 20000 22250 20052
rect 22462 20040 22468 20052
rect 22423 20012 22468 20040
rect 22462 20000 22468 20012
rect 22520 20000 22526 20052
rect 23293 20043 23351 20049
rect 23293 20009 23305 20043
rect 23339 20040 23351 20043
rect 23750 20040 23756 20052
rect 23339 20012 23756 20040
rect 23339 20009 23351 20012
rect 23293 20003 23351 20009
rect 23750 20000 23756 20012
rect 23808 20000 23814 20052
rect 27338 20040 27344 20052
rect 27299 20012 27344 20040
rect 27338 20000 27344 20012
rect 27396 20000 27402 20052
rect 31662 20000 31668 20052
rect 31720 20040 31726 20052
rect 31757 20043 31815 20049
rect 31757 20040 31769 20043
rect 31720 20012 31769 20040
rect 31720 20000 31726 20012
rect 31757 20009 31769 20012
rect 31803 20009 31815 20043
rect 31757 20003 31815 20009
rect 33778 20000 33784 20052
rect 33836 20040 33842 20052
rect 34885 20043 34943 20049
rect 34885 20040 34897 20043
rect 33836 20012 34897 20040
rect 33836 20000 33842 20012
rect 34885 20009 34897 20012
rect 34931 20009 34943 20043
rect 37918 20040 37924 20052
rect 34885 20003 34943 20009
rect 35084 20012 37924 20040
rect 8294 19972 8300 19984
rect 7852 19944 8300 19972
rect 5077 19907 5135 19913
rect 5077 19873 5089 19907
rect 5123 19904 5135 19907
rect 5718 19904 5724 19916
rect 5123 19876 5724 19904
rect 5123 19873 5135 19876
rect 5077 19867 5135 19873
rect 5718 19864 5724 19876
rect 5776 19864 5782 19916
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19836 5043 19839
rect 5534 19836 5540 19848
rect 5031 19808 5540 19836
rect 5031 19805 5043 19808
rect 4985 19799 5043 19805
rect 5534 19796 5540 19808
rect 5592 19796 5598 19848
rect 6089 19839 6147 19845
rect 6089 19805 6101 19839
rect 6135 19836 6147 19839
rect 7098 19836 7104 19848
rect 6135 19808 7104 19836
rect 6135 19805 6147 19808
rect 6089 19799 6147 19805
rect 7098 19796 7104 19808
rect 7156 19796 7162 19848
rect 7852 19845 7880 19944
rect 8294 19932 8300 19944
rect 8352 19932 8358 19984
rect 14182 19972 14188 19984
rect 14143 19944 14188 19972
rect 14182 19932 14188 19944
rect 14240 19932 14246 19984
rect 16669 19975 16727 19981
rect 16669 19941 16681 19975
rect 16715 19941 16727 19975
rect 17126 19972 17132 19984
rect 17087 19944 17132 19972
rect 16669 19935 16727 19941
rect 8478 19904 8484 19916
rect 8036 19876 8484 19904
rect 8036 19845 8064 19876
rect 8478 19864 8484 19876
rect 8536 19904 8542 19916
rect 8941 19907 8999 19913
rect 8941 19904 8953 19907
rect 8536 19876 8953 19904
rect 8536 19864 8542 19876
rect 8941 19873 8953 19876
rect 8987 19873 8999 19907
rect 8941 19867 8999 19873
rect 11146 19864 11152 19916
rect 11204 19904 11210 19916
rect 12250 19904 12256 19916
rect 11204 19876 12256 19904
rect 11204 19864 11210 19876
rect 12250 19864 12256 19876
rect 12308 19904 12314 19916
rect 12529 19907 12587 19913
rect 12529 19904 12541 19907
rect 12308 19876 12541 19904
rect 12308 19864 12314 19876
rect 12529 19873 12541 19876
rect 12575 19873 12587 19907
rect 12529 19867 12587 19873
rect 14458 19864 14464 19916
rect 14516 19904 14522 19916
rect 15289 19907 15347 19913
rect 15289 19904 15301 19907
rect 14516 19876 15301 19904
rect 14516 19864 14522 19876
rect 15289 19873 15301 19876
rect 15335 19873 15347 19907
rect 16684 19904 16712 19935
rect 17126 19932 17132 19944
rect 17184 19932 17190 19984
rect 18046 19972 18052 19984
rect 18007 19944 18052 19972
rect 18046 19932 18052 19944
rect 18104 19932 18110 19984
rect 18782 19932 18788 19984
rect 18840 19972 18846 19984
rect 20806 19972 20812 19984
rect 18840 19944 20812 19972
rect 18840 19932 18846 19944
rect 19613 19907 19671 19913
rect 16684 19876 18552 19904
rect 15289 19867 15347 19873
rect 18524 19848 18552 19876
rect 18616 19876 19288 19904
rect 7837 19839 7895 19845
rect 7837 19805 7849 19839
rect 7883 19805 7895 19839
rect 7837 19799 7895 19805
rect 8021 19839 8079 19845
rect 8021 19805 8033 19839
rect 8067 19805 8079 19839
rect 8021 19799 8079 19805
rect 8113 19839 8171 19845
rect 8113 19805 8125 19839
rect 8159 19836 8171 19839
rect 8202 19836 8208 19848
rect 8159 19808 8208 19836
rect 8159 19805 8171 19808
rect 8113 19799 8171 19805
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19836 9183 19839
rect 9490 19836 9496 19848
rect 9171 19808 9496 19836
rect 9171 19805 9183 19808
rect 9125 19799 9183 19805
rect 9490 19796 9496 19808
rect 9548 19796 9554 19848
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19836 10195 19839
rect 11514 19836 11520 19848
rect 10183 19808 11520 19836
rect 10183 19805 10195 19808
rect 10137 19799 10195 19805
rect 4614 19728 4620 19780
rect 4672 19768 4678 19780
rect 10152 19768 10180 19799
rect 11514 19796 11520 19808
rect 11572 19796 11578 19848
rect 12342 19796 12348 19848
rect 12400 19836 12406 19848
rect 12437 19839 12495 19845
rect 12437 19836 12449 19839
rect 12400 19808 12449 19836
rect 12400 19796 12406 19808
rect 12437 19805 12449 19808
rect 12483 19805 12495 19839
rect 14826 19836 14832 19848
rect 14787 19808 14832 19836
rect 12437 19799 12495 19805
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 18506 19836 18512 19848
rect 18467 19808 18512 19836
rect 18506 19796 18512 19808
rect 18564 19796 18570 19848
rect 4672 19740 10180 19768
rect 10404 19771 10462 19777
rect 4672 19728 4678 19740
rect 10404 19737 10416 19771
rect 10450 19768 10462 19771
rect 10778 19768 10784 19780
rect 10450 19740 10784 19768
rect 10450 19737 10462 19740
rect 10404 19731 10462 19737
rect 10778 19728 10784 19740
rect 10836 19728 10842 19780
rect 15556 19771 15614 19777
rect 15556 19737 15568 19771
rect 15602 19768 15614 19771
rect 15930 19768 15936 19780
rect 15602 19740 15936 19768
rect 15602 19737 15614 19740
rect 15556 19731 15614 19737
rect 15930 19728 15936 19740
rect 15988 19728 15994 19780
rect 18616 19768 18644 19876
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 19150 19836 19156 19848
rect 18739 19808 19156 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 19150 19796 19156 19808
rect 19208 19796 19214 19848
rect 19260 19836 19288 19876
rect 19613 19873 19625 19907
rect 19659 19904 19671 19907
rect 19978 19904 19984 19916
rect 19659 19876 19984 19904
rect 19659 19873 19671 19876
rect 19613 19867 19671 19873
rect 19978 19864 19984 19876
rect 20036 19864 20042 19916
rect 19705 19839 19763 19845
rect 19705 19836 19717 19839
rect 19260 19808 19717 19836
rect 19705 19805 19717 19808
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 18524 19740 18644 19768
rect 5353 19703 5411 19709
rect 5353 19669 5365 19703
rect 5399 19700 5411 19703
rect 5442 19700 5448 19712
rect 5399 19672 5448 19700
rect 5399 19669 5411 19672
rect 5353 19663 5411 19669
rect 5442 19660 5448 19672
rect 5500 19660 5506 19712
rect 6546 19700 6552 19712
rect 6507 19672 6552 19700
rect 6546 19660 6552 19672
rect 6604 19660 6610 19712
rect 7098 19700 7104 19712
rect 7059 19672 7104 19700
rect 7098 19660 7104 19672
rect 7156 19660 7162 19712
rect 9030 19660 9036 19712
rect 9088 19700 9094 19712
rect 9306 19700 9312 19712
rect 9088 19672 9312 19700
rect 9088 19660 9094 19672
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 11054 19660 11060 19712
rect 11112 19700 11118 19712
rect 11517 19703 11575 19709
rect 11517 19700 11529 19703
rect 11112 19672 11529 19700
rect 11112 19660 11118 19672
rect 11517 19669 11529 19672
rect 11563 19700 11575 19703
rect 12345 19703 12403 19709
rect 12345 19700 12357 19703
rect 11563 19672 12357 19700
rect 11563 19669 11575 19672
rect 11517 19663 11575 19669
rect 12345 19669 12357 19672
rect 12391 19669 12403 19703
rect 14642 19700 14648 19712
rect 14603 19672 14648 19700
rect 12345 19663 12403 19669
rect 14642 19660 14648 19672
rect 14700 19660 14706 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 18524 19700 18552 19740
rect 18874 19728 18880 19780
rect 18932 19768 18938 19780
rect 19518 19768 19524 19780
rect 18932 19740 19524 19768
rect 18932 19728 18938 19740
rect 19518 19728 19524 19740
rect 19576 19728 19582 19780
rect 18690 19700 18696 19712
rect 15528 19672 18552 19700
rect 18651 19672 18696 19700
rect 15528 19660 15534 19672
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 19426 19700 19432 19712
rect 19387 19672 19432 19700
rect 19426 19660 19432 19672
rect 19484 19660 19490 19712
rect 19720 19700 19748 19799
rect 19794 19796 19800 19848
rect 19852 19836 19858 19848
rect 20732 19845 20760 19944
rect 20806 19932 20812 19944
rect 20864 19932 20870 19984
rect 20898 19932 20904 19984
rect 20956 19972 20962 19984
rect 21177 19975 21235 19981
rect 21177 19972 21189 19975
rect 20956 19944 21189 19972
rect 20956 19932 20962 19944
rect 21177 19941 21189 19944
rect 21223 19941 21235 19975
rect 26050 19972 26056 19984
rect 26011 19944 26056 19972
rect 21177 19935 21235 19941
rect 26050 19932 26056 19944
rect 26108 19972 26114 19984
rect 30469 19975 30527 19981
rect 26108 19944 27108 19972
rect 26108 19932 26114 19944
rect 25774 19904 25780 19916
rect 25735 19876 25780 19904
rect 25774 19864 25780 19876
rect 25832 19864 25838 19916
rect 20073 19839 20131 19845
rect 20073 19836 20085 19839
rect 19852 19808 20085 19836
rect 19852 19796 19858 19808
rect 20073 19805 20085 19808
rect 20119 19836 20131 19839
rect 20533 19839 20591 19845
rect 20533 19836 20545 19839
rect 20119 19808 20545 19836
rect 20119 19805 20131 19808
rect 20073 19799 20131 19805
rect 20533 19805 20545 19808
rect 20579 19805 20591 19839
rect 20533 19799 20591 19805
rect 20717 19839 20775 19845
rect 20717 19805 20729 19839
rect 20763 19805 20775 19839
rect 22278 19836 22284 19848
rect 22239 19808 22284 19836
rect 20717 19799 20775 19805
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 23014 19796 23020 19848
rect 23072 19836 23078 19848
rect 23109 19839 23167 19845
rect 23109 19836 23121 19839
rect 23072 19808 23121 19836
rect 23072 19796 23078 19808
rect 23109 19805 23121 19808
rect 23155 19805 23167 19839
rect 23109 19799 23167 19805
rect 25685 19839 25743 19845
rect 25685 19805 25697 19839
rect 25731 19836 25743 19839
rect 26234 19836 26240 19848
rect 25731 19808 26240 19836
rect 25731 19805 25743 19808
rect 25685 19799 25743 19805
rect 26234 19796 26240 19808
rect 26292 19796 26298 19848
rect 27080 19845 27108 19944
rect 30469 19941 30481 19975
rect 30515 19972 30527 19975
rect 32490 19972 32496 19984
rect 30515 19944 32496 19972
rect 30515 19941 30527 19944
rect 30469 19935 30527 19941
rect 32490 19932 32496 19944
rect 32548 19932 32554 19984
rect 27154 19864 27160 19916
rect 27212 19904 27218 19916
rect 27338 19904 27344 19916
rect 27212 19876 27344 19904
rect 27212 19864 27218 19876
rect 27338 19864 27344 19876
rect 27396 19864 27402 19916
rect 29270 19864 29276 19916
rect 29328 19904 29334 19916
rect 29822 19904 29828 19916
rect 29328 19876 29828 19904
rect 29328 19864 29334 19876
rect 29822 19864 29828 19876
rect 29880 19904 29886 19916
rect 30009 19907 30067 19913
rect 30009 19904 30021 19907
rect 29880 19876 30021 19904
rect 29880 19864 29886 19876
rect 30009 19873 30021 19876
rect 30055 19873 30067 19907
rect 30009 19867 30067 19873
rect 32125 19907 32183 19913
rect 32125 19873 32137 19907
rect 32171 19904 32183 19907
rect 35084 19904 35112 20012
rect 37918 20000 37924 20012
rect 37976 20000 37982 20052
rect 40034 20040 40040 20052
rect 39995 20012 40040 20040
rect 40034 20000 40040 20012
rect 40092 20000 40098 20052
rect 41414 20000 41420 20052
rect 41472 20040 41478 20052
rect 41601 20043 41659 20049
rect 41472 20012 41517 20040
rect 41472 20000 41478 20012
rect 41601 20009 41613 20043
rect 41647 20040 41659 20043
rect 42702 20040 42708 20052
rect 41647 20012 42708 20040
rect 41647 20009 41659 20012
rect 41601 20003 41659 20009
rect 42702 20000 42708 20012
rect 42760 20000 42766 20052
rect 45465 20043 45523 20049
rect 45465 20009 45477 20043
rect 45511 20040 45523 20043
rect 45646 20040 45652 20052
rect 45511 20012 45652 20040
rect 45511 20009 45523 20012
rect 45465 20003 45523 20009
rect 45646 20000 45652 20012
rect 45704 20000 45710 20052
rect 37829 19975 37887 19981
rect 37829 19941 37841 19975
rect 37875 19972 37887 19975
rect 39942 19972 39948 19984
rect 37875 19944 39948 19972
rect 37875 19941 37887 19944
rect 37829 19935 37887 19941
rect 39942 19932 39948 19944
rect 40000 19932 40006 19984
rect 40310 19972 40316 19984
rect 40236 19944 40316 19972
rect 35434 19904 35440 19916
rect 32171 19876 35112 19904
rect 35395 19876 35440 19904
rect 32171 19873 32183 19876
rect 32125 19867 32183 19873
rect 35434 19864 35440 19876
rect 35492 19864 35498 19916
rect 37553 19907 37611 19913
rect 37553 19873 37565 19907
rect 37599 19904 37611 19907
rect 38010 19904 38016 19916
rect 37599 19876 38016 19904
rect 37599 19873 37611 19876
rect 37553 19867 37611 19873
rect 38010 19864 38016 19876
rect 38068 19864 38074 19916
rect 40236 19913 40264 19944
rect 40310 19932 40316 19944
rect 40368 19932 40374 19984
rect 43806 19932 43812 19984
rect 43864 19972 43870 19984
rect 45094 19972 45100 19984
rect 43864 19944 45100 19972
rect 43864 19932 43870 19944
rect 45094 19932 45100 19944
rect 45152 19972 45158 19984
rect 45281 19975 45339 19981
rect 45281 19972 45293 19975
rect 45152 19944 45293 19972
rect 45152 19932 45158 19944
rect 45281 19941 45293 19944
rect 45327 19941 45339 19975
rect 45281 19935 45339 19941
rect 40221 19907 40279 19913
rect 40221 19873 40233 19907
rect 40267 19873 40279 19907
rect 42794 19904 42800 19916
rect 42755 19876 42800 19904
rect 40221 19867 40279 19873
rect 42794 19864 42800 19876
rect 42852 19864 42858 19916
rect 44910 19864 44916 19916
rect 44968 19904 44974 19916
rect 45005 19907 45063 19913
rect 45005 19904 45017 19907
rect 44968 19876 45017 19904
rect 44968 19864 44974 19876
rect 45005 19873 45017 19876
rect 45051 19873 45063 19907
rect 45005 19867 45063 19873
rect 27065 19839 27123 19845
rect 27065 19805 27077 19839
rect 27111 19805 27123 19839
rect 30098 19836 30104 19848
rect 30059 19808 30104 19836
rect 27065 19799 27123 19805
rect 30098 19796 30104 19808
rect 30156 19796 30162 19848
rect 31665 19839 31723 19845
rect 31665 19836 31677 19839
rect 31128 19808 31677 19836
rect 19886 19728 19892 19780
rect 19944 19768 19950 19780
rect 19981 19771 20039 19777
rect 19981 19768 19993 19771
rect 19944 19740 19993 19768
rect 19944 19728 19950 19740
rect 19981 19737 19993 19740
rect 20027 19737 20039 19771
rect 19981 19731 20039 19737
rect 31128 19712 31156 19808
rect 31665 19805 31677 19808
rect 31711 19805 31723 19839
rect 31665 19799 31723 19805
rect 32769 19839 32827 19845
rect 32769 19805 32781 19839
rect 32815 19836 32827 19839
rect 33318 19836 33324 19848
rect 32815 19808 33324 19836
rect 32815 19805 32827 19808
rect 32769 19799 32827 19805
rect 33318 19796 33324 19808
rect 33376 19796 33382 19848
rect 35345 19839 35403 19845
rect 35345 19805 35357 19839
rect 35391 19836 35403 19839
rect 35802 19836 35808 19848
rect 35391 19808 35808 19836
rect 35391 19805 35403 19808
rect 35345 19799 35403 19805
rect 35802 19796 35808 19808
rect 35860 19836 35866 19848
rect 37461 19839 37519 19845
rect 37461 19836 37473 19839
rect 35860 19808 37473 19836
rect 35860 19796 35866 19808
rect 37461 19805 37473 19808
rect 37507 19805 37519 19839
rect 37461 19799 37519 19805
rect 40313 19839 40371 19845
rect 40313 19805 40325 19839
rect 40359 19836 40371 19839
rect 40402 19836 40408 19848
rect 40359 19808 40408 19836
rect 40359 19805 40371 19808
rect 40313 19799 40371 19805
rect 40402 19796 40408 19808
rect 40460 19796 40466 19848
rect 43070 19836 43076 19848
rect 43031 19808 43076 19836
rect 43070 19796 43076 19808
rect 43128 19796 43134 19848
rect 34149 19771 34207 19777
rect 34149 19737 34161 19771
rect 34195 19768 34207 19771
rect 35253 19771 35311 19777
rect 35253 19768 35265 19771
rect 34195 19740 35265 19768
rect 34195 19737 34207 19740
rect 34149 19731 34207 19737
rect 35253 19737 35265 19740
rect 35299 19768 35311 19771
rect 35526 19768 35532 19780
rect 35299 19740 35532 19768
rect 35299 19737 35311 19740
rect 35253 19731 35311 19737
rect 35526 19728 35532 19740
rect 35584 19728 35590 19780
rect 40586 19768 40592 19780
rect 40547 19740 40592 19768
rect 40586 19728 40592 19740
rect 40644 19728 40650 19780
rect 40678 19728 40684 19780
rect 40736 19768 40742 19780
rect 40736 19740 40781 19768
rect 40736 19728 40742 19740
rect 41138 19728 41144 19780
rect 41196 19768 41202 19780
rect 41233 19771 41291 19777
rect 41233 19768 41245 19771
rect 41196 19740 41245 19768
rect 41196 19728 41202 19740
rect 41233 19737 41245 19740
rect 41279 19737 41291 19771
rect 41233 19731 41291 19737
rect 41449 19771 41507 19777
rect 41449 19737 41461 19771
rect 41495 19768 41507 19771
rect 42426 19768 42432 19780
rect 41495 19740 42432 19768
rect 41495 19737 41507 19740
rect 41449 19731 41507 19737
rect 42426 19728 42432 19740
rect 42484 19728 42490 19780
rect 20070 19700 20076 19712
rect 19720 19672 20076 19700
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20622 19700 20628 19712
rect 20583 19672 20628 19700
rect 20622 19660 20628 19672
rect 20680 19660 20686 19712
rect 31110 19700 31116 19712
rect 31071 19672 31116 19700
rect 31110 19660 31116 19672
rect 31168 19660 31174 19712
rect 32490 19660 32496 19712
rect 32548 19700 32554 19712
rect 32585 19703 32643 19709
rect 32585 19700 32597 19703
rect 32548 19672 32597 19700
rect 32548 19660 32554 19672
rect 32585 19669 32597 19672
rect 32631 19669 32643 19703
rect 32585 19663 32643 19669
rect 43622 19660 43628 19712
rect 43680 19700 43686 19712
rect 43809 19703 43867 19709
rect 43809 19700 43821 19703
rect 43680 19672 43821 19700
rect 43680 19660 43686 19672
rect 43809 19669 43821 19672
rect 43855 19669 43867 19703
rect 43809 19663 43867 19669
rect 1104 19610 68816 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 68816 19610
rect 1104 19536 68816 19558
rect 3881 19499 3939 19505
rect 3881 19465 3893 19499
rect 3927 19465 3939 19499
rect 5718 19496 5724 19508
rect 5679 19468 5724 19496
rect 3881 19459 3939 19465
rect 3896 19428 3924 19459
rect 5718 19456 5724 19468
rect 5776 19456 5782 19508
rect 6825 19499 6883 19505
rect 6825 19465 6837 19499
rect 6871 19496 6883 19499
rect 15470 19496 15476 19508
rect 6871 19468 7604 19496
rect 15431 19468 15476 19496
rect 6871 19465 6883 19468
rect 6825 19459 6883 19465
rect 4586 19431 4644 19437
rect 4586 19428 4598 19431
rect 3896 19400 4598 19428
rect 4586 19397 4598 19400
rect 4632 19397 4644 19431
rect 4586 19391 4644 19397
rect 6365 19431 6423 19437
rect 6365 19397 6377 19431
rect 6411 19428 6423 19431
rect 7098 19428 7104 19440
rect 6411 19400 7104 19428
rect 6411 19397 6423 19400
rect 6365 19391 6423 19397
rect 7098 19388 7104 19400
rect 7156 19388 7162 19440
rect 7576 19437 7604 19468
rect 15470 19456 15476 19468
rect 15528 19456 15534 19508
rect 15930 19496 15936 19508
rect 15891 19468 15936 19496
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 20622 19496 20628 19508
rect 19352 19468 20628 19496
rect 7561 19431 7619 19437
rect 7561 19397 7573 19431
rect 7607 19397 7619 19431
rect 7561 19391 7619 19397
rect 14360 19431 14418 19437
rect 14360 19397 14372 19431
rect 14406 19428 14418 19431
rect 14642 19428 14648 19440
rect 14406 19400 14648 19428
rect 14406 19397 14418 19400
rect 14360 19391 14418 19397
rect 14642 19388 14648 19400
rect 14700 19388 14706 19440
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19360 3755 19363
rect 4341 19363 4399 19369
rect 3743 19332 4292 19360
rect 3743 19329 3755 19332
rect 3697 19323 3755 19329
rect 4264 19156 4292 19332
rect 4341 19329 4353 19363
rect 4387 19360 4399 19363
rect 4430 19360 4436 19372
rect 4387 19332 4436 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 6546 19320 6552 19372
rect 6604 19360 6610 19372
rect 7285 19363 7343 19369
rect 7285 19360 7297 19363
rect 6604 19332 7297 19360
rect 6604 19320 6610 19332
rect 7285 19329 7297 19332
rect 7331 19329 7343 19363
rect 7285 19323 7343 19329
rect 7374 19320 7380 19372
rect 7432 19360 7438 19372
rect 8294 19360 8300 19372
rect 7432 19332 7477 19360
rect 7576 19332 8300 19360
rect 7432 19320 7438 19332
rect 5718 19184 5724 19236
rect 5776 19224 5782 19236
rect 7576 19233 7604 19332
rect 8294 19320 8300 19332
rect 8352 19320 8358 19372
rect 10505 19363 10563 19369
rect 10505 19329 10517 19363
rect 10551 19360 10563 19363
rect 11054 19360 11060 19372
rect 10551 19332 11060 19360
rect 10551 19329 10563 19332
rect 10505 19323 10563 19329
rect 11054 19320 11060 19332
rect 11112 19320 11118 19372
rect 11514 19320 11520 19372
rect 11572 19360 11578 19372
rect 14093 19363 14151 19369
rect 14093 19360 14105 19363
rect 11572 19332 14105 19360
rect 11572 19320 11578 19332
rect 14093 19329 14105 19332
rect 14139 19329 14151 19363
rect 16114 19360 16120 19372
rect 16075 19332 16120 19360
rect 14093 19323 14151 19329
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 18782 19360 18788 19372
rect 18743 19332 18788 19360
rect 18782 19320 18788 19332
rect 18840 19320 18846 19372
rect 19352 19360 19380 19468
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 23658 19456 23664 19508
rect 23716 19496 23722 19508
rect 30374 19496 30380 19508
rect 23716 19468 30380 19496
rect 23716 19456 23722 19468
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 31573 19499 31631 19505
rect 31573 19465 31585 19499
rect 31619 19496 31631 19499
rect 31754 19496 31760 19508
rect 31619 19468 31760 19496
rect 31619 19465 31631 19468
rect 31573 19459 31631 19465
rect 31754 19456 31760 19468
rect 31812 19456 31818 19508
rect 33594 19496 33600 19508
rect 33555 19468 33600 19496
rect 33594 19456 33600 19468
rect 33652 19456 33658 19508
rect 40678 19456 40684 19508
rect 40736 19496 40742 19508
rect 40865 19499 40923 19505
rect 40865 19496 40877 19499
rect 40736 19468 40877 19496
rect 40736 19456 40742 19468
rect 40865 19465 40877 19468
rect 40911 19465 40923 19499
rect 45094 19496 45100 19508
rect 45055 19468 45100 19496
rect 40865 19459 40923 19465
rect 45094 19456 45100 19468
rect 45152 19456 45158 19508
rect 19426 19388 19432 19440
rect 19484 19428 19490 19440
rect 19978 19428 19984 19440
rect 19484 19400 19656 19428
rect 19484 19388 19490 19400
rect 19628 19369 19656 19400
rect 19812 19400 19984 19428
rect 19812 19369 19840 19400
rect 19978 19388 19984 19400
rect 20036 19388 20042 19440
rect 20901 19431 20959 19437
rect 20901 19397 20913 19431
rect 20947 19428 20959 19431
rect 20990 19428 20996 19440
rect 20947 19400 20996 19428
rect 20947 19397 20959 19400
rect 20901 19391 20959 19397
rect 20990 19388 20996 19400
rect 21048 19388 21054 19440
rect 22465 19431 22523 19437
rect 22465 19397 22477 19431
rect 22511 19428 22523 19431
rect 22922 19428 22928 19440
rect 22511 19400 22928 19428
rect 22511 19397 22523 19400
rect 22465 19391 22523 19397
rect 22922 19388 22928 19400
rect 22980 19388 22986 19440
rect 25222 19428 25228 19440
rect 23216 19400 25228 19428
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19352 19332 19533 19360
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19329 19671 19363
rect 19613 19323 19671 19329
rect 19797 19363 19855 19369
rect 19797 19329 19809 19363
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19360 19947 19363
rect 20070 19360 20076 19372
rect 19935 19332 20076 19360
rect 19935 19329 19947 19332
rect 19889 19323 19947 19329
rect 9582 19252 9588 19304
rect 9640 19292 9646 19304
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 9640 19264 9689 19292
rect 9640 19252 9646 19264
rect 9677 19261 9689 19264
rect 9723 19261 9735 19295
rect 10594 19292 10600 19304
rect 10555 19264 10600 19292
rect 9677 19255 9735 19261
rect 10594 19252 10600 19264
rect 10652 19252 10658 19304
rect 11072 19292 11100 19320
rect 11609 19295 11667 19301
rect 11609 19292 11621 19295
rect 11072 19264 11621 19292
rect 11609 19261 11621 19264
rect 11655 19261 11667 19295
rect 16758 19292 16764 19304
rect 16719 19264 16764 19292
rect 11609 19255 11667 19261
rect 6641 19227 6699 19233
rect 6641 19224 6653 19227
rect 5776 19196 6653 19224
rect 5776 19184 5782 19196
rect 6641 19193 6653 19196
rect 6687 19193 6699 19227
rect 6641 19187 6699 19193
rect 7561 19227 7619 19233
rect 7561 19193 7573 19227
rect 7607 19193 7619 19227
rect 7561 19187 7619 19193
rect 4982 19156 4988 19168
rect 4264 19128 4988 19156
rect 4982 19116 4988 19128
rect 5040 19116 5046 19168
rect 11624 19156 11652 19255
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 19061 19295 19119 19301
rect 19061 19261 19073 19295
rect 19107 19292 19119 19295
rect 19628 19292 19656 19323
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 21174 19360 21180 19372
rect 21008 19332 21180 19360
rect 21008 19301 21036 19332
rect 21174 19320 21180 19332
rect 21232 19360 21238 19372
rect 21821 19363 21879 19369
rect 21821 19360 21833 19363
rect 21232 19332 21833 19360
rect 21232 19320 21238 19332
rect 21821 19329 21833 19332
rect 21867 19360 21879 19363
rect 23216 19360 23244 19400
rect 25222 19388 25228 19400
rect 25280 19388 25286 19440
rect 33502 19428 33508 19440
rect 32232 19400 33508 19428
rect 32232 19372 32260 19400
rect 33502 19388 33508 19400
rect 33560 19388 33566 19440
rect 39298 19388 39304 19440
rect 39356 19428 39362 19440
rect 43622 19428 43628 19440
rect 39356 19400 41414 19428
rect 43583 19400 43628 19428
rect 39356 19388 39362 19400
rect 23382 19360 23388 19372
rect 21867 19332 23244 19360
rect 23343 19332 23388 19360
rect 21867 19329 21879 19332
rect 21821 19323 21879 19329
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 24394 19360 24400 19372
rect 24355 19332 24400 19360
rect 24394 19320 24400 19332
rect 24452 19320 24458 19372
rect 24670 19369 24676 19372
rect 24664 19323 24676 19369
rect 24728 19360 24734 19372
rect 31389 19363 31447 19369
rect 24728 19332 24764 19360
rect 24670 19320 24676 19323
rect 24728 19320 24734 19332
rect 31389 19329 31401 19363
rect 31435 19360 31447 19363
rect 32030 19360 32036 19372
rect 31435 19332 32036 19360
rect 31435 19329 31447 19332
rect 31389 19323 31447 19329
rect 32030 19320 32036 19332
rect 32088 19320 32094 19372
rect 32214 19360 32220 19372
rect 32127 19332 32220 19360
rect 32214 19320 32220 19332
rect 32272 19320 32278 19372
rect 32490 19369 32496 19372
rect 32484 19360 32496 19369
rect 32451 19332 32496 19360
rect 32484 19323 32496 19332
rect 32490 19320 32496 19323
rect 32548 19320 32554 19372
rect 38838 19320 38844 19372
rect 38896 19360 38902 19372
rect 39666 19360 39672 19372
rect 38896 19332 39672 19360
rect 38896 19320 38902 19332
rect 39666 19320 39672 19332
rect 39724 19320 39730 19372
rect 40126 19360 40132 19372
rect 40039 19332 40132 19360
rect 19107 19264 19656 19292
rect 20993 19295 21051 19301
rect 19107 19261 19119 19264
rect 19061 19255 19119 19261
rect 20993 19261 21005 19295
rect 21039 19261 21051 19295
rect 20993 19255 21051 19261
rect 21082 19252 21088 19304
rect 21140 19292 21146 19304
rect 21140 19264 21185 19292
rect 21140 19252 21146 19264
rect 23014 19252 23020 19304
rect 23072 19292 23078 19304
rect 23109 19295 23167 19301
rect 23109 19292 23121 19295
rect 23072 19264 23121 19292
rect 23072 19252 23078 19264
rect 23109 19261 23121 19264
rect 23155 19261 23167 19295
rect 23109 19255 23167 19261
rect 39206 19252 39212 19304
rect 39264 19292 39270 19304
rect 39758 19292 39764 19304
rect 39264 19264 39764 19292
rect 39264 19252 39270 19264
rect 39758 19252 39764 19264
rect 39816 19252 39822 19304
rect 40052 19301 40080 19332
rect 40126 19320 40132 19332
rect 40184 19360 40190 19372
rect 40497 19363 40555 19369
rect 40497 19360 40509 19363
rect 40184 19332 40509 19360
rect 40184 19320 40190 19332
rect 40497 19329 40509 19332
rect 40543 19329 40555 19363
rect 40678 19360 40684 19372
rect 40639 19332 40684 19360
rect 40497 19323 40555 19329
rect 40678 19320 40684 19332
rect 40736 19320 40742 19372
rect 41386 19360 41414 19400
rect 43622 19388 43628 19400
rect 43680 19388 43686 19440
rect 44266 19388 44272 19440
rect 44324 19388 44330 19440
rect 43346 19360 43352 19372
rect 41386 19332 43352 19360
rect 43346 19320 43352 19332
rect 43404 19320 43410 19372
rect 40037 19295 40095 19301
rect 40037 19261 40049 19295
rect 40083 19261 40095 19295
rect 40037 19255 40095 19261
rect 20806 19224 20812 19236
rect 15396 19196 20812 19224
rect 15396 19156 15424 19196
rect 20806 19184 20812 19196
rect 20864 19184 20870 19236
rect 20898 19184 20904 19236
rect 20956 19224 20962 19236
rect 22649 19227 22707 19233
rect 22649 19224 22661 19227
rect 20956 19196 22661 19224
rect 20956 19184 20962 19196
rect 22649 19193 22661 19196
rect 22695 19224 22707 19227
rect 24302 19224 24308 19236
rect 22695 19196 24308 19224
rect 22695 19193 22707 19196
rect 22649 19187 22707 19193
rect 24302 19184 24308 19196
rect 24360 19184 24366 19236
rect 18874 19156 18880 19168
rect 11624 19128 15424 19156
rect 18835 19128 18880 19156
rect 18874 19116 18880 19128
rect 18932 19116 18938 19168
rect 18969 19159 19027 19165
rect 18969 19125 18981 19159
rect 19015 19156 19027 19159
rect 19426 19156 19432 19168
rect 19015 19128 19432 19156
rect 19015 19125 19027 19128
rect 18969 19119 19027 19125
rect 19426 19116 19432 19128
rect 19484 19116 19490 19168
rect 20073 19159 20131 19165
rect 20073 19125 20085 19159
rect 20119 19156 20131 19159
rect 20346 19156 20352 19168
rect 20119 19128 20352 19156
rect 20119 19125 20131 19128
rect 20073 19119 20131 19125
rect 20346 19116 20352 19128
rect 20404 19116 20410 19168
rect 20530 19156 20536 19168
rect 20491 19128 20536 19156
rect 20530 19116 20536 19128
rect 20588 19116 20594 19168
rect 25774 19156 25780 19168
rect 25735 19128 25780 19156
rect 25774 19116 25780 19128
rect 25832 19116 25838 19168
rect 26234 19156 26240 19168
rect 26195 19128 26240 19156
rect 26234 19116 26240 19128
rect 26292 19116 26298 19168
rect 34793 19159 34851 19165
rect 34793 19125 34805 19159
rect 34839 19156 34851 19159
rect 35434 19156 35440 19168
rect 34839 19128 35440 19156
rect 34839 19125 34851 19128
rect 34793 19119 34851 19125
rect 35434 19116 35440 19128
rect 35492 19156 35498 19168
rect 36446 19156 36452 19168
rect 35492 19128 36452 19156
rect 35492 19116 35498 19128
rect 36446 19116 36452 19128
rect 36504 19116 36510 19168
rect 1104 19066 68816 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 65654 19066
rect 65706 19014 65718 19066
rect 65770 19014 65782 19066
rect 65834 19014 65846 19066
rect 65898 19014 65910 19066
rect 65962 19014 68816 19066
rect 1104 18992 68816 19014
rect 4982 18952 4988 18964
rect 4943 18924 4988 18952
rect 4982 18912 4988 18924
rect 5040 18912 5046 18964
rect 5534 18912 5540 18964
rect 5592 18952 5598 18964
rect 17865 18955 17923 18961
rect 5592 18924 17264 18952
rect 5592 18912 5598 18924
rect 10597 18887 10655 18893
rect 10597 18884 10609 18887
rect 5644 18856 10609 18884
rect 5644 18825 5672 18856
rect 10597 18853 10609 18856
rect 10643 18884 10655 18887
rect 11146 18884 11152 18896
rect 10643 18856 11152 18884
rect 10643 18853 10655 18856
rect 10597 18847 10655 18853
rect 11146 18844 11152 18856
rect 11204 18844 11210 18896
rect 12621 18887 12679 18893
rect 12621 18853 12633 18887
rect 12667 18884 12679 18887
rect 12894 18884 12900 18896
rect 12667 18856 12900 18884
rect 12667 18853 12679 18856
rect 12621 18847 12679 18853
rect 12894 18844 12900 18856
rect 12952 18844 12958 18896
rect 17236 18884 17264 18924
rect 17865 18921 17877 18955
rect 17911 18952 17923 18955
rect 18874 18952 18880 18964
rect 17911 18924 18880 18952
rect 17911 18921 17923 18924
rect 17865 18915 17923 18921
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 19242 18912 19248 18964
rect 19300 18952 19306 18964
rect 19337 18955 19395 18961
rect 19337 18952 19349 18955
rect 19300 18924 19349 18952
rect 19300 18912 19306 18924
rect 19337 18921 19349 18924
rect 19383 18921 19395 18955
rect 23569 18955 23627 18961
rect 23569 18952 23581 18955
rect 19337 18915 19395 18921
rect 19444 18924 23581 18952
rect 19444 18884 19472 18924
rect 23569 18921 23581 18924
rect 23615 18921 23627 18955
rect 24670 18952 24676 18964
rect 24631 18924 24676 18952
rect 23569 18915 23627 18921
rect 17236 18856 19472 18884
rect 23584 18884 23612 18915
rect 24670 18912 24676 18924
rect 24728 18912 24734 18964
rect 27798 18952 27804 18964
rect 25240 18924 27804 18952
rect 25240 18884 25268 18924
rect 27798 18912 27804 18924
rect 27856 18912 27862 18964
rect 28629 18955 28687 18961
rect 28629 18952 28641 18955
rect 27908 18924 28641 18952
rect 23584 18856 25268 18884
rect 25317 18887 25375 18893
rect 25317 18853 25329 18887
rect 25363 18853 25375 18887
rect 25317 18847 25375 18853
rect 5629 18819 5687 18825
rect 5629 18785 5641 18819
rect 5675 18785 5687 18819
rect 5629 18779 5687 18785
rect 7009 18819 7067 18825
rect 7009 18785 7021 18819
rect 7055 18816 7067 18819
rect 7098 18816 7104 18828
rect 7055 18788 7104 18816
rect 7055 18785 7067 18788
rect 7009 18779 7067 18785
rect 7098 18776 7104 18788
rect 7156 18816 7162 18828
rect 7156 18788 18644 18816
rect 7156 18776 7162 18788
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18748 5411 18751
rect 5718 18748 5724 18760
rect 5399 18720 5724 18748
rect 5399 18717 5411 18720
rect 5353 18711 5411 18717
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 11790 18748 11796 18760
rect 11751 18720 11796 18748
rect 11790 18708 11796 18720
rect 11848 18708 11854 18760
rect 16942 18748 16948 18760
rect 16903 18720 16948 18748
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17773 18751 17831 18757
rect 17773 18717 17785 18751
rect 17819 18717 17831 18751
rect 17773 18711 17831 18717
rect 10781 18683 10839 18689
rect 10781 18649 10793 18683
rect 10827 18680 10839 18683
rect 10962 18680 10968 18692
rect 10827 18652 10968 18680
rect 10827 18649 10839 18652
rect 10781 18643 10839 18649
rect 10962 18640 10968 18652
rect 11020 18640 11026 18692
rect 12253 18683 12311 18689
rect 12253 18649 12265 18683
rect 12299 18680 12311 18683
rect 12299 18652 13308 18680
rect 12299 18649 12311 18652
rect 12253 18643 12311 18649
rect 5445 18615 5503 18621
rect 5445 18581 5457 18615
rect 5491 18612 5503 18615
rect 6178 18612 6184 18624
rect 5491 18584 6184 18612
rect 5491 18581 5503 18584
rect 5445 18575 5503 18581
rect 6178 18572 6184 18584
rect 6236 18612 6242 18624
rect 6273 18615 6331 18621
rect 6273 18612 6285 18615
rect 6236 18584 6285 18612
rect 6236 18572 6242 18584
rect 6273 18581 6285 18584
rect 6319 18612 6331 18615
rect 6454 18612 6460 18624
rect 6319 18584 6460 18612
rect 6319 18581 6331 18584
rect 6273 18575 6331 18581
rect 6454 18572 6460 18584
rect 6512 18572 6518 18624
rect 7742 18612 7748 18624
rect 7703 18584 7748 18612
rect 7742 18572 7748 18584
rect 7800 18612 7806 18624
rect 10318 18612 10324 18624
rect 7800 18584 10324 18612
rect 7800 18572 7806 18584
rect 10318 18572 10324 18584
rect 10376 18572 10382 18624
rect 11606 18612 11612 18624
rect 11567 18584 11612 18612
rect 11606 18572 11612 18584
rect 11664 18572 11670 18624
rect 12710 18612 12716 18624
rect 12671 18584 12716 18612
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 13280 18621 13308 18652
rect 16390 18640 16396 18692
rect 16448 18680 16454 18692
rect 17788 18680 17816 18711
rect 16448 18652 17816 18680
rect 18616 18680 18644 18788
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19521 18819 19579 18825
rect 19521 18816 19533 18819
rect 19392 18788 19533 18816
rect 19392 18776 19398 18788
rect 19521 18785 19533 18788
rect 19567 18785 19579 18819
rect 19521 18779 19579 18785
rect 18690 18708 18696 18760
rect 18748 18748 18754 18760
rect 19150 18748 19156 18760
rect 18748 18720 19156 18748
rect 18748 18708 18754 18720
rect 19150 18708 19156 18720
rect 19208 18748 19214 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 19208 18720 19257 18748
rect 19208 18708 19214 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 20530 18748 20536 18760
rect 20491 18720 20536 18748
rect 19245 18711 19303 18717
rect 20530 18708 20536 18720
rect 20588 18708 20594 18760
rect 21177 18751 21235 18757
rect 21177 18717 21189 18751
rect 21223 18748 21235 18751
rect 21266 18748 21272 18760
rect 21223 18720 21272 18748
rect 21223 18717 21235 18720
rect 21177 18711 21235 18717
rect 21266 18708 21272 18720
rect 21324 18708 21330 18760
rect 24857 18751 24915 18757
rect 24857 18717 24869 18751
rect 24903 18748 24915 18751
rect 25332 18748 25360 18847
rect 26418 18844 26424 18896
rect 26476 18884 26482 18896
rect 26973 18887 27031 18893
rect 26973 18884 26985 18887
rect 26476 18856 26985 18884
rect 26476 18844 26482 18856
rect 26973 18853 26985 18856
rect 27019 18884 27031 18887
rect 27246 18884 27252 18896
rect 27019 18856 27252 18884
rect 27019 18853 27031 18856
rect 26973 18847 27031 18853
rect 27246 18844 27252 18856
rect 27304 18844 27310 18896
rect 25774 18816 25780 18828
rect 25735 18788 25780 18816
rect 25774 18776 25780 18788
rect 25832 18776 25838 18828
rect 25961 18819 26019 18825
rect 25961 18785 25973 18819
rect 26007 18816 26019 18819
rect 27062 18816 27068 18828
rect 26007 18788 27068 18816
rect 26007 18785 26019 18788
rect 25961 18779 26019 18785
rect 27062 18776 27068 18788
rect 27120 18776 27126 18828
rect 27801 18819 27859 18825
rect 27801 18816 27813 18819
rect 27172 18788 27813 18816
rect 24903 18720 25360 18748
rect 24903 18717 24915 18720
rect 24857 18711 24915 18717
rect 25406 18708 25412 18760
rect 25464 18748 25470 18760
rect 27172 18748 27200 18788
rect 27801 18785 27813 18788
rect 27847 18816 27859 18819
rect 27908 18816 27936 18924
rect 28629 18921 28641 18924
rect 28675 18921 28687 18955
rect 28629 18915 28687 18921
rect 28997 18955 29055 18961
rect 28997 18921 29009 18955
rect 29043 18952 29055 18955
rect 29362 18952 29368 18964
rect 29043 18924 29368 18952
rect 29043 18921 29055 18924
rect 28997 18915 29055 18921
rect 29362 18912 29368 18924
rect 29420 18912 29426 18964
rect 29638 18912 29644 18964
rect 29696 18952 29702 18964
rect 32582 18952 32588 18964
rect 29696 18924 32588 18952
rect 29696 18912 29702 18924
rect 32582 18912 32588 18924
rect 32640 18952 32646 18964
rect 32861 18955 32919 18961
rect 32861 18952 32873 18955
rect 32640 18924 32873 18952
rect 32640 18912 32646 18924
rect 32861 18921 32873 18924
rect 32907 18921 32919 18955
rect 33318 18952 33324 18964
rect 33279 18924 33324 18952
rect 32861 18915 32919 18921
rect 33318 18912 33324 18924
rect 33376 18912 33382 18964
rect 40221 18955 40279 18961
rect 40221 18921 40233 18955
rect 40267 18952 40279 18955
rect 40586 18952 40592 18964
rect 40267 18924 40592 18952
rect 40267 18921 40279 18924
rect 40221 18915 40279 18921
rect 40586 18912 40592 18924
rect 40644 18912 40650 18964
rect 44266 18952 44272 18964
rect 44227 18924 44272 18952
rect 44266 18912 44272 18924
rect 44324 18912 44330 18964
rect 45002 18912 45008 18964
rect 45060 18952 45066 18964
rect 45097 18955 45155 18961
rect 45097 18952 45109 18955
rect 45060 18924 45109 18952
rect 45060 18912 45066 18924
rect 45097 18921 45109 18924
rect 45143 18921 45155 18955
rect 45097 18915 45155 18921
rect 28077 18887 28135 18893
rect 28077 18853 28089 18887
rect 28123 18884 28135 18887
rect 30098 18884 30104 18896
rect 28123 18856 30104 18884
rect 28123 18853 28135 18856
rect 28077 18847 28135 18853
rect 30098 18844 30104 18856
rect 30156 18844 30162 18896
rect 27847 18788 27936 18816
rect 27847 18785 27859 18788
rect 27801 18779 27859 18785
rect 33594 18776 33600 18828
rect 33652 18816 33658 18828
rect 33781 18819 33839 18825
rect 33781 18816 33793 18819
rect 33652 18788 33793 18816
rect 33652 18776 33658 18788
rect 33781 18785 33793 18788
rect 33827 18785 33839 18819
rect 33781 18779 33839 18785
rect 33870 18776 33876 18828
rect 33928 18816 33934 18828
rect 39298 18816 39304 18828
rect 33928 18788 33973 18816
rect 39259 18788 39304 18816
rect 33928 18776 33934 18788
rect 39298 18776 39304 18788
rect 39356 18776 39362 18828
rect 25464 18720 27200 18748
rect 25464 18708 25470 18720
rect 27246 18708 27252 18760
rect 27304 18748 27310 18760
rect 27709 18751 27767 18757
rect 27709 18748 27721 18751
rect 27304 18720 27721 18748
rect 27304 18708 27310 18720
rect 27709 18717 27721 18720
rect 27755 18717 27767 18751
rect 27709 18711 27767 18717
rect 28537 18751 28595 18757
rect 28537 18717 28549 18751
rect 28583 18717 28595 18751
rect 28537 18711 28595 18717
rect 31481 18751 31539 18757
rect 31481 18717 31493 18751
rect 31527 18748 31539 18751
rect 32214 18748 32220 18760
rect 31527 18720 32220 18748
rect 31527 18717 31539 18720
rect 31481 18711 31539 18717
rect 19334 18680 19340 18692
rect 18616 18652 19340 18680
rect 16448 18640 16454 18652
rect 19334 18640 19340 18652
rect 19392 18640 19398 18692
rect 21422 18683 21480 18689
rect 21422 18680 21434 18683
rect 20732 18652 21434 18680
rect 13265 18615 13323 18621
rect 13265 18581 13277 18615
rect 13311 18612 13323 18615
rect 13538 18612 13544 18624
rect 13311 18584 13544 18612
rect 13311 18581 13323 18584
rect 13265 18575 13323 18581
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 17126 18612 17132 18624
rect 17087 18584 17132 18612
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 19797 18615 19855 18621
rect 19797 18581 19809 18615
rect 19843 18612 19855 18615
rect 19978 18612 19984 18624
rect 19843 18584 19984 18612
rect 19843 18581 19855 18584
rect 19797 18575 19855 18581
rect 19978 18572 19984 18584
rect 20036 18572 20042 18624
rect 20732 18621 20760 18652
rect 21422 18649 21434 18652
rect 21468 18649 21480 18683
rect 23014 18680 23020 18692
rect 21422 18643 21480 18649
rect 22572 18652 23020 18680
rect 22572 18621 22600 18652
rect 23014 18640 23020 18652
rect 23072 18680 23078 18692
rect 23293 18683 23351 18689
rect 23293 18680 23305 18683
rect 23072 18652 23305 18680
rect 23072 18640 23078 18652
rect 23293 18649 23305 18652
rect 23339 18649 23351 18683
rect 23293 18643 23351 18649
rect 26234 18640 26240 18692
rect 26292 18680 26298 18692
rect 28552 18680 28580 18711
rect 32214 18708 32220 18720
rect 32272 18708 32278 18760
rect 40126 18748 40132 18760
rect 40087 18720 40132 18748
rect 40126 18708 40132 18720
rect 40184 18708 40190 18760
rect 40313 18751 40371 18757
rect 40313 18717 40325 18751
rect 40359 18748 40371 18751
rect 40678 18748 40684 18760
rect 40359 18720 40684 18748
rect 40359 18717 40371 18720
rect 40313 18711 40371 18717
rect 29178 18680 29184 18692
rect 26292 18652 29184 18680
rect 26292 18640 26298 18652
rect 29178 18640 29184 18652
rect 29236 18680 29242 18692
rect 29549 18683 29607 18689
rect 29549 18680 29561 18683
rect 29236 18652 29561 18680
rect 29236 18640 29242 18652
rect 29549 18649 29561 18652
rect 29595 18680 29607 18683
rect 31110 18680 31116 18692
rect 29595 18652 31116 18680
rect 29595 18649 29607 18652
rect 29549 18643 29607 18649
rect 31110 18640 31116 18652
rect 31168 18640 31174 18692
rect 31754 18689 31760 18692
rect 31748 18643 31760 18689
rect 31812 18680 31818 18692
rect 31812 18652 31848 18680
rect 31754 18640 31760 18643
rect 31812 18640 31818 18652
rect 32490 18640 32496 18692
rect 32548 18680 32554 18692
rect 33689 18683 33747 18689
rect 33689 18680 33701 18683
rect 32548 18652 33701 18680
rect 32548 18640 32554 18652
rect 33689 18649 33701 18652
rect 33735 18680 33747 18683
rect 38010 18680 38016 18692
rect 33735 18652 38016 18680
rect 33735 18649 33747 18652
rect 33689 18643 33747 18649
rect 38010 18640 38016 18652
rect 38068 18640 38074 18692
rect 38838 18640 38844 18692
rect 38896 18680 38902 18692
rect 39034 18683 39092 18689
rect 39034 18680 39046 18683
rect 38896 18652 39046 18680
rect 38896 18640 38902 18652
rect 39034 18649 39046 18652
rect 39080 18649 39092 18683
rect 39034 18643 39092 18649
rect 20717 18615 20775 18621
rect 20717 18581 20729 18615
rect 20763 18581 20775 18615
rect 20717 18575 20775 18581
rect 22557 18615 22615 18621
rect 22557 18581 22569 18615
rect 22603 18581 22615 18615
rect 25682 18612 25688 18624
rect 25643 18584 25688 18612
rect 22557 18575 22615 18581
rect 25682 18572 25688 18584
rect 25740 18572 25746 18624
rect 30190 18572 30196 18624
rect 30248 18612 30254 18624
rect 34514 18612 34520 18624
rect 30248 18584 34520 18612
rect 30248 18572 30254 18584
rect 34514 18572 34520 18584
rect 34572 18572 34578 18624
rect 37918 18612 37924 18624
rect 37831 18584 37924 18612
rect 37918 18572 37924 18584
rect 37976 18612 37982 18624
rect 40328 18612 40356 18711
rect 40678 18708 40684 18720
rect 40736 18708 40742 18760
rect 41874 18708 41880 18760
rect 41932 18748 41938 18760
rect 44177 18751 44235 18757
rect 44177 18748 44189 18751
rect 41932 18720 44189 18748
rect 41932 18708 41938 18720
rect 44177 18717 44189 18720
rect 44223 18748 44235 18751
rect 45005 18751 45063 18757
rect 45005 18748 45017 18751
rect 44223 18720 45017 18748
rect 44223 18717 44235 18720
rect 44177 18711 44235 18717
rect 45005 18717 45017 18720
rect 45051 18717 45063 18751
rect 67818 18748 67824 18760
rect 67779 18720 67824 18748
rect 45005 18711 45063 18717
rect 67818 18708 67824 18720
rect 67876 18708 67882 18760
rect 37976 18584 40356 18612
rect 37976 18572 37982 18584
rect 55122 18572 55128 18624
rect 55180 18612 55186 18624
rect 55766 18612 55772 18624
rect 55180 18584 55772 18612
rect 55180 18572 55186 18584
rect 55766 18572 55772 18584
rect 55824 18572 55830 18624
rect 68002 18612 68008 18624
rect 67963 18584 68008 18612
rect 68002 18572 68008 18584
rect 68060 18572 68066 18624
rect 1104 18522 68816 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 68816 18522
rect 1104 18448 68816 18470
rect 7193 18411 7251 18417
rect 7193 18377 7205 18411
rect 7239 18408 7251 18411
rect 7374 18408 7380 18420
rect 7239 18380 7380 18408
rect 7239 18377 7251 18380
rect 7193 18371 7251 18377
rect 7374 18368 7380 18380
rect 7432 18368 7438 18420
rect 8478 18408 8484 18420
rect 8439 18380 8484 18408
rect 8478 18368 8484 18380
rect 8536 18368 8542 18420
rect 15378 18368 15384 18420
rect 15436 18408 15442 18420
rect 15749 18411 15807 18417
rect 15749 18408 15761 18411
rect 15436 18380 15761 18408
rect 15436 18368 15442 18380
rect 15749 18377 15761 18380
rect 15795 18377 15807 18411
rect 15749 18371 15807 18377
rect 18417 18411 18475 18417
rect 18417 18377 18429 18411
rect 18463 18408 18475 18411
rect 18966 18408 18972 18420
rect 18463 18380 18972 18408
rect 18463 18377 18475 18380
rect 18417 18371 18475 18377
rect 18966 18368 18972 18380
rect 19024 18368 19030 18420
rect 19242 18408 19248 18420
rect 19203 18380 19248 18408
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19889 18411 19947 18417
rect 19889 18408 19901 18411
rect 19392 18380 19901 18408
rect 19392 18368 19398 18380
rect 19889 18377 19901 18380
rect 19935 18408 19947 18411
rect 19935 18380 20484 18408
rect 19935 18377 19947 18380
rect 19889 18371 19947 18377
rect 5442 18300 5448 18352
rect 5500 18340 5506 18352
rect 5500 18312 8340 18340
rect 5500 18300 5506 18312
rect 7653 18275 7711 18281
rect 7653 18241 7665 18275
rect 7699 18272 7711 18275
rect 7742 18272 7748 18284
rect 7699 18244 7748 18272
rect 7699 18241 7711 18244
rect 7653 18235 7711 18241
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 8312 18281 8340 18312
rect 11606 18300 11612 18352
rect 11664 18340 11670 18352
rect 11762 18343 11820 18349
rect 11762 18340 11774 18343
rect 11664 18312 11774 18340
rect 11664 18300 11670 18312
rect 11762 18309 11774 18312
rect 11808 18309 11820 18343
rect 11762 18303 11820 18309
rect 8297 18275 8355 18281
rect 8297 18241 8309 18275
rect 8343 18241 8355 18275
rect 11514 18272 11520 18284
rect 11475 18244 11520 18272
rect 8297 18235 8355 18241
rect 11514 18232 11520 18244
rect 11572 18232 11578 18284
rect 15657 18275 15715 18281
rect 15657 18241 15669 18275
rect 15703 18272 15715 18275
rect 16390 18272 16396 18284
rect 15703 18244 16396 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 16390 18232 16396 18244
rect 16448 18232 16454 18284
rect 17126 18232 17132 18284
rect 17184 18272 17190 18284
rect 17293 18275 17351 18281
rect 17293 18272 17305 18275
rect 17184 18244 17305 18272
rect 17184 18232 17190 18244
rect 17293 18241 17305 18244
rect 17339 18241 17351 18275
rect 17293 18235 17351 18241
rect 18874 18232 18880 18284
rect 18932 18272 18938 18284
rect 19061 18275 19119 18281
rect 19061 18272 19073 18275
rect 18932 18244 19073 18272
rect 18932 18232 18938 18244
rect 19061 18241 19073 18244
rect 19107 18241 19119 18275
rect 19061 18235 19119 18241
rect 19150 18232 19156 18284
rect 19208 18272 19214 18284
rect 20456 18281 20484 18380
rect 20714 18368 20720 18420
rect 20772 18408 20778 18420
rect 20772 18380 22094 18408
rect 20772 18368 20778 18380
rect 22066 18340 22094 18380
rect 22738 18368 22744 18420
rect 22796 18408 22802 18420
rect 22833 18411 22891 18417
rect 22833 18408 22845 18411
rect 22796 18380 22845 18408
rect 22796 18368 22802 18380
rect 22833 18377 22845 18380
rect 22879 18408 22891 18411
rect 23658 18408 23664 18420
rect 22879 18380 23664 18408
rect 22879 18377 22891 18380
rect 22833 18371 22891 18377
rect 23658 18368 23664 18380
rect 23716 18368 23722 18420
rect 25317 18411 25375 18417
rect 25317 18377 25329 18411
rect 25363 18408 25375 18411
rect 26326 18408 26332 18420
rect 25363 18380 26332 18408
rect 25363 18377 25375 18380
rect 25317 18371 25375 18377
rect 26326 18368 26332 18380
rect 26384 18368 26390 18420
rect 29178 18408 29184 18420
rect 29139 18380 29184 18408
rect 29178 18368 29184 18380
rect 29236 18368 29242 18420
rect 32030 18368 32036 18420
rect 32088 18408 32094 18420
rect 32125 18411 32183 18417
rect 32125 18408 32137 18411
rect 32088 18380 32137 18408
rect 32088 18368 32094 18380
rect 32125 18377 32137 18380
rect 32171 18377 32183 18411
rect 32582 18408 32588 18420
rect 32543 18380 32588 18408
rect 32125 18371 32183 18377
rect 32582 18368 32588 18380
rect 32640 18368 32646 18420
rect 33689 18411 33747 18417
rect 33689 18377 33701 18411
rect 33735 18408 33747 18411
rect 33870 18408 33876 18420
rect 33735 18380 33876 18408
rect 33735 18377 33747 18380
rect 33689 18371 33747 18377
rect 33870 18368 33876 18380
rect 33928 18368 33934 18420
rect 37918 18408 37924 18420
rect 37879 18380 37924 18408
rect 37918 18368 37924 18380
rect 37976 18368 37982 18420
rect 38010 18368 38016 18420
rect 38068 18408 38074 18420
rect 38381 18411 38439 18417
rect 38068 18380 38113 18408
rect 38068 18368 38074 18380
rect 38381 18377 38393 18411
rect 38427 18377 38439 18411
rect 38838 18408 38844 18420
rect 38799 18380 38844 18408
rect 38381 18371 38439 18377
rect 22066 18312 38148 18340
rect 19337 18275 19395 18281
rect 19337 18272 19349 18275
rect 19208 18244 19349 18272
rect 19208 18232 19214 18244
rect 19337 18241 19349 18244
rect 19383 18241 19395 18275
rect 19337 18235 19395 18241
rect 20441 18275 20499 18281
rect 20441 18241 20453 18275
rect 20487 18272 20499 18275
rect 23382 18272 23388 18284
rect 20487 18244 23388 18272
rect 20487 18241 20499 18244
rect 20441 18235 20499 18241
rect 23382 18232 23388 18244
rect 23440 18232 23446 18284
rect 23937 18275 23995 18281
rect 23937 18241 23949 18275
rect 23983 18272 23995 18275
rect 24946 18272 24952 18284
rect 23983 18244 24952 18272
rect 23983 18241 23995 18244
rect 23937 18235 23995 18241
rect 24946 18232 24952 18244
rect 25004 18232 25010 18284
rect 26234 18272 26240 18284
rect 25148 18244 26240 18272
rect 8110 18204 8116 18216
rect 8071 18176 8116 18204
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 12894 18164 12900 18216
rect 12952 18204 12958 18216
rect 13817 18207 13875 18213
rect 13817 18204 13829 18207
rect 12952 18176 13829 18204
rect 12952 18164 12958 18176
rect 13817 18173 13829 18176
rect 13863 18173 13875 18207
rect 15930 18204 15936 18216
rect 15891 18176 15936 18204
rect 13817 18167 13875 18173
rect 15930 18164 15936 18176
rect 15988 18164 15994 18216
rect 17037 18207 17095 18213
rect 17037 18173 17049 18207
rect 17083 18173 17095 18207
rect 17037 18167 17095 18173
rect 12526 18096 12532 18148
rect 12584 18136 12590 18148
rect 13357 18139 13415 18145
rect 13357 18136 13369 18139
rect 12584 18108 13369 18136
rect 12584 18096 12590 18108
rect 13357 18105 13369 18108
rect 13403 18105 13415 18139
rect 13357 18099 13415 18105
rect 13538 18096 13544 18148
rect 13596 18136 13602 18148
rect 14369 18139 14427 18145
rect 14369 18136 14381 18139
rect 13596 18108 14381 18136
rect 13596 18096 13602 18108
rect 14369 18105 14381 18108
rect 14415 18136 14427 18139
rect 14415 18108 15516 18136
rect 14415 18105 14427 18108
rect 14369 18099 14427 18105
rect 7466 18068 7472 18080
rect 7427 18040 7472 18068
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 12894 18068 12900 18080
rect 12855 18040 12900 18068
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 15289 18071 15347 18077
rect 15289 18037 15301 18071
rect 15335 18068 15347 18071
rect 15378 18068 15384 18080
rect 15335 18040 15384 18068
rect 15335 18037 15347 18040
rect 15289 18031 15347 18037
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 15488 18068 15516 18108
rect 15746 18096 15752 18148
rect 15804 18136 15810 18148
rect 17052 18136 17080 18167
rect 20806 18164 20812 18216
rect 20864 18204 20870 18216
rect 25038 18204 25044 18216
rect 20864 18176 24900 18204
rect 24999 18176 25044 18204
rect 20864 18164 20870 18176
rect 20898 18136 20904 18148
rect 15804 18108 17080 18136
rect 17972 18108 20904 18136
rect 15804 18096 15810 18108
rect 17972 18068 18000 18108
rect 20898 18096 20904 18108
rect 20956 18096 20962 18148
rect 22281 18139 22339 18145
rect 22281 18105 22293 18139
rect 22327 18136 22339 18139
rect 23106 18136 23112 18148
rect 22327 18108 23112 18136
rect 22327 18105 22339 18108
rect 22281 18099 22339 18105
rect 23106 18096 23112 18108
rect 23164 18096 23170 18148
rect 23474 18096 23480 18148
rect 23532 18136 23538 18148
rect 24397 18139 24455 18145
rect 24397 18136 24409 18139
rect 23532 18108 24409 18136
rect 23532 18096 23538 18108
rect 24397 18105 24409 18108
rect 24443 18105 24455 18139
rect 24872 18136 24900 18176
rect 25038 18164 25044 18176
rect 25096 18164 25102 18216
rect 25148 18136 25176 18244
rect 26234 18232 26240 18244
rect 26292 18232 26298 18284
rect 27154 18232 27160 18284
rect 27212 18272 27218 18284
rect 29365 18275 29423 18281
rect 29365 18272 29377 18275
rect 27212 18244 29377 18272
rect 27212 18232 27218 18244
rect 29365 18241 29377 18244
rect 29411 18272 29423 18275
rect 30745 18275 30803 18281
rect 30745 18272 30757 18275
rect 29411 18244 30757 18272
rect 29411 18241 29423 18244
rect 29365 18235 29423 18241
rect 30745 18241 30757 18244
rect 30791 18241 30803 18275
rect 30745 18235 30803 18241
rect 31205 18275 31263 18281
rect 31205 18241 31217 18275
rect 31251 18272 31263 18275
rect 31662 18272 31668 18284
rect 31251 18244 31668 18272
rect 31251 18241 31263 18244
rect 31205 18235 31263 18241
rect 31662 18232 31668 18244
rect 31720 18232 31726 18284
rect 32490 18272 32496 18284
rect 32451 18244 32496 18272
rect 32490 18232 32496 18244
rect 32548 18232 32554 18284
rect 33781 18275 33839 18281
rect 33781 18241 33793 18275
rect 33827 18241 33839 18275
rect 34514 18272 34520 18284
rect 34475 18244 34520 18272
rect 33781 18235 33839 18241
rect 26970 18204 26976 18216
rect 24872 18108 25176 18136
rect 25240 18176 26976 18204
rect 24397 18099 24455 18105
rect 15488 18040 18000 18068
rect 18877 18071 18935 18077
rect 18877 18037 18889 18071
rect 18923 18068 18935 18071
rect 18966 18068 18972 18080
rect 18923 18040 18972 18068
rect 18923 18037 18935 18040
rect 18877 18031 18935 18037
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 20671 18071 20729 18077
rect 20671 18037 20683 18071
rect 20717 18068 20729 18071
rect 20990 18068 20996 18080
rect 20717 18040 20996 18068
rect 20717 18037 20729 18040
rect 20671 18031 20729 18037
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 23385 18071 23443 18077
rect 23385 18037 23397 18071
rect 23431 18068 23443 18071
rect 24026 18068 24032 18080
rect 23431 18040 24032 18068
rect 23431 18037 23443 18040
rect 23385 18031 23443 18037
rect 24026 18028 24032 18040
rect 24084 18028 24090 18080
rect 24412 18068 24440 18099
rect 24949 18071 25007 18077
rect 24949 18068 24961 18071
rect 24412 18040 24961 18068
rect 24949 18037 24961 18040
rect 24995 18068 25007 18071
rect 25240 18068 25268 18176
rect 26970 18164 26976 18176
rect 27028 18164 27034 18216
rect 31573 18207 31631 18213
rect 31573 18173 31585 18207
rect 31619 18204 31631 18207
rect 32674 18204 32680 18216
rect 31619 18176 31754 18204
rect 32635 18176 32680 18204
rect 31619 18173 31631 18176
rect 31573 18167 31631 18173
rect 26326 18096 26332 18148
rect 26384 18136 26390 18148
rect 27522 18136 27528 18148
rect 26384 18108 27528 18136
rect 26384 18096 26390 18108
rect 27522 18096 27528 18108
rect 27580 18136 27586 18148
rect 31726 18136 31754 18176
rect 32674 18164 32680 18176
rect 32732 18164 32738 18216
rect 33502 18164 33508 18216
rect 33560 18204 33566 18216
rect 33796 18204 33824 18235
rect 34514 18232 34520 18244
rect 34572 18232 34578 18284
rect 34698 18204 34704 18216
rect 33560 18176 34704 18204
rect 33560 18164 33566 18176
rect 34698 18164 34704 18176
rect 34756 18164 34762 18216
rect 37826 18204 37832 18216
rect 37787 18176 37832 18204
rect 37826 18164 37832 18176
rect 37884 18164 37890 18216
rect 38120 18204 38148 18312
rect 38396 18272 38424 18371
rect 38838 18368 38844 18380
rect 38896 18368 38902 18420
rect 39025 18275 39083 18281
rect 39025 18272 39037 18275
rect 38396 18244 39037 18272
rect 39025 18241 39037 18244
rect 39071 18241 39083 18275
rect 39025 18235 39083 18241
rect 41598 18204 41604 18216
rect 38120 18176 41604 18204
rect 41598 18164 41604 18176
rect 41656 18164 41662 18216
rect 39666 18136 39672 18148
rect 27580 18108 31248 18136
rect 31726 18108 39672 18136
rect 27580 18096 27586 18108
rect 25866 18068 25872 18080
rect 24995 18040 25268 18068
rect 25827 18040 25872 18068
rect 24995 18037 25007 18040
rect 24949 18031 25007 18037
rect 25866 18028 25872 18040
rect 25924 18028 25930 18080
rect 31220 18068 31248 18108
rect 39666 18096 39672 18108
rect 39724 18096 39730 18148
rect 32582 18068 32588 18080
rect 31220 18040 32588 18068
rect 32582 18028 32588 18040
rect 32640 18028 32646 18080
rect 34698 18068 34704 18080
rect 34659 18040 34704 18068
rect 34698 18028 34704 18040
rect 34756 18028 34762 18080
rect 43530 18068 43536 18080
rect 43491 18040 43536 18068
rect 43530 18028 43536 18040
rect 43588 18028 43594 18080
rect 1104 17978 68816 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 65654 17978
rect 65706 17926 65718 17978
rect 65770 17926 65782 17978
rect 65834 17926 65846 17978
rect 65898 17926 65910 17978
rect 65962 17926 68816 17978
rect 1104 17904 68816 17926
rect 11790 17824 11796 17876
rect 11848 17864 11854 17876
rect 11977 17867 12035 17873
rect 11977 17864 11989 17867
rect 11848 17836 11989 17864
rect 11848 17824 11854 17836
rect 11977 17833 11989 17836
rect 12023 17833 12035 17867
rect 16390 17864 16396 17876
rect 16351 17836 16396 17864
rect 11977 17827 12035 17833
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 16942 17824 16948 17876
rect 17000 17864 17006 17876
rect 17037 17867 17095 17873
rect 17037 17864 17049 17867
rect 17000 17836 17049 17864
rect 17000 17824 17006 17836
rect 17037 17833 17049 17836
rect 17083 17833 17095 17867
rect 17037 17827 17095 17833
rect 20438 17824 20444 17876
rect 20496 17864 20502 17876
rect 26145 17867 26203 17873
rect 26145 17864 26157 17867
rect 20496 17836 26157 17864
rect 20496 17824 20502 17836
rect 26145 17833 26157 17836
rect 26191 17864 26203 17867
rect 30282 17864 30288 17876
rect 26191 17836 30288 17864
rect 26191 17833 26203 17836
rect 26145 17827 26203 17833
rect 30282 17824 30288 17836
rect 30340 17864 30346 17876
rect 33502 17864 33508 17876
rect 30340 17836 31156 17864
rect 33463 17836 33508 17864
rect 30340 17824 30346 17836
rect 6454 17756 6460 17808
rect 6512 17796 6518 17808
rect 6512 17768 13492 17796
rect 6512 17756 6518 17768
rect 5442 17728 5448 17740
rect 5403 17700 5448 17728
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 7285 17731 7343 17737
rect 7285 17697 7297 17731
rect 7331 17728 7343 17731
rect 7374 17728 7380 17740
rect 7331 17700 7380 17728
rect 7331 17697 7343 17700
rect 7285 17691 7343 17697
rect 7374 17688 7380 17700
rect 7432 17688 7438 17740
rect 7650 17728 7656 17740
rect 7563 17700 7656 17728
rect 7650 17688 7656 17700
rect 7708 17728 7714 17740
rect 8110 17728 8116 17740
rect 7708 17700 8116 17728
rect 7708 17688 7714 17700
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 10962 17688 10968 17740
rect 11020 17728 11026 17740
rect 12529 17731 12587 17737
rect 12529 17728 12541 17731
rect 11020 17700 12541 17728
rect 11020 17688 11026 17700
rect 12529 17697 12541 17700
rect 12575 17697 12587 17731
rect 12529 17691 12587 17697
rect 5353 17663 5411 17669
rect 5353 17629 5365 17663
rect 5399 17660 5411 17663
rect 5718 17660 5724 17672
rect 5399 17632 5724 17660
rect 5399 17629 5411 17632
rect 5353 17623 5411 17629
rect 5718 17620 5724 17632
rect 5776 17620 5782 17672
rect 7745 17663 7803 17669
rect 7745 17629 7757 17663
rect 7791 17660 7803 17663
rect 7791 17632 8156 17660
rect 7791 17629 7803 17632
rect 7745 17623 7803 17629
rect 8128 17604 8156 17632
rect 10410 17620 10416 17672
rect 10468 17660 10474 17672
rect 11057 17663 11115 17669
rect 11057 17660 11069 17663
rect 10468 17632 11069 17660
rect 10468 17620 10474 17632
rect 11057 17629 11069 17632
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 11333 17663 11391 17669
rect 11333 17629 11345 17663
rect 11379 17629 11391 17663
rect 11333 17623 11391 17629
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17660 12403 17663
rect 12894 17660 12900 17672
rect 12391 17632 12900 17660
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 8110 17552 8116 17604
rect 8168 17552 8174 17604
rect 11348 17592 11376 17623
rect 12894 17620 12900 17632
rect 12952 17620 12958 17672
rect 12526 17592 12532 17604
rect 11348 17564 12532 17592
rect 12526 17552 12532 17564
rect 12584 17552 12590 17604
rect 13464 17601 13492 17768
rect 17402 17756 17408 17808
rect 17460 17796 17466 17808
rect 19889 17799 19947 17805
rect 17460 17768 17632 17796
rect 17460 17756 17466 17768
rect 17604 17737 17632 17768
rect 19889 17765 19901 17799
rect 19935 17796 19947 17799
rect 21082 17796 21088 17808
rect 19935 17768 21088 17796
rect 19935 17765 19947 17768
rect 19889 17759 19947 17765
rect 21082 17756 21088 17768
rect 21140 17756 21146 17808
rect 23014 17796 23020 17808
rect 22975 17768 23020 17796
rect 23014 17756 23020 17768
rect 23072 17756 23078 17808
rect 27246 17756 27252 17808
rect 27304 17796 27310 17808
rect 27341 17799 27399 17805
rect 27341 17796 27353 17799
rect 27304 17768 27353 17796
rect 27304 17756 27310 17768
rect 27341 17765 27353 17768
rect 27387 17765 27399 17799
rect 27341 17759 27399 17765
rect 17589 17731 17647 17737
rect 17589 17697 17601 17731
rect 17635 17728 17647 17731
rect 17635 17700 19748 17728
rect 17635 17697 17647 17700
rect 17589 17691 17647 17697
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17660 15071 17663
rect 15746 17660 15752 17672
rect 15059 17632 15752 17660
rect 15059 17629 15071 17632
rect 15013 17623 15071 17629
rect 15746 17620 15752 17632
rect 15804 17620 15810 17672
rect 17405 17663 17463 17669
rect 17405 17629 17417 17663
rect 17451 17660 17463 17663
rect 17862 17660 17868 17672
rect 17451 17632 17868 17660
rect 17451 17629 17463 17632
rect 17405 17623 17463 17629
rect 17862 17620 17868 17632
rect 17920 17620 17926 17672
rect 19720 17669 19748 17700
rect 20254 17688 20260 17740
rect 20312 17728 20318 17740
rect 25866 17728 25872 17740
rect 20312 17700 25872 17728
rect 20312 17688 20318 17700
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17629 19763 17663
rect 20622 17660 20628 17672
rect 20583 17632 20628 17660
rect 19705 17623 19763 17629
rect 20622 17620 20628 17632
rect 20680 17620 20686 17672
rect 20806 17660 20812 17672
rect 20767 17632 20812 17660
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 21266 17660 21272 17672
rect 21227 17632 21272 17660
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 23658 17660 23664 17672
rect 23619 17632 23664 17660
rect 23658 17620 23664 17632
rect 23716 17620 23722 17672
rect 24872 17669 24900 17700
rect 25866 17688 25872 17700
rect 25924 17688 25930 17740
rect 24857 17663 24915 17669
rect 24857 17629 24869 17663
rect 24903 17629 24915 17663
rect 24857 17623 24915 17629
rect 25130 17620 25136 17672
rect 25188 17660 25194 17672
rect 25682 17660 25688 17672
rect 25188 17632 25688 17660
rect 25188 17620 25194 17632
rect 25682 17620 25688 17632
rect 25740 17660 25746 17672
rect 30101 17663 30159 17669
rect 25740 17632 27476 17660
rect 25740 17620 25746 17632
rect 13265 17595 13323 17601
rect 13265 17561 13277 17595
rect 13311 17561 13323 17595
rect 13265 17555 13323 17561
rect 13449 17595 13507 17601
rect 13449 17561 13461 17595
rect 13495 17592 13507 17595
rect 15102 17592 15108 17604
rect 13495 17564 15108 17592
rect 13495 17561 13507 17564
rect 13449 17555 13507 17561
rect 5721 17527 5779 17533
rect 5721 17493 5733 17527
rect 5767 17524 5779 17527
rect 6914 17524 6920 17536
rect 5767 17496 6920 17524
rect 5767 17493 5779 17496
rect 5721 17487 5779 17493
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 7006 17484 7012 17536
rect 7064 17524 7070 17536
rect 7929 17527 7987 17533
rect 7929 17524 7941 17527
rect 7064 17496 7941 17524
rect 7064 17484 7070 17496
rect 7929 17493 7941 17496
rect 7975 17493 7987 17527
rect 7929 17487 7987 17493
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 11149 17527 11207 17533
rect 11149 17524 11161 17527
rect 10836 17496 11161 17524
rect 10836 17484 10842 17496
rect 11149 17493 11161 17496
rect 11195 17493 11207 17527
rect 11149 17487 11207 17493
rect 11517 17527 11575 17533
rect 11517 17493 11529 17527
rect 11563 17524 11575 17527
rect 11790 17524 11796 17536
rect 11563 17496 11796 17524
rect 11563 17493 11575 17496
rect 11517 17487 11575 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 12342 17484 12348 17536
rect 12400 17524 12406 17536
rect 12437 17527 12495 17533
rect 12437 17524 12449 17527
rect 12400 17496 12449 17524
rect 12400 17484 12406 17496
rect 12437 17493 12449 17496
rect 12483 17493 12495 17527
rect 13280 17524 13308 17555
rect 15102 17552 15108 17564
rect 15160 17552 15166 17604
rect 15286 17601 15292 17604
rect 15280 17555 15292 17601
rect 15344 17592 15350 17604
rect 15344 17564 15380 17592
rect 15286 17552 15292 17555
rect 15344 17552 15350 17564
rect 16482 17552 16488 17604
rect 16540 17592 16546 17604
rect 20717 17595 20775 17601
rect 16540 17564 20668 17592
rect 16540 17552 16546 17564
rect 13354 17524 13360 17536
rect 13267 17496 13360 17524
rect 12437 17487 12495 17493
rect 13354 17484 13360 17496
rect 13412 17524 13418 17536
rect 14182 17524 14188 17536
rect 13412 17496 14188 17524
rect 13412 17484 13418 17496
rect 14182 17484 14188 17496
rect 14240 17484 14246 17536
rect 17310 17484 17316 17536
rect 17368 17524 17374 17536
rect 17497 17527 17555 17533
rect 17497 17524 17509 17527
rect 17368 17496 17509 17524
rect 17368 17484 17374 17496
rect 17497 17493 17509 17496
rect 17543 17524 17555 17527
rect 18233 17527 18291 17533
rect 18233 17524 18245 17527
rect 17543 17496 18245 17524
rect 17543 17493 17555 17496
rect 17497 17487 17555 17493
rect 18233 17493 18245 17496
rect 18279 17524 18291 17527
rect 18598 17524 18604 17536
rect 18279 17496 18604 17524
rect 18279 17493 18291 17496
rect 18233 17487 18291 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 20640 17524 20668 17564
rect 20717 17561 20729 17595
rect 20763 17592 20775 17595
rect 21545 17595 21603 17601
rect 21545 17592 21557 17595
rect 20763 17564 21557 17592
rect 20763 17561 20775 17564
rect 20717 17555 20775 17561
rect 21545 17561 21557 17564
rect 21591 17561 21603 17595
rect 21545 17555 21603 17561
rect 22554 17552 22560 17604
rect 22612 17552 22618 17604
rect 26234 17552 26240 17604
rect 26292 17592 26298 17604
rect 27154 17592 27160 17604
rect 26292 17564 27160 17592
rect 26292 17552 26298 17564
rect 27154 17552 27160 17564
rect 27212 17552 27218 17604
rect 21174 17524 21180 17536
rect 20640 17496 21180 17524
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 23382 17484 23388 17536
rect 23440 17524 23446 17536
rect 23477 17527 23535 17533
rect 23477 17524 23489 17527
rect 23440 17496 23489 17524
rect 23440 17484 23446 17496
rect 23477 17493 23489 17496
rect 23523 17493 23535 17527
rect 27448 17524 27476 17632
rect 30101 17629 30113 17663
rect 30147 17660 30159 17663
rect 31128 17660 31156 17836
rect 33502 17824 33508 17836
rect 33560 17824 33566 17876
rect 36817 17867 36875 17873
rect 36817 17833 36829 17867
rect 36863 17864 36875 17867
rect 37826 17864 37832 17876
rect 36863 17836 37832 17864
rect 36863 17833 36875 17836
rect 36817 17827 36875 17833
rect 37826 17824 37832 17836
rect 37884 17824 37890 17876
rect 31481 17799 31539 17805
rect 31481 17765 31493 17799
rect 31527 17765 31539 17799
rect 31481 17759 31539 17765
rect 31496 17728 31524 17759
rect 31662 17728 31668 17740
rect 31496 17700 31668 17728
rect 31662 17688 31668 17700
rect 31720 17728 31726 17740
rect 32401 17731 32459 17737
rect 32401 17728 32413 17731
rect 31720 17700 32413 17728
rect 31720 17688 31726 17700
rect 32401 17697 32413 17700
rect 32447 17697 32459 17731
rect 32401 17691 32459 17697
rect 32585 17731 32643 17737
rect 32585 17697 32597 17731
rect 32631 17728 32643 17731
rect 35066 17728 35072 17740
rect 32631 17700 35072 17728
rect 32631 17697 32643 17700
rect 32585 17691 32643 17697
rect 35066 17688 35072 17700
rect 35124 17688 35130 17740
rect 43806 17688 43812 17740
rect 43864 17728 43870 17740
rect 44269 17731 44327 17737
rect 44269 17728 44281 17731
rect 43864 17700 44281 17728
rect 43864 17688 43870 17700
rect 44269 17697 44281 17700
rect 44315 17697 44327 17731
rect 44269 17691 44327 17697
rect 32030 17660 32036 17672
rect 30147 17632 30972 17660
rect 31128 17632 32036 17660
rect 30147 17629 30159 17632
rect 30101 17623 30159 17629
rect 30368 17595 30426 17601
rect 30368 17561 30380 17595
rect 30414 17592 30426 17595
rect 30742 17592 30748 17604
rect 30414 17564 30748 17592
rect 30414 17561 30426 17564
rect 30368 17555 30426 17561
rect 30742 17552 30748 17564
rect 30800 17552 30806 17604
rect 30944 17592 30972 17632
rect 32030 17620 32036 17632
rect 32088 17620 32094 17672
rect 34698 17620 34704 17672
rect 34756 17660 34762 17672
rect 35814 17663 35872 17669
rect 35814 17660 35826 17663
rect 34756 17632 35826 17660
rect 34756 17620 34762 17632
rect 35814 17629 35826 17632
rect 35860 17629 35872 17663
rect 36078 17660 36084 17672
rect 35991 17632 36084 17660
rect 35814 17623 35872 17629
rect 36078 17620 36084 17632
rect 36136 17660 36142 17672
rect 37553 17663 37611 17669
rect 37553 17660 37565 17663
rect 36136 17632 37565 17660
rect 36136 17620 36142 17632
rect 37553 17629 37565 17632
rect 37599 17660 37611 17663
rect 38654 17660 38660 17672
rect 37599 17632 38660 17660
rect 37599 17629 37611 17632
rect 37553 17623 37611 17629
rect 38654 17620 38660 17632
rect 38712 17660 38718 17672
rect 39298 17660 39304 17672
rect 38712 17632 39304 17660
rect 38712 17620 38718 17632
rect 39298 17620 39304 17632
rect 39356 17620 39362 17672
rect 40037 17663 40095 17669
rect 40037 17629 40049 17663
rect 40083 17660 40095 17663
rect 40126 17660 40132 17672
rect 40083 17632 40132 17660
rect 40083 17629 40095 17632
rect 40037 17623 40095 17629
rect 40126 17620 40132 17632
rect 40184 17620 40190 17672
rect 43070 17660 43076 17672
rect 43031 17632 43076 17660
rect 43070 17620 43076 17632
rect 43128 17620 43134 17672
rect 54662 17620 54668 17672
rect 54720 17660 54726 17672
rect 55309 17663 55367 17669
rect 55309 17660 55321 17663
rect 54720 17632 55321 17660
rect 54720 17620 54726 17632
rect 55309 17629 55321 17632
rect 55355 17660 55367 17663
rect 55953 17663 56011 17669
rect 55953 17660 55965 17663
rect 55355 17632 55965 17660
rect 55355 17629 55367 17632
rect 55309 17623 55367 17629
rect 55953 17629 55965 17632
rect 55999 17629 56011 17663
rect 55953 17623 56011 17629
rect 31754 17592 31760 17604
rect 30944 17564 31760 17592
rect 31754 17552 31760 17564
rect 31812 17592 31818 17604
rect 32214 17592 32220 17604
rect 31812 17564 32220 17592
rect 31812 17552 31818 17564
rect 32214 17552 32220 17564
rect 32272 17552 32278 17604
rect 32309 17595 32367 17601
rect 32309 17561 32321 17595
rect 32355 17592 32367 17595
rect 32490 17592 32496 17604
rect 32355 17564 32496 17592
rect 32355 17561 32367 17564
rect 32309 17555 32367 17561
rect 32490 17552 32496 17564
rect 32548 17552 32554 17604
rect 33778 17552 33784 17604
rect 33836 17592 33842 17604
rect 33836 17564 34928 17592
rect 33836 17552 33842 17564
rect 31018 17524 31024 17536
rect 27448 17496 31024 17524
rect 23477 17487 23535 17493
rect 31018 17484 31024 17496
rect 31076 17484 31082 17536
rect 31938 17524 31944 17536
rect 31899 17496 31944 17524
rect 31938 17484 31944 17496
rect 31996 17484 32002 17536
rect 34701 17527 34759 17533
rect 34701 17493 34713 17527
rect 34747 17524 34759 17527
rect 34790 17524 34796 17536
rect 34747 17496 34796 17524
rect 34747 17493 34759 17496
rect 34701 17487 34759 17493
rect 34790 17484 34796 17496
rect 34848 17484 34854 17536
rect 34900 17524 34928 17564
rect 36446 17552 36452 17604
rect 36504 17592 36510 17604
rect 36725 17595 36783 17601
rect 36725 17592 36737 17595
rect 36504 17564 36737 17592
rect 36504 17552 36510 17564
rect 36725 17561 36737 17564
rect 36771 17561 36783 17595
rect 36725 17555 36783 17561
rect 37458 17552 37464 17604
rect 37516 17592 37522 17604
rect 37798 17595 37856 17601
rect 37798 17592 37810 17595
rect 37516 17564 37810 17592
rect 37516 17552 37522 17564
rect 37798 17561 37810 17564
rect 37844 17561 37856 17595
rect 43530 17592 43536 17604
rect 37798 17555 37856 17561
rect 37936 17564 43536 17592
rect 37936 17524 37964 17564
rect 43530 17552 43536 17564
rect 43588 17592 43594 17604
rect 44085 17595 44143 17601
rect 44085 17592 44097 17595
rect 43588 17564 44097 17592
rect 43588 17552 43594 17564
rect 44085 17561 44097 17564
rect 44131 17561 44143 17595
rect 67818 17592 67824 17604
rect 44085 17555 44143 17561
rect 55508 17564 67824 17592
rect 38930 17524 38936 17536
rect 34900 17496 37964 17524
rect 38891 17496 38936 17524
rect 38930 17484 38936 17496
rect 38988 17484 38994 17536
rect 39850 17524 39856 17536
rect 39811 17496 39856 17524
rect 39850 17484 39856 17496
rect 39908 17484 39914 17536
rect 41598 17484 41604 17536
rect 41656 17524 41662 17536
rect 41966 17524 41972 17536
rect 41656 17496 41972 17524
rect 41656 17484 41662 17496
rect 41966 17484 41972 17496
rect 42024 17524 42030 17536
rect 42061 17527 42119 17533
rect 42061 17524 42073 17527
rect 42024 17496 42073 17524
rect 42024 17484 42030 17496
rect 42061 17493 42073 17496
rect 42107 17524 42119 17527
rect 42702 17524 42708 17536
rect 42107 17496 42708 17524
rect 42107 17493 42119 17496
rect 42061 17487 42119 17493
rect 42702 17484 42708 17496
rect 42760 17484 42766 17536
rect 43254 17524 43260 17536
rect 43215 17496 43260 17524
rect 43254 17484 43260 17496
rect 43312 17484 43318 17536
rect 43714 17524 43720 17536
rect 43675 17496 43720 17524
rect 43714 17484 43720 17496
rect 43772 17484 43778 17536
rect 44177 17527 44235 17533
rect 44177 17493 44189 17527
rect 44223 17524 44235 17527
rect 45554 17524 45560 17536
rect 44223 17496 45560 17524
rect 44223 17493 44235 17496
rect 44177 17487 44235 17493
rect 45554 17484 45560 17496
rect 45612 17484 45618 17536
rect 55508 17533 55536 17564
rect 67818 17552 67824 17564
rect 67876 17552 67882 17604
rect 55493 17527 55551 17533
rect 55493 17493 55505 17527
rect 55539 17493 55551 17527
rect 55493 17487 55551 17493
rect 1104 17434 68816 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 68816 17434
rect 1104 17360 68816 17382
rect 4617 17323 4675 17329
rect 4617 17289 4629 17323
rect 4663 17289 4675 17323
rect 4617 17283 4675 17289
rect 5077 17323 5135 17329
rect 5077 17289 5089 17323
rect 5123 17320 5135 17323
rect 6454 17320 6460 17332
rect 5123 17292 6460 17320
rect 5123 17289 5135 17292
rect 5077 17283 5135 17289
rect 3973 17187 4031 17193
rect 3973 17153 3985 17187
rect 4019 17184 4031 17187
rect 4632 17184 4660 17283
rect 6454 17280 6460 17292
rect 6512 17280 6518 17332
rect 7650 17320 7656 17332
rect 7611 17292 7656 17320
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 15197 17323 15255 17329
rect 15197 17289 15209 17323
rect 15243 17320 15255 17323
rect 15286 17320 15292 17332
rect 15243 17292 15292 17320
rect 15243 17289 15255 17292
rect 15197 17283 15255 17289
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 19426 17280 19432 17332
rect 19484 17320 19490 17332
rect 20073 17323 20131 17329
rect 20073 17320 20085 17323
rect 19484 17292 20085 17320
rect 19484 17280 19490 17292
rect 20073 17289 20085 17292
rect 20119 17289 20131 17323
rect 20073 17283 20131 17289
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 21913 17323 21971 17329
rect 21913 17320 21925 17323
rect 20864 17292 21925 17320
rect 20864 17280 20870 17292
rect 21913 17289 21925 17292
rect 21959 17289 21971 17323
rect 22554 17320 22560 17332
rect 22515 17292 22560 17320
rect 21913 17283 21971 17289
rect 22554 17280 22560 17292
rect 22612 17280 22618 17332
rect 24397 17323 24455 17329
rect 24397 17289 24409 17323
rect 24443 17320 24455 17323
rect 27706 17320 27712 17332
rect 24443 17292 27712 17320
rect 24443 17289 24455 17292
rect 24397 17283 24455 17289
rect 27706 17280 27712 17292
rect 27764 17280 27770 17332
rect 27893 17323 27951 17329
rect 27893 17289 27905 17323
rect 27939 17289 27951 17323
rect 27893 17283 27951 17289
rect 7558 17252 7564 17264
rect 7116 17224 7564 17252
rect 4019 17156 4660 17184
rect 4985 17187 5043 17193
rect 4019 17153 4031 17156
rect 3973 17147 4031 17153
rect 4985 17153 4997 17187
rect 5031 17184 5043 17187
rect 5718 17184 5724 17196
rect 5031 17156 5724 17184
rect 5031 17153 5043 17156
rect 4985 17147 5043 17153
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 7116 17128 7144 17224
rect 7558 17212 7564 17224
rect 7616 17212 7622 17264
rect 11054 17252 11060 17264
rect 8128 17224 11060 17252
rect 8128 17193 8156 17224
rect 11054 17212 11060 17224
rect 11112 17212 11118 17264
rect 12618 17252 12624 17264
rect 12406 17224 12624 17252
rect 7285 17187 7343 17193
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 8113 17187 8171 17193
rect 8113 17184 8125 17187
rect 7331 17156 8125 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 8113 17153 8125 17156
rect 8159 17153 8171 17187
rect 10778 17184 10784 17196
rect 10739 17156 10784 17184
rect 8113 17147 8171 17153
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17184 11943 17187
rect 12406 17184 12434 17224
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 13265 17255 13323 17261
rect 13265 17221 13277 17255
rect 13311 17252 13323 17255
rect 16574 17252 16580 17264
rect 13311 17224 16580 17252
rect 13311 17221 13323 17224
rect 13265 17215 13323 17221
rect 12526 17184 12532 17196
rect 11931 17156 12434 17184
rect 12487 17156 12532 17184
rect 11931 17153 11943 17156
rect 11885 17147 11943 17153
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12710 17184 12716 17196
rect 12671 17156 12716 17184
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 5261 17119 5319 17125
rect 5261 17085 5273 17119
rect 5307 17116 5319 17119
rect 7098 17116 7104 17128
rect 5307 17088 7104 17116
rect 5307 17085 5319 17088
rect 5261 17079 5319 17085
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 7377 17119 7435 17125
rect 7377 17085 7389 17119
rect 7423 17116 7435 17119
rect 7466 17116 7472 17128
rect 7423 17088 7472 17116
rect 7423 17085 7435 17088
rect 7377 17079 7435 17085
rect 7466 17076 7472 17088
rect 7524 17076 7530 17128
rect 10410 17076 10416 17128
rect 10468 17116 10474 17128
rect 10689 17119 10747 17125
rect 10689 17116 10701 17119
rect 10468 17088 10701 17116
rect 10468 17076 10474 17088
rect 10689 17085 10701 17088
rect 10735 17085 10747 17119
rect 11790 17116 11796 17128
rect 11751 17088 11796 17116
rect 10689 17079 10747 17085
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 12342 17076 12348 17128
rect 12400 17116 12406 17128
rect 13280 17116 13308 17215
rect 16574 17212 16580 17224
rect 16632 17212 16638 17264
rect 19889 17255 19947 17261
rect 17788 17224 19472 17252
rect 15378 17184 15384 17196
rect 15339 17156 15384 17184
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 16850 17184 16856 17196
rect 16811 17156 16856 17184
rect 16850 17144 16856 17156
rect 16908 17144 16914 17196
rect 17678 17116 17684 17128
rect 12400 17088 13308 17116
rect 17639 17088 17684 17116
rect 12400 17076 12406 17088
rect 17678 17076 17684 17088
rect 17736 17076 17742 17128
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 12529 17051 12587 17057
rect 12529 17048 12541 17051
rect 10836 17020 12541 17048
rect 10836 17008 10842 17020
rect 12529 17017 12541 17020
rect 12575 17017 12587 17051
rect 12529 17011 12587 17017
rect 12618 17008 12624 17060
rect 12676 17048 12682 17060
rect 17788 17048 17816 17224
rect 19444 17196 19472 17224
rect 19889 17221 19901 17255
rect 19935 17252 19947 17255
rect 19978 17252 19984 17264
rect 19935 17224 19984 17252
rect 19935 17221 19947 17224
rect 19889 17215 19947 17221
rect 19978 17212 19984 17224
rect 20036 17212 20042 17264
rect 24486 17252 24492 17264
rect 21008 17224 22048 17252
rect 18785 17187 18843 17193
rect 18785 17153 18797 17187
rect 18831 17153 18843 17187
rect 18966 17184 18972 17196
rect 18927 17156 18972 17184
rect 18785 17147 18843 17153
rect 12676 17020 17816 17048
rect 12676 17008 12682 17020
rect 17862 17008 17868 17060
rect 17920 17048 17926 17060
rect 17957 17051 18015 17057
rect 17957 17048 17969 17051
rect 17920 17020 17969 17048
rect 17920 17008 17926 17020
rect 17957 17017 17969 17020
rect 18003 17017 18015 17051
rect 17957 17011 18015 17017
rect 4157 16983 4215 16989
rect 4157 16949 4169 16983
rect 4203 16980 4215 16983
rect 4706 16980 4712 16992
rect 4203 16952 4712 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 10502 16980 10508 16992
rect 10463 16952 10508 16980
rect 10502 16940 10508 16952
rect 10560 16940 10566 16992
rect 11609 16983 11667 16989
rect 11609 16949 11621 16983
rect 11655 16980 11667 16983
rect 11790 16980 11796 16992
rect 11655 16952 11796 16980
rect 11655 16949 11667 16952
rect 11609 16943 11667 16949
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 16666 16980 16672 16992
rect 16627 16952 16672 16980
rect 16666 16940 16672 16952
rect 16724 16940 16730 16992
rect 18141 16983 18199 16989
rect 18141 16949 18153 16983
rect 18187 16980 18199 16983
rect 18230 16980 18236 16992
rect 18187 16952 18236 16980
rect 18187 16949 18199 16952
rect 18141 16943 18199 16949
rect 18230 16940 18236 16952
rect 18288 16940 18294 16992
rect 18800 16980 18828 17147
rect 18966 17144 18972 17156
rect 19024 17144 19030 17196
rect 19150 17144 19156 17196
rect 19208 17184 19214 17196
rect 19245 17187 19303 17193
rect 19245 17184 19257 17187
rect 19208 17156 19257 17184
rect 19208 17144 19214 17156
rect 19245 17153 19257 17156
rect 19291 17153 19303 17187
rect 19245 17147 19303 17153
rect 19426 17144 19432 17196
rect 19484 17184 19490 17196
rect 20070 17184 20076 17196
rect 19484 17156 20076 17184
rect 19484 17144 19490 17156
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 20162 17144 20168 17196
rect 20220 17184 20226 17196
rect 20220 17156 20265 17184
rect 20220 17144 20226 17156
rect 20622 17144 20628 17196
rect 20680 17184 20686 17196
rect 21008 17193 21036 17224
rect 20809 17187 20867 17193
rect 20809 17184 20821 17187
rect 20680 17156 20821 17184
rect 20680 17144 20686 17156
rect 20809 17153 20821 17156
rect 20855 17153 20867 17187
rect 20809 17147 20867 17153
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 21082 17144 21088 17196
rect 21140 17184 21146 17196
rect 22020 17193 22048 17224
rect 22572 17224 24492 17252
rect 21821 17187 21879 17193
rect 21821 17184 21833 17187
rect 21140 17156 21833 17184
rect 21140 17144 21146 17156
rect 21821 17153 21833 17156
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17184 22063 17187
rect 22278 17184 22284 17196
rect 22051 17156 22284 17184
rect 22051 17153 22063 17156
rect 22005 17147 22063 17153
rect 22278 17144 22284 17156
rect 22336 17144 22342 17196
rect 19429 17051 19487 17057
rect 19429 17017 19441 17051
rect 19475 17048 19487 17051
rect 22572 17048 22600 17224
rect 24486 17212 24492 17224
rect 24544 17212 24550 17264
rect 26176 17255 26234 17261
rect 26176 17221 26188 17255
rect 26222 17252 26234 17255
rect 26222 17224 27108 17252
rect 26222 17221 26234 17224
rect 26176 17215 26234 17221
rect 22649 17187 22707 17193
rect 22649 17153 22661 17187
rect 22695 17153 22707 17187
rect 23106 17184 23112 17196
rect 23067 17156 23112 17184
rect 22649 17147 22707 17153
rect 22664 17116 22692 17147
rect 23106 17144 23112 17156
rect 23164 17144 23170 17196
rect 23293 17187 23351 17193
rect 23293 17153 23305 17187
rect 23339 17184 23351 17187
rect 23382 17184 23388 17196
rect 23339 17156 23388 17184
rect 23339 17153 23351 17156
rect 23293 17147 23351 17153
rect 23382 17144 23388 17156
rect 23440 17184 23446 17196
rect 24213 17187 24271 17193
rect 24213 17184 24225 17187
rect 23440 17156 24225 17184
rect 23440 17144 23446 17156
rect 24213 17153 24225 17156
rect 24259 17184 24271 17187
rect 25038 17184 25044 17196
rect 24259 17156 25044 17184
rect 24259 17153 24271 17156
rect 24213 17147 24271 17153
rect 25038 17144 25044 17156
rect 25096 17184 25102 17196
rect 26970 17184 26976 17196
rect 25096 17156 26556 17184
rect 26931 17156 26976 17184
rect 25096 17144 25102 17156
rect 23750 17116 23756 17128
rect 22664 17088 23756 17116
rect 23750 17076 23756 17088
rect 23808 17076 23814 17128
rect 24578 17116 24584 17128
rect 24539 17088 24584 17116
rect 24578 17076 24584 17088
rect 24636 17076 24642 17128
rect 26418 17116 26424 17128
rect 26379 17088 26424 17116
rect 26418 17076 26424 17088
rect 26476 17076 26482 17128
rect 26528 17116 26556 17156
rect 26970 17144 26976 17156
rect 27028 17144 27034 17196
rect 27080 17184 27108 17224
rect 27908 17184 27936 17283
rect 27982 17280 27988 17332
rect 28040 17320 28046 17332
rect 28040 17292 34468 17320
rect 28040 17280 28046 17292
rect 32582 17252 32588 17264
rect 32543 17224 32588 17252
rect 32582 17212 32588 17224
rect 32640 17212 32646 17264
rect 34440 17252 34468 17292
rect 34514 17280 34520 17332
rect 34572 17320 34578 17332
rect 34885 17323 34943 17329
rect 34885 17320 34897 17323
rect 34572 17292 34897 17320
rect 34572 17280 34578 17292
rect 34885 17289 34897 17292
rect 34931 17289 34943 17323
rect 34885 17283 34943 17289
rect 35066 17280 35072 17332
rect 35124 17320 35130 17332
rect 35529 17323 35587 17329
rect 35529 17320 35541 17323
rect 35124 17292 35541 17320
rect 35124 17280 35130 17292
rect 35529 17289 35541 17292
rect 35575 17320 35587 17323
rect 37182 17320 37188 17332
rect 35575 17292 37188 17320
rect 35575 17289 35587 17292
rect 35529 17283 35587 17289
rect 37182 17280 37188 17292
rect 37240 17280 37246 17332
rect 37458 17320 37464 17332
rect 37419 17292 37464 17320
rect 37458 17280 37464 17292
rect 37516 17280 37522 17332
rect 42610 17320 42616 17332
rect 37568 17292 42616 17320
rect 35342 17252 35348 17264
rect 34440 17224 35348 17252
rect 35342 17212 35348 17224
rect 35400 17252 35406 17264
rect 35400 17224 35480 17252
rect 35400 17212 35406 17224
rect 28074 17184 28080 17196
rect 27080 17156 27936 17184
rect 28035 17156 28080 17184
rect 28074 17144 28080 17156
rect 28132 17144 28138 17196
rect 30929 17187 30987 17193
rect 30929 17153 30941 17187
rect 30975 17184 30987 17187
rect 31938 17184 31944 17196
rect 30975 17156 31944 17184
rect 30975 17153 30987 17156
rect 30929 17147 30987 17153
rect 31938 17144 31944 17156
rect 31996 17144 32002 17196
rect 35452 17193 35480 17224
rect 33689 17187 33747 17193
rect 33689 17153 33701 17187
rect 33735 17184 33747 17187
rect 34517 17188 34575 17193
rect 34517 17187 34652 17188
rect 34517 17184 34529 17187
rect 33735 17156 34529 17184
rect 33735 17153 33747 17156
rect 33689 17147 33747 17153
rect 34517 17153 34529 17156
rect 34563 17184 34652 17187
rect 35437 17187 35495 17193
rect 34563 17156 35296 17184
rect 34563 17153 34575 17156
rect 34517 17147 34575 17153
rect 27065 17119 27123 17125
rect 27065 17116 27077 17119
rect 26528 17088 27077 17116
rect 27065 17085 27077 17088
rect 27111 17085 27123 17119
rect 28537 17119 28595 17125
rect 28537 17116 28549 17119
rect 27065 17079 27123 17085
rect 27172 17088 28549 17116
rect 23474 17048 23480 17060
rect 19475 17020 22600 17048
rect 23435 17020 23480 17048
rect 19475 17017 19487 17020
rect 19429 17011 19487 17017
rect 23474 17008 23480 17020
rect 23532 17008 23538 17060
rect 25041 17051 25099 17057
rect 25041 17017 25053 17051
rect 25087 17048 25099 17051
rect 25406 17048 25412 17060
rect 25087 17020 25412 17048
rect 25087 17017 25099 17020
rect 25041 17011 25099 17017
rect 25406 17008 25412 17020
rect 25464 17008 25470 17060
rect 27172 17048 27200 17088
rect 28537 17085 28549 17088
rect 28583 17085 28595 17119
rect 28537 17079 28595 17085
rect 31018 17076 31024 17128
rect 31076 17116 31082 17128
rect 32490 17116 32496 17128
rect 31076 17088 32496 17116
rect 31076 17076 31082 17088
rect 32490 17076 32496 17088
rect 32548 17076 32554 17128
rect 30742 17048 30748 17060
rect 26988 17020 27200 17048
rect 30703 17020 30748 17048
rect 19889 16983 19947 16989
rect 19889 16980 19901 16983
rect 18800 16952 19901 16980
rect 19889 16949 19901 16952
rect 19935 16949 19947 16983
rect 19889 16943 19947 16949
rect 22922 16940 22928 16992
rect 22980 16980 22986 16992
rect 23109 16983 23167 16989
rect 23109 16980 23121 16983
rect 22980 16952 23121 16980
rect 22980 16940 22986 16952
rect 23109 16949 23121 16952
rect 23155 16980 23167 16983
rect 23290 16980 23296 16992
rect 23155 16952 23296 16980
rect 23155 16949 23167 16952
rect 23109 16943 23167 16949
rect 23290 16940 23296 16952
rect 23348 16940 23354 16992
rect 24026 16980 24032 16992
rect 23987 16952 24032 16980
rect 24026 16940 24032 16952
rect 24084 16980 24090 16992
rect 26988 16989 27016 17020
rect 30742 17008 30748 17020
rect 30800 17008 30806 17060
rect 32398 17048 32404 17060
rect 30852 17020 32404 17048
rect 26973 16983 27031 16989
rect 26973 16980 26985 16983
rect 24084 16952 26985 16980
rect 24084 16940 24090 16952
rect 26973 16949 26985 16952
rect 27019 16949 27031 16983
rect 26973 16943 27031 16949
rect 27341 16983 27399 16989
rect 27341 16949 27353 16983
rect 27387 16980 27399 16983
rect 30852 16980 30880 17020
rect 32398 17008 32404 17020
rect 32456 17008 32462 17060
rect 33704 17048 33732 17147
rect 34241 17119 34299 17125
rect 34241 17116 34253 17119
rect 32600 17020 33732 17048
rect 33796 17088 34253 17116
rect 27387 16952 30880 16980
rect 27387 16949 27399 16952
rect 27341 16943 27399 16949
rect 31202 16940 31208 16992
rect 31260 16980 31266 16992
rect 32600 16980 32628 17020
rect 31260 16952 32628 16980
rect 31260 16940 31266 16952
rect 32674 16940 32680 16992
rect 32732 16980 32738 16992
rect 33796 16980 33824 17088
rect 34241 17085 34253 17088
rect 34287 17085 34299 17119
rect 34241 17079 34299 17085
rect 34425 17119 34483 17125
rect 34425 17085 34437 17119
rect 34471 17116 34483 17119
rect 34790 17116 34796 17128
rect 34471 17088 34796 17116
rect 34471 17085 34483 17088
rect 34425 17079 34483 17085
rect 34790 17076 34796 17088
rect 34848 17076 34854 17128
rect 35268 17116 35296 17156
rect 35437 17153 35449 17187
rect 35483 17153 35495 17187
rect 37274 17184 37280 17196
rect 37235 17156 37280 17184
rect 35437 17147 35495 17153
rect 37274 17144 37280 17156
rect 37332 17144 37338 17196
rect 37568 17116 37596 17292
rect 42610 17280 42616 17292
rect 42668 17280 42674 17332
rect 38654 17252 38660 17264
rect 37936 17224 38660 17252
rect 37936 17193 37964 17224
rect 38654 17212 38660 17224
rect 38712 17212 38718 17264
rect 38930 17212 38936 17264
rect 38988 17252 38994 17264
rect 38988 17224 42656 17252
rect 38988 17212 38994 17224
rect 37921 17187 37979 17193
rect 37921 17153 37933 17187
rect 37967 17153 37979 17187
rect 37921 17147 37979 17153
rect 38188 17187 38246 17193
rect 38188 17153 38200 17187
rect 38234 17184 38246 17187
rect 39850 17184 39856 17196
rect 38234 17156 39856 17184
rect 38234 17153 38246 17156
rect 38188 17147 38246 17153
rect 39850 17144 39856 17156
rect 39908 17144 39914 17196
rect 41598 17184 41604 17196
rect 41559 17156 41604 17184
rect 41598 17144 41604 17156
rect 41656 17144 41662 17196
rect 42628 17193 42656 17224
rect 43254 17212 43260 17264
rect 43312 17252 43318 17264
rect 43870 17255 43928 17261
rect 43870 17252 43882 17255
rect 43312 17224 43882 17252
rect 43312 17212 43318 17224
rect 43870 17221 43882 17224
rect 43916 17221 43928 17255
rect 43870 17215 43928 17221
rect 44726 17212 44732 17264
rect 44784 17252 44790 17264
rect 55306 17252 55312 17264
rect 44784 17224 51074 17252
rect 44784 17212 44790 17224
rect 42613 17187 42671 17193
rect 42613 17153 42625 17187
rect 42659 17153 42671 17187
rect 42613 17147 42671 17153
rect 43346 17144 43352 17196
rect 43404 17184 43410 17196
rect 43625 17187 43683 17193
rect 43625 17184 43637 17187
rect 43404 17156 43637 17184
rect 43404 17144 43410 17156
rect 43625 17153 43637 17156
rect 43671 17153 43683 17187
rect 45649 17187 45707 17193
rect 43625 17147 43683 17153
rect 43732 17156 44680 17184
rect 35268 17088 37596 17116
rect 41782 17076 41788 17128
rect 41840 17116 41846 17128
rect 42521 17119 42579 17125
rect 42521 17116 42533 17119
rect 41840 17088 42533 17116
rect 41840 17076 41846 17088
rect 42521 17085 42533 17088
rect 42567 17085 42579 17119
rect 43732 17116 43760 17156
rect 42521 17079 42579 17085
rect 42628 17088 43760 17116
rect 44652 17116 44680 17156
rect 45649 17153 45661 17187
rect 45695 17153 45707 17187
rect 45649 17147 45707 17153
rect 45557 17119 45615 17125
rect 45557 17116 45569 17119
rect 44652 17088 45569 17116
rect 42150 17008 42156 17060
rect 42208 17048 42214 17060
rect 42628 17048 42656 17088
rect 45557 17085 45569 17088
rect 45603 17085 45615 17119
rect 45557 17079 45615 17085
rect 45664 17048 45692 17147
rect 51046 17116 51074 17224
rect 55186 17224 55312 17252
rect 55186 17116 55214 17224
rect 55306 17212 55312 17224
rect 55364 17212 55370 17264
rect 51046 17088 55214 17116
rect 46014 17048 46020 17060
rect 42208 17020 42656 17048
rect 45020 17020 45692 17048
rect 45975 17020 46020 17048
rect 42208 17008 42214 17020
rect 45020 16992 45048 17020
rect 46014 17008 46020 17020
rect 46072 17008 46078 17060
rect 36446 16980 36452 16992
rect 32732 16952 33824 16980
rect 36407 16952 36452 16980
rect 32732 16940 32738 16952
rect 36446 16940 36452 16952
rect 36504 16940 36510 16992
rect 39301 16983 39359 16989
rect 39301 16949 39313 16983
rect 39347 16980 39359 16983
rect 40034 16980 40040 16992
rect 39347 16952 40040 16980
rect 39347 16949 39359 16952
rect 39301 16943 39359 16949
rect 40034 16940 40040 16952
rect 40092 16940 40098 16992
rect 41785 16983 41843 16989
rect 41785 16949 41797 16983
rect 41831 16980 41843 16983
rect 41874 16980 41880 16992
rect 41831 16952 41880 16980
rect 41831 16949 41843 16952
rect 41785 16943 41843 16949
rect 41874 16940 41880 16952
rect 41932 16940 41938 16992
rect 42889 16983 42947 16989
rect 42889 16949 42901 16983
rect 42935 16980 42947 16983
rect 44910 16980 44916 16992
rect 42935 16952 44916 16980
rect 42935 16949 42947 16952
rect 42889 16943 42947 16949
rect 44910 16940 44916 16952
rect 44968 16940 44974 16992
rect 45002 16940 45008 16992
rect 45060 16980 45066 16992
rect 45060 16952 45105 16980
rect 45060 16940 45066 16952
rect 1104 16890 68816 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 65654 16890
rect 65706 16838 65718 16890
rect 65770 16838 65782 16890
rect 65834 16838 65846 16890
rect 65898 16838 65910 16890
rect 65962 16838 68816 16890
rect 1104 16816 68816 16838
rect 4614 16776 4620 16788
rect 4356 16748 4620 16776
rect 4356 16652 4384 16748
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 5718 16776 5724 16788
rect 5679 16748 5724 16776
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 7285 16779 7343 16785
rect 7285 16745 7297 16779
rect 7331 16776 7343 16779
rect 8941 16779 8999 16785
rect 8941 16776 8953 16779
rect 7331 16748 8953 16776
rect 7331 16745 7343 16748
rect 7285 16739 7343 16745
rect 8941 16745 8953 16748
rect 8987 16745 8999 16779
rect 8941 16739 8999 16745
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 11517 16779 11575 16785
rect 11517 16776 11529 16779
rect 11204 16748 11529 16776
rect 11204 16736 11210 16748
rect 11517 16745 11529 16748
rect 11563 16745 11575 16779
rect 12618 16776 12624 16788
rect 12579 16748 12624 16776
rect 11517 16739 11575 16745
rect 12618 16736 12624 16748
rect 12676 16736 12682 16788
rect 16482 16736 16488 16788
rect 16540 16776 16546 16788
rect 16540 16748 16896 16776
rect 16540 16736 16546 16748
rect 9674 16668 9680 16720
rect 9732 16708 9738 16720
rect 10962 16708 10968 16720
rect 9732 16680 10968 16708
rect 9732 16668 9738 16680
rect 10962 16668 10968 16680
rect 11020 16708 11026 16720
rect 12434 16708 12440 16720
rect 11020 16680 12440 16708
rect 11020 16668 11026 16680
rect 12434 16668 12440 16680
rect 12492 16668 12498 16720
rect 4338 16640 4344 16652
rect 4251 16612 4344 16640
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 6914 16640 6920 16652
rect 6875 16612 6920 16640
rect 6914 16600 6920 16612
rect 6972 16600 6978 16652
rect 8110 16640 8116 16652
rect 8071 16612 8116 16640
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 9030 16640 9036 16652
rect 8991 16612 9036 16640
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 11609 16643 11667 16649
rect 11609 16640 11621 16643
rect 10520 16612 11621 16640
rect 7006 16572 7012 16584
rect 6967 16544 7012 16572
rect 7006 16532 7012 16544
rect 7064 16532 7070 16584
rect 7650 16532 7656 16584
rect 7708 16572 7714 16584
rect 8205 16575 8263 16581
rect 8205 16572 8217 16575
rect 7708 16544 8217 16572
rect 7708 16532 7714 16544
rect 8205 16541 8217 16544
rect 8251 16541 8263 16575
rect 9214 16572 9220 16584
rect 9175 16544 9220 16572
rect 8205 16535 8263 16541
rect 9214 16532 9220 16544
rect 9272 16532 9278 16584
rect 10520 16572 10548 16612
rect 11609 16609 11621 16612
rect 11655 16609 11667 16643
rect 16868 16640 16896 16748
rect 18230 16736 18236 16788
rect 18288 16776 18294 16788
rect 18874 16776 18880 16788
rect 18288 16748 18880 16776
rect 18288 16736 18294 16748
rect 18874 16736 18880 16748
rect 18932 16776 18938 16788
rect 19245 16779 19303 16785
rect 19245 16776 19257 16779
rect 18932 16748 19257 16776
rect 18932 16736 18938 16748
rect 19245 16745 19257 16748
rect 19291 16745 19303 16779
rect 23382 16776 23388 16788
rect 23343 16748 23388 16776
rect 19245 16739 19303 16745
rect 23382 16736 23388 16748
rect 23440 16736 23446 16788
rect 26418 16736 26424 16788
rect 26476 16776 26482 16788
rect 26476 16748 30972 16776
rect 26476 16736 26482 16748
rect 17034 16668 17040 16720
rect 17092 16708 17098 16720
rect 17678 16708 17684 16720
rect 17092 16680 17684 16708
rect 17092 16668 17098 16680
rect 17678 16668 17684 16680
rect 17736 16708 17742 16720
rect 17957 16711 18015 16717
rect 17957 16708 17969 16711
rect 17736 16680 17969 16708
rect 17736 16668 17742 16680
rect 17957 16677 17969 16680
rect 18003 16677 18015 16711
rect 17957 16671 18015 16677
rect 18141 16711 18199 16717
rect 18141 16677 18153 16711
rect 18187 16708 18199 16711
rect 19150 16708 19156 16720
rect 18187 16680 19156 16708
rect 18187 16677 18199 16680
rect 18141 16671 18199 16677
rect 19150 16668 19156 16680
rect 19208 16708 19214 16720
rect 20901 16711 20959 16717
rect 20901 16708 20913 16711
rect 19208 16680 19380 16708
rect 19208 16668 19214 16680
rect 19352 16649 19380 16680
rect 19444 16680 20913 16708
rect 19337 16643 19395 16649
rect 16868 16612 19288 16640
rect 11609 16603 11667 16609
rect 9416 16544 10548 16572
rect 4608 16507 4666 16513
rect 4608 16473 4620 16507
rect 4654 16504 4666 16507
rect 4706 16504 4712 16516
rect 4654 16476 4712 16504
rect 4654 16473 4666 16476
rect 4608 16467 4666 16473
rect 4706 16464 4712 16476
rect 4764 16464 4770 16516
rect 8941 16507 8999 16513
rect 8941 16473 8953 16507
rect 8987 16504 8999 16507
rect 9122 16504 9128 16516
rect 8987 16476 9128 16504
rect 8987 16473 8999 16476
rect 8941 16467 8999 16473
rect 9122 16464 9128 16476
rect 9180 16464 9186 16516
rect 7834 16436 7840 16448
rect 7795 16408 7840 16436
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 9416 16445 9444 16544
rect 11422 16532 11428 16584
rect 11480 16572 11486 16584
rect 11517 16575 11575 16581
rect 11517 16572 11529 16575
rect 11480 16544 11529 16572
rect 11480 16532 11486 16544
rect 11517 16541 11529 16544
rect 11563 16541 11575 16575
rect 11790 16572 11796 16584
rect 11751 16544 11796 16572
rect 11517 16535 11575 16541
rect 11790 16532 11796 16544
rect 11848 16532 11854 16584
rect 15746 16532 15752 16584
rect 15804 16572 15810 16584
rect 15841 16575 15899 16581
rect 15841 16572 15853 16575
rect 15804 16544 15853 16572
rect 15804 16532 15810 16544
rect 15841 16541 15853 16544
rect 15887 16572 15899 16575
rect 18138 16572 18144 16584
rect 15887 16544 18144 16572
rect 15887 16541 15899 16544
rect 15841 16535 15899 16541
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 19260 16572 19288 16612
rect 19337 16609 19349 16643
rect 19383 16609 19395 16643
rect 19337 16603 19395 16609
rect 19444 16572 19472 16680
rect 20901 16677 20913 16680
rect 20947 16708 20959 16711
rect 23106 16708 23112 16720
rect 20947 16680 23112 16708
rect 20947 16677 20959 16680
rect 20901 16671 20959 16677
rect 23106 16668 23112 16680
rect 23164 16708 23170 16720
rect 23164 16680 23336 16708
rect 23164 16668 23170 16680
rect 22186 16640 22192 16652
rect 22147 16612 22192 16640
rect 22186 16600 22192 16612
rect 22244 16600 22250 16652
rect 23308 16649 23336 16680
rect 23293 16643 23351 16649
rect 23293 16609 23305 16643
rect 23339 16609 23351 16643
rect 25130 16640 25136 16652
rect 25091 16612 25136 16640
rect 23293 16603 23351 16609
rect 25130 16600 25136 16612
rect 25188 16600 25194 16652
rect 27540 16649 27568 16748
rect 30944 16708 30972 16748
rect 32398 16736 32404 16788
rect 32456 16776 32462 16788
rect 36446 16776 36452 16788
rect 32456 16748 36452 16776
rect 32456 16736 32462 16748
rect 36446 16736 36452 16748
rect 36504 16736 36510 16788
rect 37274 16776 37280 16788
rect 37235 16748 37280 16776
rect 37274 16736 37280 16748
rect 37332 16736 37338 16788
rect 38562 16736 38568 16788
rect 38620 16776 38626 16788
rect 42426 16776 42432 16788
rect 38620 16748 42288 16776
rect 42387 16748 42432 16776
rect 38620 16736 38626 16748
rect 31754 16708 31760 16720
rect 30944 16680 31760 16708
rect 30944 16649 30972 16680
rect 31754 16668 31760 16680
rect 31812 16668 31818 16720
rect 31849 16711 31907 16717
rect 31849 16677 31861 16711
rect 31895 16708 31907 16711
rect 34514 16708 34520 16720
rect 31895 16680 33640 16708
rect 31895 16677 31907 16680
rect 31849 16671 31907 16677
rect 27525 16643 27583 16649
rect 27525 16609 27537 16643
rect 27571 16609 27583 16643
rect 27525 16603 27583 16609
rect 30929 16643 30987 16649
rect 30929 16609 30941 16643
rect 30975 16609 30987 16643
rect 30929 16603 30987 16609
rect 32674 16600 32680 16652
rect 32732 16640 32738 16652
rect 33505 16643 33563 16649
rect 33505 16640 33517 16643
rect 32732 16612 33517 16640
rect 32732 16600 32738 16612
rect 33505 16609 33517 16612
rect 33551 16609 33563 16643
rect 33505 16603 33563 16609
rect 19260 16544 19472 16572
rect 19521 16575 19579 16581
rect 19521 16541 19533 16575
rect 19567 16572 19579 16575
rect 19978 16572 19984 16584
rect 19567 16544 19984 16572
rect 19567 16541 19579 16544
rect 19521 16535 19579 16541
rect 19978 16532 19984 16544
rect 20036 16532 20042 16584
rect 21634 16532 21640 16584
rect 21692 16572 21698 16584
rect 21913 16575 21971 16581
rect 21913 16572 21925 16575
rect 21692 16544 21925 16572
rect 21692 16532 21698 16544
rect 21913 16541 21925 16544
rect 21959 16541 21971 16575
rect 23566 16572 23572 16584
rect 23479 16544 23572 16572
rect 21913 16535 21971 16541
rect 23566 16532 23572 16544
rect 23624 16572 23630 16584
rect 24854 16572 24860 16584
rect 23624 16544 24624 16572
rect 24815 16544 24860 16572
rect 23624 16532 23630 16544
rect 24596 16516 24624 16544
rect 24854 16532 24860 16544
rect 24912 16532 24918 16584
rect 27706 16532 27712 16584
rect 27764 16572 27770 16584
rect 28169 16575 28227 16581
rect 28169 16572 28181 16575
rect 27764 16544 28181 16572
rect 27764 16532 27770 16544
rect 28169 16541 28181 16544
rect 28215 16541 28227 16575
rect 28169 16535 28227 16541
rect 28813 16575 28871 16581
rect 28813 16541 28825 16575
rect 28859 16572 28871 16575
rect 29454 16572 29460 16584
rect 28859 16544 29460 16572
rect 28859 16541 28871 16544
rect 28813 16535 28871 16541
rect 29454 16532 29460 16544
rect 29512 16532 29518 16584
rect 32306 16572 32312 16584
rect 32267 16544 32312 16572
rect 32306 16532 32312 16544
rect 32364 16532 32370 16584
rect 33612 16572 33640 16680
rect 33704 16680 34520 16708
rect 33704 16649 33732 16680
rect 34514 16668 34520 16680
rect 34572 16708 34578 16720
rect 34701 16711 34759 16717
rect 34701 16708 34713 16711
rect 34572 16680 34713 16708
rect 34572 16668 34578 16680
rect 34701 16677 34713 16680
rect 34747 16677 34759 16711
rect 38930 16708 38936 16720
rect 34701 16671 34759 16677
rect 37752 16680 38936 16708
rect 33689 16643 33747 16649
rect 33689 16609 33701 16643
rect 33735 16609 33747 16643
rect 36078 16640 36084 16652
rect 36039 16612 36084 16640
rect 33689 16603 33747 16609
rect 36078 16600 36084 16612
rect 36136 16600 36142 16652
rect 37752 16649 37780 16680
rect 38930 16668 38936 16680
rect 38988 16668 38994 16720
rect 40405 16711 40463 16717
rect 40405 16677 40417 16711
rect 40451 16708 40463 16711
rect 41417 16711 41475 16717
rect 40451 16680 41000 16708
rect 40451 16677 40463 16680
rect 40405 16671 40463 16677
rect 37737 16643 37795 16649
rect 37737 16609 37749 16643
rect 37783 16609 37795 16643
rect 37737 16603 37795 16609
rect 37826 16600 37832 16652
rect 37884 16640 37890 16652
rect 37921 16643 37979 16649
rect 37921 16640 37933 16643
rect 37884 16612 37933 16640
rect 37884 16600 37890 16612
rect 37921 16609 37933 16612
rect 37967 16640 37979 16643
rect 38562 16640 38568 16652
rect 37967 16612 38568 16640
rect 37967 16609 37979 16612
rect 37921 16603 37979 16609
rect 38562 16600 38568 16612
rect 38620 16600 38626 16652
rect 38749 16643 38807 16649
rect 38749 16609 38761 16643
rect 38795 16640 38807 16643
rect 40129 16643 40187 16649
rect 38795 16612 39896 16640
rect 38795 16609 38807 16612
rect 38749 16603 38807 16609
rect 33778 16572 33784 16584
rect 33612 16544 33784 16572
rect 33778 16532 33784 16544
rect 33836 16532 33842 16584
rect 39868 16572 39896 16612
rect 40129 16609 40141 16643
rect 40175 16640 40187 16643
rect 40310 16640 40316 16652
rect 40175 16612 40316 16640
rect 40175 16609 40187 16612
rect 40129 16603 40187 16609
rect 40310 16600 40316 16612
rect 40368 16600 40374 16652
rect 40972 16649 41000 16680
rect 41417 16677 41429 16711
rect 41463 16677 41475 16711
rect 41417 16671 41475 16677
rect 40957 16643 41015 16649
rect 40957 16609 40969 16643
rect 41003 16609 41015 16643
rect 41432 16640 41460 16671
rect 41506 16668 41512 16720
rect 41564 16708 41570 16720
rect 41877 16711 41935 16717
rect 41877 16708 41889 16711
rect 41564 16680 41889 16708
rect 41564 16668 41570 16680
rect 41877 16677 41889 16680
rect 41923 16677 41935 16711
rect 42260 16708 42288 16748
rect 42426 16736 42432 16748
rect 42484 16736 42490 16788
rect 43070 16736 43076 16788
rect 43128 16776 43134 16788
rect 43257 16779 43315 16785
rect 43257 16776 43269 16779
rect 43128 16748 43269 16776
rect 43128 16736 43134 16748
rect 43257 16745 43269 16748
rect 43303 16745 43315 16779
rect 43806 16776 43812 16788
rect 43257 16739 43315 16745
rect 43456 16748 43812 16776
rect 43456 16708 43484 16748
rect 43806 16736 43812 16748
rect 43864 16736 43870 16788
rect 42260 16680 43484 16708
rect 43640 16680 45140 16708
rect 41877 16671 41935 16677
rect 43640 16640 43668 16680
rect 41432 16612 43668 16640
rect 43717 16643 43775 16649
rect 40957 16603 41015 16609
rect 43717 16609 43729 16643
rect 43763 16609 43775 16643
rect 43717 16603 43775 16609
rect 40034 16572 40040 16584
rect 39868 16544 40040 16572
rect 40034 16532 40040 16544
rect 40092 16532 40098 16584
rect 41046 16572 41052 16584
rect 41007 16544 41052 16572
rect 41046 16532 41052 16544
rect 41104 16532 41110 16584
rect 42061 16575 42119 16581
rect 42061 16572 42073 16575
rect 41386 16544 42073 16572
rect 16108 16507 16166 16513
rect 16108 16473 16120 16507
rect 16154 16504 16166 16507
rect 16666 16504 16672 16516
rect 16154 16476 16672 16504
rect 16154 16473 16166 16476
rect 16108 16467 16166 16473
rect 16666 16464 16672 16476
rect 16724 16464 16730 16516
rect 17681 16507 17739 16513
rect 17681 16473 17693 16507
rect 17727 16504 17739 16507
rect 17862 16504 17868 16516
rect 17727 16476 17868 16504
rect 17727 16473 17739 16476
rect 17681 16467 17739 16473
rect 17862 16464 17868 16476
rect 17920 16464 17926 16516
rect 19245 16507 19303 16513
rect 19245 16473 19257 16507
rect 19291 16504 19303 16507
rect 19334 16504 19340 16516
rect 19291 16476 19340 16504
rect 19291 16473 19303 16476
rect 19245 16467 19303 16473
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 24578 16464 24584 16516
rect 24636 16504 24642 16516
rect 25038 16504 25044 16516
rect 24636 16476 25044 16504
rect 24636 16464 24642 16476
rect 25038 16464 25044 16476
rect 25096 16464 25102 16516
rect 27280 16507 27338 16513
rect 27280 16473 27292 16507
rect 27326 16504 27338 16507
rect 30662 16507 30720 16513
rect 30662 16504 30674 16507
rect 27326 16476 28028 16504
rect 27326 16473 27338 16476
rect 27280 16467 27338 16473
rect 9401 16439 9459 16445
rect 9401 16405 9413 16439
rect 9447 16405 9459 16439
rect 9401 16399 9459 16405
rect 10594 16396 10600 16448
rect 10652 16436 10658 16448
rect 11422 16436 11428 16448
rect 10652 16408 11428 16436
rect 10652 16396 10658 16408
rect 11422 16396 11428 16408
rect 11480 16396 11486 16448
rect 11977 16439 12035 16445
rect 11977 16405 11989 16439
rect 12023 16436 12035 16439
rect 12158 16436 12164 16448
rect 12023 16408 12164 16436
rect 12023 16405 12035 16408
rect 11977 16399 12035 16405
rect 12158 16396 12164 16408
rect 12216 16396 12222 16448
rect 17034 16396 17040 16448
rect 17092 16436 17098 16448
rect 17221 16439 17279 16445
rect 17221 16436 17233 16439
rect 17092 16408 17233 16436
rect 17092 16396 17098 16408
rect 17221 16405 17233 16408
rect 17267 16405 17279 16439
rect 17221 16399 17279 16405
rect 19705 16439 19763 16445
rect 19705 16405 19717 16439
rect 19751 16436 19763 16439
rect 20070 16436 20076 16448
rect 19751 16408 20076 16436
rect 19751 16405 19763 16408
rect 19705 16399 19763 16405
rect 20070 16396 20076 16408
rect 20128 16396 20134 16448
rect 22830 16396 22836 16448
rect 22888 16436 22894 16448
rect 23017 16439 23075 16445
rect 23017 16436 23029 16439
rect 22888 16408 23029 16436
rect 22888 16396 22894 16408
rect 23017 16405 23029 16408
rect 23063 16405 23075 16439
rect 26142 16436 26148 16448
rect 26103 16408 26148 16436
rect 23017 16399 23075 16405
rect 26142 16396 26148 16408
rect 26200 16396 26206 16448
rect 28000 16445 28028 16476
rect 29012 16476 30674 16504
rect 29012 16445 29040 16476
rect 30662 16473 30674 16476
rect 30708 16473 30720 16507
rect 30662 16467 30720 16473
rect 33962 16464 33968 16516
rect 34020 16504 34026 16516
rect 35814 16507 35872 16513
rect 35814 16504 35826 16507
rect 34020 16476 35826 16504
rect 34020 16464 34026 16476
rect 35814 16473 35826 16476
rect 35860 16473 35872 16507
rect 35814 16467 35872 16473
rect 27985 16439 28043 16445
rect 27985 16405 27997 16439
rect 28031 16405 28043 16439
rect 27985 16399 28043 16405
rect 28997 16439 29055 16445
rect 28997 16405 29009 16439
rect 29043 16405 29055 16439
rect 28997 16399 29055 16405
rect 29549 16439 29607 16445
rect 29549 16405 29561 16439
rect 29595 16436 29607 16439
rect 29914 16436 29920 16448
rect 29595 16408 29920 16436
rect 29595 16405 29607 16408
rect 29549 16399 29607 16405
rect 29914 16396 29920 16408
rect 29972 16396 29978 16448
rect 32490 16436 32496 16448
rect 32451 16408 32496 16436
rect 32490 16396 32496 16408
rect 32548 16396 32554 16448
rect 34146 16436 34152 16448
rect 34107 16408 34152 16436
rect 34146 16396 34152 16408
rect 34204 16396 34210 16448
rect 34422 16396 34428 16448
rect 34480 16436 34486 16448
rect 36725 16439 36783 16445
rect 36725 16436 36737 16439
rect 34480 16408 36737 16436
rect 34480 16396 34486 16408
rect 36725 16405 36737 16408
rect 36771 16436 36783 16439
rect 37645 16439 37703 16445
rect 37645 16436 37657 16439
rect 36771 16408 37657 16436
rect 36771 16405 36783 16408
rect 36725 16399 36783 16405
rect 37645 16405 37657 16408
rect 37691 16436 37703 16439
rect 38102 16436 38108 16448
rect 37691 16408 38108 16436
rect 37691 16405 37703 16408
rect 37645 16399 37703 16405
rect 38102 16396 38108 16408
rect 38160 16396 38166 16448
rect 38838 16436 38844 16448
rect 38799 16408 38844 16436
rect 38838 16396 38844 16408
rect 38896 16396 38902 16448
rect 39209 16439 39267 16445
rect 39209 16405 39221 16439
rect 39255 16436 39267 16439
rect 40126 16436 40132 16448
rect 39255 16408 40132 16436
rect 39255 16405 39267 16408
rect 39209 16399 39267 16405
rect 40126 16396 40132 16408
rect 40184 16396 40190 16448
rect 40402 16396 40408 16448
rect 40460 16436 40466 16448
rect 41386 16436 41414 16544
rect 42061 16541 42073 16544
rect 42107 16541 42119 16575
rect 42061 16535 42119 16541
rect 42150 16532 42156 16584
rect 42208 16572 42214 16584
rect 43732 16572 43760 16603
rect 43806 16600 43812 16652
rect 43864 16640 43870 16652
rect 45002 16640 45008 16652
rect 43864 16612 43909 16640
rect 44008 16612 45008 16640
rect 43864 16600 43870 16612
rect 44008 16572 44036 16612
rect 45002 16600 45008 16612
rect 45060 16600 45066 16652
rect 45112 16649 45140 16680
rect 45186 16668 45192 16720
rect 45244 16708 45250 16720
rect 46017 16711 46075 16717
rect 46017 16708 46029 16711
rect 45244 16680 45289 16708
rect 45388 16680 46029 16708
rect 45244 16668 45250 16680
rect 45097 16643 45155 16649
rect 45097 16609 45109 16643
rect 45143 16609 45155 16643
rect 45097 16603 45155 16609
rect 45281 16643 45339 16649
rect 45281 16609 45293 16643
rect 45327 16640 45339 16643
rect 45388 16640 45416 16680
rect 46017 16677 46029 16680
rect 46063 16677 46075 16711
rect 46017 16671 46075 16677
rect 45554 16640 45560 16652
rect 45327 16612 45416 16640
rect 45515 16612 45560 16640
rect 45327 16609 45339 16612
rect 45281 16603 45339 16609
rect 45554 16600 45560 16612
rect 45612 16640 45618 16652
rect 45612 16612 46244 16640
rect 45612 16600 45618 16612
rect 45370 16572 45376 16584
rect 42208 16544 42253 16572
rect 43732 16544 44036 16572
rect 45331 16544 45376 16572
rect 42208 16532 42214 16544
rect 45370 16532 45376 16544
rect 45428 16532 45434 16584
rect 46014 16572 46020 16584
rect 45975 16544 46020 16572
rect 46014 16532 46020 16544
rect 46072 16532 46078 16584
rect 46216 16581 46244 16612
rect 46201 16575 46259 16581
rect 46201 16541 46213 16575
rect 46247 16541 46259 16575
rect 46201 16535 46259 16541
rect 46293 16575 46351 16581
rect 46293 16541 46305 16575
rect 46339 16541 46351 16575
rect 46293 16535 46351 16541
rect 42610 16464 42616 16516
rect 42668 16504 42674 16516
rect 43625 16507 43683 16513
rect 43625 16504 43637 16507
rect 42668 16476 43637 16504
rect 42668 16464 42674 16476
rect 43625 16473 43637 16476
rect 43671 16473 43683 16507
rect 43625 16467 43683 16473
rect 44910 16464 44916 16516
rect 44968 16504 44974 16516
rect 45189 16507 45247 16513
rect 45189 16504 45201 16507
rect 44968 16476 45201 16504
rect 44968 16464 44974 16476
rect 45189 16473 45201 16476
rect 45235 16473 45247 16507
rect 45388 16504 45416 16532
rect 46308 16504 46336 16535
rect 45388 16476 46336 16504
rect 45189 16467 45247 16473
rect 40460 16408 41414 16436
rect 42245 16439 42303 16445
rect 40460 16396 40466 16408
rect 42245 16405 42257 16439
rect 42291 16436 42303 16439
rect 43254 16436 43260 16448
rect 42291 16408 43260 16436
rect 42291 16405 42303 16408
rect 42245 16399 42303 16405
rect 43254 16396 43260 16408
rect 43312 16396 43318 16448
rect 1104 16346 68816 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 68816 16346
rect 1104 16272 68816 16294
rect 5813 16235 5871 16241
rect 5813 16201 5825 16235
rect 5859 16232 5871 16235
rect 6733 16235 6791 16241
rect 6733 16232 6745 16235
rect 5859 16204 6745 16232
rect 5859 16201 5871 16204
rect 5813 16195 5871 16201
rect 6733 16201 6745 16204
rect 6779 16232 6791 16235
rect 7466 16232 7472 16244
rect 6779 16204 7472 16232
rect 6779 16201 6791 16204
rect 6733 16195 6791 16201
rect 7466 16192 7472 16204
rect 7524 16192 7530 16244
rect 8113 16235 8171 16241
rect 8113 16201 8125 16235
rect 8159 16232 8171 16235
rect 9030 16232 9036 16244
rect 8159 16204 9036 16232
rect 8159 16201 8171 16204
rect 8113 16195 8171 16201
rect 9030 16192 9036 16204
rect 9088 16192 9094 16244
rect 10965 16235 11023 16241
rect 10965 16201 10977 16235
rect 11011 16232 11023 16235
rect 11146 16232 11152 16244
rect 11011 16204 11152 16232
rect 11011 16201 11023 16204
rect 10965 16195 11023 16201
rect 11146 16192 11152 16204
rect 11204 16192 11210 16244
rect 14829 16235 14887 16241
rect 14829 16201 14841 16235
rect 14875 16232 14887 16235
rect 15102 16232 15108 16244
rect 14875 16204 15108 16232
rect 14875 16201 14887 16204
rect 14829 16195 14887 16201
rect 15102 16192 15108 16204
rect 15160 16232 15166 16244
rect 15749 16235 15807 16241
rect 15749 16232 15761 16235
rect 15160 16204 15761 16232
rect 15160 16192 15166 16204
rect 15749 16201 15761 16204
rect 15795 16201 15807 16235
rect 18230 16232 18236 16244
rect 15749 16195 15807 16201
rect 17328 16204 18236 16232
rect 11514 16124 11520 16176
rect 11572 16164 11578 16176
rect 11974 16164 11980 16176
rect 11572 16136 11980 16164
rect 11572 16124 11578 16136
rect 11974 16124 11980 16136
rect 12032 16124 12038 16176
rect 12802 16164 12808 16176
rect 12715 16136 12808 16164
rect 12802 16124 12808 16136
rect 12860 16164 12866 16176
rect 17328 16173 17356 16204
rect 18230 16192 18236 16204
rect 18288 16232 18294 16244
rect 18785 16235 18843 16241
rect 18785 16232 18797 16235
rect 18288 16204 18797 16232
rect 18288 16192 18294 16204
rect 18785 16201 18797 16204
rect 18831 16232 18843 16235
rect 20438 16232 20444 16244
rect 18831 16204 20444 16232
rect 18831 16201 18843 16204
rect 18785 16195 18843 16201
rect 20438 16192 20444 16204
rect 20496 16192 20502 16244
rect 22189 16235 22247 16241
rect 22189 16201 22201 16235
rect 22235 16232 22247 16235
rect 22741 16235 22799 16241
rect 22741 16232 22753 16235
rect 22235 16204 22753 16232
rect 22235 16201 22247 16204
rect 22189 16195 22247 16201
rect 22741 16201 22753 16204
rect 22787 16232 22799 16235
rect 23566 16232 23572 16244
rect 22787 16204 23572 16232
rect 22787 16201 22799 16204
rect 22741 16195 22799 16201
rect 23566 16192 23572 16204
rect 23624 16192 23630 16244
rect 24673 16235 24731 16241
rect 24673 16201 24685 16235
rect 24719 16232 24731 16235
rect 25406 16232 25412 16244
rect 24719 16204 25412 16232
rect 24719 16201 24731 16204
rect 24673 16195 24731 16201
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 26142 16192 26148 16244
rect 26200 16232 26206 16244
rect 27249 16235 27307 16241
rect 27249 16232 27261 16235
rect 26200 16204 27261 16232
rect 26200 16192 26206 16204
rect 27249 16201 27261 16204
rect 27295 16201 27307 16235
rect 27706 16232 27712 16244
rect 27667 16204 27712 16232
rect 27249 16195 27307 16201
rect 13357 16167 13415 16173
rect 13357 16164 13369 16167
rect 12860 16136 13369 16164
rect 12860 16124 12866 16136
rect 13357 16133 13369 16136
rect 13403 16164 13415 16167
rect 17313 16167 17371 16173
rect 17313 16164 17325 16167
rect 13403 16136 17325 16164
rect 13403 16133 13415 16136
rect 13357 16127 13415 16133
rect 17313 16133 17325 16136
rect 17359 16133 17371 16167
rect 17313 16127 17371 16133
rect 22830 16124 22836 16176
rect 22888 16164 22894 16176
rect 23293 16167 23351 16173
rect 23293 16164 23305 16167
rect 22888 16136 23305 16164
rect 22888 16124 22894 16136
rect 23293 16133 23305 16136
rect 23339 16133 23351 16167
rect 27264 16164 27292 16195
rect 27706 16192 27712 16204
rect 27764 16192 27770 16244
rect 29454 16232 29460 16244
rect 29415 16204 29460 16232
rect 29454 16192 29460 16204
rect 29512 16192 29518 16244
rect 29914 16232 29920 16244
rect 29875 16204 29920 16232
rect 29914 16192 29920 16204
rect 29972 16192 29978 16244
rect 32306 16232 32312 16244
rect 32267 16204 32312 16232
rect 32306 16192 32312 16204
rect 32364 16192 32370 16244
rect 33962 16232 33968 16244
rect 33923 16204 33968 16232
rect 33962 16192 33968 16204
rect 34020 16192 34026 16244
rect 42610 16192 42616 16244
rect 42668 16232 42674 16244
rect 42705 16235 42763 16241
rect 42705 16232 42717 16235
rect 42668 16204 42717 16232
rect 42668 16192 42674 16204
rect 42705 16201 42717 16204
rect 42751 16201 42763 16235
rect 42705 16195 42763 16201
rect 43441 16235 43499 16241
rect 43441 16201 43453 16235
rect 43487 16201 43499 16235
rect 43441 16195 43499 16201
rect 45281 16235 45339 16241
rect 45281 16201 45293 16235
rect 45327 16232 45339 16235
rect 45554 16232 45560 16244
rect 45327 16204 45560 16232
rect 45327 16201 45339 16204
rect 45281 16195 45339 16201
rect 31573 16167 31631 16173
rect 27264 16136 28212 16164
rect 23293 16127 23351 16133
rect 4338 16056 4344 16108
rect 4396 16096 4402 16108
rect 4433 16099 4491 16105
rect 4433 16096 4445 16099
rect 4396 16068 4445 16096
rect 4396 16056 4402 16068
rect 4433 16065 4445 16068
rect 4479 16065 4491 16099
rect 4433 16059 4491 16065
rect 4700 16099 4758 16105
rect 4700 16065 4712 16099
rect 4746 16096 4758 16099
rect 5166 16096 5172 16108
rect 4746 16068 5172 16096
rect 4746 16065 4758 16068
rect 4700 16059 4758 16065
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 7742 16096 7748 16108
rect 7703 16068 7748 16096
rect 7742 16056 7748 16068
rect 7800 16056 7806 16108
rect 10594 16096 10600 16108
rect 10555 16068 10600 16096
rect 10594 16056 10600 16068
rect 10652 16056 10658 16108
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 16942 16096 16948 16108
rect 15703 16068 16948 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 16942 16056 16948 16068
rect 17000 16056 17006 16108
rect 24762 16096 24768 16108
rect 24723 16068 24768 16096
rect 24762 16056 24768 16068
rect 24820 16096 24826 16108
rect 28184 16105 28212 16136
rect 31573 16133 31585 16167
rect 31619 16164 31631 16167
rect 32677 16167 32735 16173
rect 32677 16164 32689 16167
rect 31619 16136 32689 16164
rect 31619 16133 31631 16136
rect 31573 16127 31631 16133
rect 32677 16133 32689 16136
rect 32723 16164 32735 16167
rect 33502 16164 33508 16176
rect 32723 16136 33508 16164
rect 32723 16133 32735 16136
rect 32677 16127 32735 16133
rect 33502 16124 33508 16136
rect 33560 16164 33566 16176
rect 34422 16164 34428 16176
rect 33560 16136 34428 16164
rect 33560 16124 33566 16136
rect 34422 16124 34428 16136
rect 34480 16124 34486 16176
rect 43456 16164 43484 16195
rect 45554 16192 45560 16204
rect 45612 16192 45618 16244
rect 44146 16167 44204 16173
rect 44146 16164 44158 16167
rect 43456 16136 44158 16164
rect 44146 16133 44158 16136
rect 44192 16133 44204 16167
rect 44146 16127 44204 16133
rect 25593 16099 25651 16105
rect 25593 16096 25605 16099
rect 24820 16068 25605 16096
rect 24820 16056 24826 16068
rect 25593 16065 25605 16068
rect 25639 16065 25651 16099
rect 25593 16059 25651 16065
rect 27341 16099 27399 16105
rect 27341 16065 27353 16099
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 28169 16099 28227 16105
rect 28169 16065 28181 16099
rect 28215 16065 28227 16099
rect 29822 16096 29828 16108
rect 29783 16068 29828 16096
rect 28169 16059 28227 16065
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 5442 15920 5448 15972
rect 5500 15960 5506 15972
rect 6365 15963 6423 15969
rect 6365 15960 6377 15963
rect 5500 15932 6377 15960
rect 5500 15920 5506 15932
rect 6365 15929 6377 15932
rect 6411 15929 6423 15963
rect 6365 15923 6423 15929
rect 6840 15892 6868 15991
rect 6914 15988 6920 16040
rect 6972 16028 6978 16040
rect 7834 16028 7840 16040
rect 6972 16000 7017 16028
rect 7795 16000 7840 16028
rect 6972 15988 6978 16000
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 10502 16028 10508 16040
rect 10463 16000 10508 16028
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 15930 16028 15936 16040
rect 15891 16000 15936 16028
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 18138 16028 18144 16040
rect 18099 16000 18144 16028
rect 18138 15988 18144 16000
rect 18196 15988 18202 16040
rect 22646 15988 22652 16040
rect 22704 16028 22710 16040
rect 23477 16031 23535 16037
rect 23477 16028 23489 16031
rect 22704 16000 23489 16028
rect 22704 15988 22710 16000
rect 23477 15997 23489 16000
rect 23523 16028 23535 16031
rect 24489 16031 24547 16037
rect 24489 16028 24501 16031
rect 23523 16000 24501 16028
rect 23523 15997 23535 16000
rect 23477 15991 23535 15997
rect 24489 15997 24501 16000
rect 24535 15997 24547 16031
rect 27062 16028 27068 16040
rect 27023 16000 27068 16028
rect 24489 15991 24547 15997
rect 27062 15988 27068 16000
rect 27120 15988 27126 16040
rect 27356 16028 27384 16059
rect 29822 16056 29828 16068
rect 29880 16056 29886 16108
rect 33781 16099 33839 16105
rect 33781 16065 33793 16099
rect 33827 16096 33839 16099
rect 34146 16096 34152 16108
rect 33827 16068 34152 16096
rect 33827 16065 33839 16068
rect 33781 16059 33839 16065
rect 34146 16056 34152 16068
rect 34204 16056 34210 16108
rect 34790 16096 34796 16108
rect 34751 16068 34796 16096
rect 34790 16056 34796 16068
rect 34848 16056 34854 16108
rect 43257 16099 43315 16105
rect 43257 16065 43269 16099
rect 43303 16096 43315 16099
rect 43714 16096 43720 16108
rect 43303 16068 43720 16096
rect 43303 16065 43315 16068
rect 43257 16059 43315 16065
rect 43714 16056 43720 16068
rect 43772 16056 43778 16108
rect 29840 16028 29868 16056
rect 27356 16000 29868 16028
rect 30101 16031 30159 16037
rect 30101 15997 30113 16031
rect 30147 15997 30159 16031
rect 32766 16028 32772 16040
rect 32727 16000 32772 16028
rect 30101 15991 30159 15997
rect 12158 15920 12164 15972
rect 12216 15960 12222 15972
rect 24670 15960 24676 15972
rect 12216 15932 24676 15960
rect 12216 15920 12222 15932
rect 24670 15920 24676 15932
rect 24728 15920 24734 15972
rect 25133 15963 25191 15969
rect 25133 15929 25145 15963
rect 25179 15960 25191 15963
rect 28074 15960 28080 15972
rect 25179 15932 28080 15960
rect 25179 15929 25191 15932
rect 25133 15923 25191 15929
rect 28074 15920 28080 15932
rect 28132 15920 28138 15972
rect 30116 15960 30144 15991
rect 32766 15988 32772 16000
rect 32824 15988 32830 16040
rect 32861 16031 32919 16037
rect 32861 15997 32873 16031
rect 32907 15997 32919 16031
rect 32861 15991 32919 15997
rect 32674 15960 32680 15972
rect 30116 15932 32680 15960
rect 32674 15920 32680 15932
rect 32732 15960 32738 15972
rect 32876 15960 32904 15991
rect 34606 15988 34612 16040
rect 34664 16028 34670 16040
rect 34701 16031 34759 16037
rect 34701 16028 34713 16031
rect 34664 16000 34713 16028
rect 34664 15988 34670 16000
rect 34701 15997 34713 16000
rect 34747 15997 34759 16031
rect 34701 15991 34759 15997
rect 42426 15988 42432 16040
rect 42484 16028 42490 16040
rect 43901 16031 43959 16037
rect 43901 16028 43913 16031
rect 42484 16000 43913 16028
rect 42484 15988 42490 16000
rect 43901 15997 43913 16000
rect 43947 15997 43959 16031
rect 43901 15991 43959 15997
rect 32732 15932 32904 15960
rect 32732 15920 32738 15932
rect 8570 15892 8576 15904
rect 6840 15864 8576 15892
rect 8570 15852 8576 15864
rect 8628 15852 8634 15904
rect 14090 15852 14096 15904
rect 14148 15892 14154 15904
rect 14185 15895 14243 15901
rect 14185 15892 14197 15895
rect 14148 15864 14197 15892
rect 14148 15852 14154 15864
rect 14185 15861 14197 15864
rect 14231 15861 14243 15895
rect 15286 15892 15292 15904
rect 15247 15864 15292 15892
rect 14185 15855 14243 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 28258 15892 28264 15904
rect 28219 15864 28264 15892
rect 28258 15852 28264 15864
rect 28316 15852 28322 15904
rect 28902 15892 28908 15904
rect 28863 15864 28908 15892
rect 28902 15852 28908 15864
rect 28960 15852 28966 15904
rect 34422 15892 34428 15904
rect 34383 15864 34428 15892
rect 34422 15852 34428 15864
rect 34480 15852 34486 15904
rect 1104 15802 68816 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 65654 15802
rect 65706 15750 65718 15802
rect 65770 15750 65782 15802
rect 65834 15750 65846 15802
rect 65898 15750 65910 15802
rect 65962 15750 68816 15802
rect 1104 15728 68816 15750
rect 5166 15688 5172 15700
rect 5127 15660 5172 15688
rect 5166 15648 5172 15660
rect 5224 15648 5230 15700
rect 6454 15648 6460 15700
rect 6512 15688 6518 15700
rect 6512 15660 6868 15688
rect 6512 15648 6518 15660
rect 6840 15632 6868 15660
rect 7006 15648 7012 15700
rect 7064 15688 7070 15700
rect 7193 15691 7251 15697
rect 7193 15688 7205 15691
rect 7064 15660 7205 15688
rect 7064 15648 7070 15660
rect 7193 15657 7205 15660
rect 7239 15688 7251 15691
rect 7742 15688 7748 15700
rect 7239 15660 7748 15688
rect 7239 15657 7251 15660
rect 7193 15651 7251 15657
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 15746 15688 15752 15700
rect 14752 15660 15752 15688
rect 6822 15580 6828 15632
rect 6880 15620 6886 15632
rect 9493 15623 9551 15629
rect 9493 15620 9505 15623
rect 6880 15592 9505 15620
rect 6880 15580 6886 15592
rect 9493 15589 9505 15592
rect 9539 15589 9551 15623
rect 9493 15583 9551 15589
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 5813 15555 5871 15561
rect 5813 15552 5825 15555
rect 4672 15524 5825 15552
rect 4672 15512 4678 15524
rect 5813 15521 5825 15524
rect 5859 15521 5871 15555
rect 5813 15515 5871 15521
rect 5353 15487 5411 15493
rect 5353 15453 5365 15487
rect 5399 15484 5411 15487
rect 5442 15484 5448 15496
rect 5399 15456 5448 15484
rect 5399 15453 5411 15456
rect 5353 15447 5411 15453
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 5828 15484 5856 15515
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 14752 15561 14780 15660
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 16669 15691 16727 15697
rect 16669 15657 16681 15691
rect 16715 15688 16727 15691
rect 16850 15688 16856 15700
rect 16715 15660 16856 15688
rect 16715 15657 16727 15660
rect 16669 15651 16727 15657
rect 16850 15648 16856 15660
rect 16908 15648 16914 15700
rect 21821 15691 21879 15697
rect 21821 15657 21833 15691
rect 21867 15688 21879 15691
rect 22186 15688 22192 15700
rect 21867 15660 22192 15688
rect 21867 15657 21879 15660
rect 21821 15651 21879 15657
rect 22186 15648 22192 15660
rect 22244 15648 22250 15700
rect 24026 15688 24032 15700
rect 23492 15660 24032 15688
rect 16758 15580 16764 15632
rect 16816 15620 16822 15632
rect 23492 15620 23520 15660
rect 24026 15648 24032 15660
rect 24084 15648 24090 15700
rect 28074 15648 28080 15700
rect 28132 15688 28138 15700
rect 28169 15691 28227 15697
rect 28169 15688 28181 15691
rect 28132 15660 28181 15688
rect 28132 15648 28138 15660
rect 28169 15657 28181 15660
rect 28215 15688 28227 15691
rect 28258 15688 28264 15700
rect 28215 15660 28264 15688
rect 28215 15657 28227 15660
rect 28169 15651 28227 15657
rect 28258 15648 28264 15660
rect 28316 15648 28322 15700
rect 28902 15648 28908 15700
rect 28960 15688 28966 15700
rect 38378 15688 38384 15700
rect 28960 15660 38384 15688
rect 28960 15648 28966 15660
rect 38378 15648 38384 15660
rect 38436 15688 38442 15700
rect 39209 15691 39267 15697
rect 39209 15688 39221 15691
rect 38436 15660 39221 15688
rect 38436 15648 38442 15660
rect 39209 15657 39221 15660
rect 39255 15688 39267 15691
rect 40034 15688 40040 15700
rect 39255 15660 40040 15688
rect 39255 15657 39267 15660
rect 39209 15651 39267 15657
rect 40034 15648 40040 15660
rect 40092 15648 40098 15700
rect 41322 15648 41328 15700
rect 41380 15688 41386 15700
rect 42337 15691 42395 15697
rect 41380 15660 42104 15688
rect 41380 15648 41386 15660
rect 16816 15592 23520 15620
rect 16816 15580 16822 15592
rect 23566 15580 23572 15632
rect 23624 15620 23630 15632
rect 28920 15620 28948 15648
rect 23624 15592 28948 15620
rect 40221 15623 40279 15629
rect 23624 15580 23630 15592
rect 7653 15555 7711 15561
rect 7653 15552 7665 15555
rect 7156 15524 7665 15552
rect 7156 15512 7162 15524
rect 7653 15521 7665 15524
rect 7699 15521 7711 15555
rect 7653 15515 7711 15521
rect 10873 15555 10931 15561
rect 10873 15521 10885 15555
rect 10919 15521 10931 15555
rect 10873 15515 10931 15521
rect 14737 15555 14795 15561
rect 14737 15521 14749 15555
rect 14783 15521 14795 15555
rect 17218 15552 17224 15564
rect 17179 15524 17224 15552
rect 14737 15515 14795 15521
rect 8294 15484 8300 15496
rect 5828 15456 8300 15484
rect 8294 15444 8300 15456
rect 8352 15444 8358 15496
rect 10594 15484 10600 15496
rect 10555 15456 10600 15484
rect 10594 15444 10600 15456
rect 10652 15444 10658 15496
rect 6080 15419 6138 15425
rect 6080 15385 6092 15419
rect 6126 15416 6138 15419
rect 6362 15416 6368 15428
rect 6126 15388 6368 15416
rect 6126 15385 6138 15388
rect 6080 15379 6138 15385
rect 6362 15376 6368 15388
rect 6420 15376 6426 15428
rect 7837 15419 7895 15425
rect 7837 15385 7849 15419
rect 7883 15385 7895 15419
rect 7837 15379 7895 15385
rect 7852 15348 7880 15379
rect 9674 15376 9680 15428
rect 9732 15416 9738 15428
rect 10888 15416 10916 15515
rect 17218 15512 17224 15524
rect 17276 15512 17282 15564
rect 26142 15512 26148 15564
rect 26200 15552 26206 15564
rect 28092 15561 28120 15592
rect 40221 15589 40233 15623
rect 40267 15620 40279 15623
rect 40310 15620 40316 15632
rect 40267 15592 40316 15620
rect 40267 15589 40279 15592
rect 40221 15583 40279 15589
rect 40310 15580 40316 15592
rect 40368 15580 40374 15632
rect 41782 15620 41788 15632
rect 41743 15592 41788 15620
rect 41782 15580 41788 15592
rect 41840 15580 41846 15632
rect 42076 15620 42104 15660
rect 42337 15657 42349 15691
rect 42383 15688 42395 15691
rect 42610 15688 42616 15700
rect 42383 15660 42616 15688
rect 42383 15657 42395 15660
rect 42337 15651 42395 15657
rect 42610 15648 42616 15660
rect 42668 15648 42674 15700
rect 42981 15623 43039 15629
rect 42981 15620 42993 15623
rect 42076 15592 42993 15620
rect 42981 15589 42993 15592
rect 43027 15589 43039 15623
rect 42981 15583 43039 15589
rect 44453 15623 44511 15629
rect 44453 15589 44465 15623
rect 44499 15620 44511 15623
rect 45370 15620 45376 15632
rect 44499 15592 45376 15620
rect 44499 15589 44511 15592
rect 44453 15583 44511 15589
rect 45370 15580 45376 15592
rect 45428 15580 45434 15632
rect 26697 15555 26755 15561
rect 26697 15552 26709 15555
rect 26200 15524 26709 15552
rect 26200 15512 26206 15524
rect 26697 15521 26709 15524
rect 26743 15521 26755 15555
rect 26697 15515 26755 15521
rect 28077 15555 28135 15561
rect 28077 15521 28089 15555
rect 28123 15521 28135 15555
rect 28077 15515 28135 15521
rect 28166 15512 28172 15564
rect 28224 15552 28230 15564
rect 29825 15555 29883 15561
rect 29825 15552 29837 15555
rect 28224 15524 29837 15552
rect 28224 15512 28230 15524
rect 29825 15521 29837 15524
rect 29871 15521 29883 15555
rect 29825 15515 29883 15521
rect 41417 15555 41475 15561
rect 41417 15521 41429 15555
rect 41463 15552 41475 15555
rect 41598 15552 41604 15564
rect 41463 15524 41604 15552
rect 41463 15521 41475 15524
rect 41417 15515 41475 15521
rect 41598 15512 41604 15524
rect 41656 15512 41662 15564
rect 43993 15555 44051 15561
rect 43993 15552 44005 15555
rect 43272 15524 44005 15552
rect 43272 15496 43300 15524
rect 43993 15521 44005 15524
rect 44039 15521 44051 15555
rect 43993 15515 44051 15521
rect 11974 15444 11980 15496
rect 12032 15484 12038 15496
rect 12805 15487 12863 15493
rect 12805 15484 12817 15487
rect 12032 15456 12817 15484
rect 12032 15444 12038 15456
rect 12805 15453 12817 15456
rect 12851 15453 12863 15487
rect 12805 15447 12863 15453
rect 14093 15487 14151 15493
rect 14093 15453 14105 15487
rect 14139 15484 14151 15487
rect 15286 15484 15292 15496
rect 14139 15456 15292 15484
rect 14139 15453 14151 15456
rect 14093 15447 14151 15453
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 17034 15484 17040 15496
rect 16995 15456 17040 15484
rect 17034 15444 17040 15456
rect 17092 15444 17098 15496
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 19978 15484 19984 15496
rect 19392 15456 19984 15484
rect 19392 15444 19398 15456
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 22278 15484 22284 15496
rect 22239 15456 22284 15484
rect 22278 15444 22284 15456
rect 22336 15444 22342 15496
rect 22462 15484 22468 15496
rect 22423 15456 22468 15484
rect 22462 15444 22468 15456
rect 22520 15444 22526 15496
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15484 23719 15487
rect 23750 15484 23756 15496
rect 23707 15456 23756 15484
rect 23707 15453 23719 15456
rect 23661 15447 23719 15453
rect 23750 15444 23756 15456
rect 23808 15444 23814 15496
rect 26789 15487 26847 15493
rect 26789 15484 26801 15487
rect 26068 15456 26801 15484
rect 12526 15416 12532 15428
rect 12584 15425 12590 15428
rect 9732 15388 9777 15416
rect 9876 15388 12434 15416
rect 12496 15388 12532 15416
rect 9732 15376 9738 15388
rect 8202 15348 8208 15360
rect 7852 15320 8208 15348
rect 8202 15308 8208 15320
rect 8260 15348 8266 15360
rect 9876 15348 9904 15388
rect 8260 15320 9904 15348
rect 8260 15308 8266 15320
rect 10134 15308 10140 15360
rect 10192 15348 10198 15360
rect 10229 15351 10287 15357
rect 10229 15348 10241 15351
rect 10192 15320 10241 15348
rect 10192 15308 10198 15320
rect 10229 15317 10241 15320
rect 10275 15317 10287 15351
rect 10229 15311 10287 15317
rect 10689 15351 10747 15357
rect 10689 15317 10701 15351
rect 10735 15348 10747 15351
rect 11054 15348 11060 15360
rect 10735 15320 11060 15348
rect 10735 15317 10747 15320
rect 10689 15311 10747 15317
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11422 15348 11428 15360
rect 11383 15320 11428 15348
rect 11422 15308 11428 15320
rect 11480 15308 11486 15360
rect 12406 15348 12434 15388
rect 12526 15376 12532 15388
rect 12584 15379 12596 15425
rect 14982 15419 15040 15425
rect 14982 15416 14994 15419
rect 14292 15388 14994 15416
rect 12584 15376 12590 15379
rect 13722 15348 13728 15360
rect 12406 15320 13728 15348
rect 13722 15308 13728 15320
rect 13780 15308 13786 15360
rect 14292 15357 14320 15388
rect 14982 15385 14994 15388
rect 15028 15385 15040 15419
rect 14982 15379 15040 15385
rect 16574 15376 16580 15428
rect 16632 15416 16638 15428
rect 17129 15419 17187 15425
rect 17129 15416 17141 15419
rect 16632 15388 17141 15416
rect 16632 15376 16638 15388
rect 17129 15385 17141 15388
rect 17175 15416 17187 15419
rect 17865 15419 17923 15425
rect 17865 15416 17877 15419
rect 17175 15388 17877 15416
rect 17175 15385 17187 15388
rect 17129 15379 17187 15385
rect 17865 15385 17877 15388
rect 17911 15385 17923 15419
rect 17865 15379 17923 15385
rect 23382 15376 23388 15428
rect 23440 15416 23446 15428
rect 24673 15419 24731 15425
rect 24673 15416 24685 15419
rect 23440 15388 24685 15416
rect 23440 15376 23446 15388
rect 24673 15385 24685 15388
rect 24719 15416 24731 15419
rect 24854 15416 24860 15428
rect 24719 15388 24860 15416
rect 24719 15385 24731 15388
rect 24673 15379 24731 15385
rect 24854 15376 24860 15388
rect 24912 15376 24918 15428
rect 14277 15351 14335 15357
rect 14277 15317 14289 15351
rect 14323 15317 14335 15351
rect 14277 15311 14335 15317
rect 16117 15351 16175 15357
rect 16117 15317 16129 15351
rect 16163 15348 16175 15351
rect 16942 15348 16948 15360
rect 16163 15320 16948 15348
rect 16163 15317 16175 15320
rect 16117 15311 16175 15317
rect 16942 15308 16948 15320
rect 17000 15308 17006 15360
rect 19334 15348 19340 15360
rect 19247 15320 19340 15348
rect 19334 15308 19340 15320
rect 19392 15348 19398 15360
rect 20622 15348 20628 15360
rect 19392 15320 20628 15348
rect 19392 15308 19398 15320
rect 20622 15308 20628 15320
rect 20680 15308 20686 15360
rect 22370 15348 22376 15360
rect 22331 15320 22376 15348
rect 22370 15308 22376 15320
rect 22428 15308 22434 15360
rect 22922 15348 22928 15360
rect 22883 15320 22928 15348
rect 22922 15308 22928 15320
rect 22980 15308 22986 15360
rect 23658 15308 23664 15360
rect 23716 15348 23722 15360
rect 23753 15351 23811 15357
rect 23753 15348 23765 15351
rect 23716 15320 23765 15348
rect 23716 15308 23722 15320
rect 23753 15317 23765 15320
rect 23799 15317 23811 15351
rect 23753 15311 23811 15317
rect 25682 15308 25688 15360
rect 25740 15348 25746 15360
rect 26068 15357 26096 15456
rect 26789 15453 26801 15456
rect 26835 15453 26847 15487
rect 26789 15447 26847 15453
rect 28353 15487 28411 15493
rect 28353 15453 28365 15487
rect 28399 15484 28411 15487
rect 29362 15484 29368 15496
rect 28399 15456 29368 15484
rect 28399 15453 28411 15456
rect 28353 15447 28411 15453
rect 29362 15444 29368 15456
rect 29420 15444 29426 15496
rect 29914 15484 29920 15496
rect 29875 15456 29920 15484
rect 29914 15444 29920 15456
rect 29972 15444 29978 15496
rect 32125 15487 32183 15493
rect 32125 15453 32137 15487
rect 32171 15484 32183 15487
rect 32858 15484 32864 15496
rect 32171 15456 32864 15484
rect 32171 15453 32183 15456
rect 32125 15447 32183 15453
rect 32858 15444 32864 15456
rect 32916 15444 32922 15496
rect 41495 15487 41553 15493
rect 41495 15484 41507 15487
rect 41386 15456 41507 15484
rect 32392 15419 32450 15425
rect 32392 15385 32404 15419
rect 32438 15416 32450 15419
rect 32490 15416 32496 15428
rect 32438 15388 32496 15416
rect 32438 15385 32450 15388
rect 32392 15379 32450 15385
rect 32490 15376 32496 15388
rect 32548 15376 32554 15428
rect 39666 15376 39672 15428
rect 39724 15416 39730 15428
rect 39853 15419 39911 15425
rect 39853 15416 39865 15419
rect 39724 15388 39865 15416
rect 39724 15376 39730 15388
rect 39853 15385 39865 15388
rect 39899 15416 39911 15419
rect 41386 15416 41414 15456
rect 41495 15453 41507 15456
rect 41541 15453 41553 15487
rect 41495 15447 41553 15453
rect 42981 15487 43039 15493
rect 42981 15453 42993 15487
rect 43027 15484 43039 15487
rect 43162 15484 43168 15496
rect 43027 15456 43168 15484
rect 43027 15453 43039 15456
rect 42981 15447 43039 15453
rect 43162 15444 43168 15456
rect 43220 15444 43226 15496
rect 43254 15444 43260 15496
rect 43312 15484 43318 15496
rect 44085 15487 44143 15493
rect 44085 15484 44097 15487
rect 43312 15456 43357 15484
rect 43548 15456 44097 15484
rect 43312 15444 43318 15456
rect 39899 15388 41414 15416
rect 39899 15385 39911 15388
rect 39853 15379 39911 15385
rect 26053 15351 26111 15357
rect 26053 15348 26065 15351
rect 25740 15320 26065 15348
rect 25740 15308 25746 15320
rect 26053 15317 26065 15320
rect 26099 15317 26111 15351
rect 26053 15311 26111 15317
rect 27157 15351 27215 15357
rect 27157 15317 27169 15351
rect 27203 15348 27215 15351
rect 28166 15348 28172 15360
rect 27203 15320 28172 15348
rect 27203 15317 27215 15320
rect 27157 15311 27215 15317
rect 28166 15308 28172 15320
rect 28224 15308 28230 15360
rect 28534 15348 28540 15360
rect 28495 15320 28540 15348
rect 28534 15308 28540 15320
rect 28592 15308 28598 15360
rect 29546 15348 29552 15360
rect 29507 15320 29552 15348
rect 29546 15308 29552 15320
rect 29604 15308 29610 15360
rect 32766 15308 32772 15360
rect 32824 15348 32830 15360
rect 33505 15351 33563 15357
rect 33505 15348 33517 15351
rect 32824 15320 33517 15348
rect 32824 15308 32830 15320
rect 33505 15317 33517 15320
rect 33551 15317 33563 15351
rect 33505 15311 33563 15317
rect 40313 15351 40371 15357
rect 40313 15317 40325 15351
rect 40359 15348 40371 15351
rect 40402 15348 40408 15360
rect 40359 15320 40408 15348
rect 40359 15317 40371 15320
rect 40313 15311 40371 15317
rect 40402 15308 40408 15320
rect 40460 15308 40466 15360
rect 41386 15348 41414 15388
rect 43548 15360 43576 15456
rect 44085 15453 44097 15456
rect 44131 15453 44143 15487
rect 44085 15447 44143 15453
rect 41506 15348 41512 15360
rect 41386 15320 41512 15348
rect 41506 15308 41512 15320
rect 41564 15308 41570 15360
rect 43165 15351 43223 15357
rect 43165 15317 43177 15351
rect 43211 15348 43223 15351
rect 43530 15348 43536 15360
rect 43211 15320 43536 15348
rect 43211 15317 43223 15320
rect 43165 15311 43223 15317
rect 43530 15308 43536 15320
rect 43588 15308 43594 15360
rect 1104 15258 68816 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 68816 15258
rect 1104 15184 68816 15206
rect 7006 15144 7012 15156
rect 6967 15116 7012 15144
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 10594 15144 10600 15156
rect 10555 15116 10600 15144
rect 10594 15104 10600 15116
rect 10652 15104 10658 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11609 15147 11667 15153
rect 11609 15144 11621 15147
rect 11112 15116 11621 15144
rect 11112 15104 11118 15116
rect 11609 15113 11621 15116
rect 11655 15144 11667 15147
rect 12342 15144 12348 15156
rect 11655 15116 12348 15144
rect 11655 15113 11667 15116
rect 11609 15107 11667 15113
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 12526 15144 12532 15156
rect 12487 15116 12532 15144
rect 12526 15104 12532 15116
rect 12584 15104 12590 15156
rect 13173 15147 13231 15153
rect 13173 15113 13185 15147
rect 13219 15113 13231 15147
rect 13173 15107 13231 15113
rect 20533 15147 20591 15153
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 20622 15144 20628 15156
rect 20579 15116 20628 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 8294 14968 8300 15020
rect 8352 15008 8358 15020
rect 9217 15011 9275 15017
rect 9217 15008 9229 15011
rect 8352 14980 9229 15008
rect 8352 14968 8358 14980
rect 9217 14977 9229 14980
rect 9263 14977 9275 15011
rect 9217 14971 9275 14977
rect 9484 15011 9542 15017
rect 9484 14977 9496 15011
rect 9530 15008 9542 15011
rect 9950 15008 9956 15020
rect 9530 14980 9956 15008
rect 9530 14977 9542 14980
rect 9484 14971 9542 14977
rect 9950 14968 9956 14980
rect 10008 14968 10014 15020
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 15008 12403 15011
rect 13188 15008 13216 15107
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 22189 15147 22247 15153
rect 22189 15113 22201 15147
rect 22235 15144 22247 15147
rect 22278 15144 22284 15156
rect 22235 15116 22284 15144
rect 22235 15113 22247 15116
rect 22189 15107 22247 15113
rect 22278 15104 22284 15116
rect 22336 15104 22342 15156
rect 24397 15147 24455 15153
rect 24397 15113 24409 15147
rect 24443 15144 24455 15147
rect 24857 15147 24915 15153
rect 24857 15144 24869 15147
rect 24443 15116 24869 15144
rect 24443 15113 24455 15116
rect 24397 15107 24455 15113
rect 24857 15113 24869 15116
rect 24903 15144 24915 15147
rect 26234 15144 26240 15156
rect 24903 15116 26240 15144
rect 24903 15113 24915 15116
rect 24857 15107 24915 15113
rect 26234 15104 26240 15116
rect 26292 15104 26298 15156
rect 27062 15104 27068 15156
rect 27120 15144 27126 15156
rect 27246 15144 27252 15156
rect 27120 15116 27252 15144
rect 27120 15104 27126 15116
rect 27246 15104 27252 15116
rect 27304 15104 27310 15156
rect 27338 15104 27344 15156
rect 27396 15144 27402 15156
rect 27893 15147 27951 15153
rect 27893 15144 27905 15147
rect 27396 15116 27905 15144
rect 27396 15104 27402 15116
rect 27893 15113 27905 15116
rect 27939 15113 27951 15147
rect 27893 15107 27951 15113
rect 34149 15147 34207 15153
rect 34149 15113 34161 15147
rect 34195 15144 34207 15147
rect 34514 15144 34520 15156
rect 34195 15116 34520 15144
rect 34195 15113 34207 15116
rect 34149 15107 34207 15113
rect 13446 15036 13452 15088
rect 13504 15076 13510 15088
rect 13633 15079 13691 15085
rect 13633 15076 13645 15079
rect 13504 15048 13645 15076
rect 13504 15036 13510 15048
rect 13633 15045 13645 15048
rect 13679 15076 13691 15079
rect 13679 15048 15516 15076
rect 13679 15045 13691 15048
rect 13633 15039 13691 15045
rect 15488 15020 15516 15048
rect 15930 15036 15936 15088
rect 15988 15076 15994 15088
rect 17037 15079 17095 15085
rect 17037 15076 17049 15079
rect 15988 15048 17049 15076
rect 15988 15036 15994 15048
rect 17037 15045 17049 15048
rect 17083 15045 17095 15079
rect 17037 15039 17095 15045
rect 18248 15048 21312 15076
rect 12391 14980 13216 15008
rect 13541 15011 13599 15017
rect 12391 14977 12403 14980
rect 12345 14971 12403 14977
rect 13541 14977 13553 15011
rect 13587 14977 13599 15011
rect 13541 14971 13599 14977
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14909 7159 14943
rect 7101 14903 7159 14909
rect 7285 14943 7343 14949
rect 7285 14909 7297 14943
rect 7331 14940 7343 14943
rect 7374 14940 7380 14952
rect 7331 14912 7380 14940
rect 7331 14909 7343 14912
rect 7285 14903 7343 14909
rect 7116 14872 7144 14903
rect 7374 14900 7380 14912
rect 7432 14900 7438 14952
rect 11422 14900 11428 14952
rect 11480 14940 11486 14952
rect 13556 14940 13584 14971
rect 14090 14968 14096 15020
rect 14148 15008 14154 15020
rect 14369 15011 14427 15017
rect 14369 15008 14381 15011
rect 14148 14980 14381 15008
rect 14148 14968 14154 14980
rect 14369 14977 14381 14980
rect 14415 14977 14427 15011
rect 14369 14971 14427 14977
rect 14458 14968 14464 15020
rect 14516 15008 14522 15020
rect 14553 15011 14611 15017
rect 14553 15008 14565 15011
rect 14516 14980 14565 15008
rect 14516 14968 14522 14980
rect 14553 14977 14565 14980
rect 14599 14977 14611 15011
rect 15470 15008 15476 15020
rect 15431 14980 15476 15008
rect 14553 14971 14611 14977
rect 15470 14968 15476 14980
rect 15528 14968 15534 15020
rect 17218 15008 17224 15020
rect 17179 14980 17224 15008
rect 17218 14968 17224 14980
rect 17276 14968 17282 15020
rect 11480 14912 13584 14940
rect 13817 14943 13875 14949
rect 11480 14900 11486 14912
rect 13817 14909 13829 14943
rect 13863 14940 13875 14943
rect 14734 14940 14740 14952
rect 13863 14912 14740 14940
rect 13863 14909 13875 14912
rect 13817 14903 13875 14909
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 18138 14940 18144 14952
rect 18051 14912 18144 14940
rect 18138 14900 18144 14912
rect 18196 14940 18202 14952
rect 18248 14940 18276 15048
rect 21284 15020 21312 15048
rect 21634 15036 21640 15088
rect 21692 15076 21698 15088
rect 21821 15079 21879 15085
rect 21821 15076 21833 15079
rect 21692 15048 21833 15076
rect 21692 15036 21698 15048
rect 21821 15045 21833 15048
rect 21867 15045 21879 15079
rect 21821 15039 21879 15045
rect 22002 15036 22008 15088
rect 22060 15085 22066 15088
rect 22060 15079 22079 15085
rect 22067 15045 22079 15079
rect 22060 15039 22079 15045
rect 22060 15036 22066 15039
rect 22370 15036 22376 15088
rect 22428 15076 22434 15088
rect 22925 15079 22983 15085
rect 22925 15076 22937 15079
rect 22428 15048 22937 15076
rect 22428 15036 22434 15048
rect 22925 15045 22937 15048
rect 22971 15045 22983 15079
rect 22925 15039 22983 15045
rect 23658 15036 23664 15088
rect 23716 15036 23722 15088
rect 27522 15076 27528 15088
rect 26252 15048 27528 15076
rect 18414 15017 18420 15020
rect 18408 14971 18420 15017
rect 18472 15008 18478 15020
rect 18472 14980 18508 15008
rect 18414 14968 18420 14971
rect 18472 14968 18478 14980
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 20257 15011 20315 15017
rect 20257 15008 20269 15011
rect 19484 14980 20269 15008
rect 19484 14968 19490 14980
rect 20257 14977 20269 14980
rect 20303 15008 20315 15011
rect 20530 15008 20536 15020
rect 20303 14980 20536 15008
rect 20303 14977 20315 14980
rect 20257 14971 20315 14977
rect 20530 14968 20536 14980
rect 20588 15008 20594 15020
rect 21085 15011 21143 15017
rect 21085 15008 21097 15011
rect 20588 14980 21097 15008
rect 20588 14968 20594 14980
rect 21085 14977 21097 14980
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 21266 14968 21272 15020
rect 21324 15008 21330 15020
rect 22649 15011 22707 15017
rect 22649 15008 22661 15011
rect 21324 14980 22661 15008
rect 21324 14968 21330 14980
rect 22649 14977 22661 14980
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 24210 14968 24216 15020
rect 24268 15008 24274 15020
rect 26252 15017 26280 15048
rect 27522 15036 27528 15048
rect 27580 15076 27586 15088
rect 32858 15076 32864 15088
rect 27580 15048 32864 15076
rect 27580 15036 27586 15048
rect 32858 15036 32864 15048
rect 32916 15036 32922 15088
rect 34164 15076 34192 15107
rect 34514 15104 34520 15116
rect 34572 15104 34578 15156
rect 38838 15144 38844 15156
rect 38799 15116 38844 15144
rect 38838 15104 38844 15116
rect 38896 15104 38902 15156
rect 39758 15144 39764 15156
rect 39719 15116 39764 15144
rect 39758 15104 39764 15116
rect 39816 15104 39822 15156
rect 40402 15144 40408 15156
rect 40144 15116 40408 15144
rect 33612 15048 34192 15076
rect 34333 15079 34391 15085
rect 25970 15011 26028 15017
rect 25970 15008 25982 15011
rect 24268 14980 25982 15008
rect 24268 14968 24274 14980
rect 25970 14977 25982 14980
rect 26016 14977 26028 15011
rect 25970 14971 26028 14977
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 26786 14968 26792 15020
rect 26844 15008 26850 15020
rect 28074 15017 28080 15020
rect 27157 15011 27215 15017
rect 27157 15008 27169 15011
rect 26844 14980 27169 15008
rect 26844 14968 26850 14980
rect 27157 14977 27169 14980
rect 27203 14977 27215 15011
rect 28072 15008 28080 15017
rect 28035 14980 28080 15008
rect 27157 14971 27215 14977
rect 28072 14971 28080 14980
rect 28074 14968 28080 14971
rect 28132 14968 28138 15020
rect 28169 15011 28227 15017
rect 28169 14977 28181 15011
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 18196 14912 18276 14940
rect 18196 14900 18202 14912
rect 26510 14900 26516 14952
rect 26568 14940 26574 14952
rect 28184 14940 28212 14971
rect 28258 14968 28264 15020
rect 28316 15008 28322 15020
rect 28444 15011 28502 15017
rect 28316 14980 28361 15008
rect 28316 14968 28322 14980
rect 28444 14977 28456 15011
rect 28490 14977 28502 15011
rect 28444 14971 28502 14977
rect 26568 14912 28212 14940
rect 26568 14900 26574 14912
rect 7116 14844 7972 14872
rect 6546 14764 6552 14816
rect 6604 14804 6610 14816
rect 7944 14813 7972 14844
rect 12434 14832 12440 14884
rect 12492 14872 12498 14884
rect 14369 14875 14427 14881
rect 14369 14872 14381 14875
rect 12492 14844 14381 14872
rect 12492 14832 12498 14844
rect 14369 14841 14381 14844
rect 14415 14841 14427 14875
rect 28460 14872 28488 14971
rect 28534 14968 28540 15020
rect 28592 15008 28598 15020
rect 29454 15008 29460 15020
rect 28592 14980 28637 15008
rect 29415 14980 29460 15008
rect 28592 14968 28598 14980
rect 29454 14968 29460 14980
rect 29512 14968 29518 15020
rect 30098 14968 30104 15020
rect 30156 15008 30162 15020
rect 30469 15011 30527 15017
rect 30469 15008 30481 15011
rect 30156 14980 30481 15008
rect 30156 14968 30162 14980
rect 30469 14977 30481 14980
rect 30515 14977 30527 15011
rect 30469 14971 30527 14977
rect 32306 14968 32312 15020
rect 32364 15008 32370 15020
rect 32585 15011 32643 15017
rect 32585 15008 32597 15011
rect 32364 14980 32597 15008
rect 32364 14968 32370 14980
rect 32585 14977 32597 14980
rect 32631 14977 32643 15011
rect 32585 14971 32643 14977
rect 32769 15011 32827 15017
rect 32769 14977 32781 15011
rect 32815 14977 32827 15011
rect 32769 14971 32827 14977
rect 33137 15011 33195 15017
rect 33137 14977 33149 15011
rect 33183 14977 33195 15011
rect 33137 14971 33195 14977
rect 29546 14940 29552 14952
rect 29507 14912 29552 14940
rect 29546 14900 29552 14912
rect 29604 14900 29610 14952
rect 30558 14940 30564 14952
rect 29656 14912 30564 14940
rect 29656 14872 29684 14912
rect 30558 14900 30564 14912
rect 30616 14940 30622 14952
rect 31478 14940 31484 14952
rect 30616 14912 31484 14940
rect 30616 14900 30622 14912
rect 31478 14900 31484 14912
rect 31536 14900 31542 14952
rect 31846 14900 31852 14952
rect 31904 14940 31910 14952
rect 32677 14943 32735 14949
rect 32677 14940 32689 14943
rect 31904 14912 32689 14940
rect 31904 14900 31910 14912
rect 32677 14909 32689 14912
rect 32723 14909 32735 14943
rect 32677 14903 32735 14909
rect 28460 14844 29684 14872
rect 29825 14875 29883 14881
rect 14369 14835 14427 14841
rect 29825 14841 29837 14875
rect 29871 14872 29883 14875
rect 32784 14872 32812 14971
rect 29871 14844 32812 14872
rect 33152 14872 33180 14971
rect 33226 14968 33232 15020
rect 33284 15008 33290 15020
rect 33612 15017 33640 15048
rect 34333 15045 34345 15079
rect 34379 15076 34391 15079
rect 34422 15076 34428 15088
rect 34379 15048 34428 15076
rect 34379 15045 34391 15048
rect 34333 15039 34391 15045
rect 34422 15036 34428 15048
rect 34480 15036 34486 15088
rect 40034 15076 40040 15088
rect 39995 15048 40040 15076
rect 40034 15036 40040 15048
rect 40092 15036 40098 15088
rect 40144 15085 40172 15116
rect 40402 15104 40408 15116
rect 40460 15104 40466 15156
rect 40865 15147 40923 15153
rect 40865 15113 40877 15147
rect 40911 15144 40923 15147
rect 41046 15144 41052 15156
rect 40911 15116 41052 15144
rect 40911 15113 40923 15116
rect 40865 15107 40923 15113
rect 41046 15104 41052 15116
rect 41104 15104 41110 15156
rect 40129 15079 40187 15085
rect 40129 15045 40141 15079
rect 40175 15045 40187 15079
rect 41598 15076 41604 15088
rect 40129 15039 40187 15045
rect 40328 15048 41604 15076
rect 33597 15011 33655 15017
rect 33284 14980 33329 15008
rect 33284 14968 33290 14980
rect 33597 14977 33609 15011
rect 33643 14977 33655 15011
rect 33597 14971 33655 14977
rect 34057 15011 34115 15017
rect 34057 14977 34069 15011
rect 34103 14977 34115 15011
rect 34057 14971 34115 14977
rect 33244 14940 33272 14968
rect 34072 14940 34100 14971
rect 37182 14968 37188 15020
rect 37240 15008 37246 15020
rect 37240 14980 38608 15008
rect 37240 14968 37246 14980
rect 37274 14940 37280 14952
rect 33244 14912 34100 14940
rect 37235 14912 37280 14940
rect 37274 14900 37280 14912
rect 37332 14900 37338 14952
rect 38580 14949 38608 14980
rect 39206 14968 39212 15020
rect 39264 15008 39270 15020
rect 40328 15017 40356 15048
rect 41598 15036 41604 15048
rect 41656 15076 41662 15088
rect 42889 15079 42947 15085
rect 42889 15076 42901 15079
rect 41656 15048 42901 15076
rect 41656 15036 41662 15048
rect 42889 15045 42901 15048
rect 42935 15045 42947 15079
rect 42889 15039 42947 15045
rect 43257 15079 43315 15085
rect 43257 15045 43269 15079
rect 43303 15076 43315 15079
rect 43530 15076 43536 15088
rect 43303 15048 43536 15076
rect 43303 15045 43315 15048
rect 43257 15039 43315 15045
rect 43530 15036 43536 15048
rect 43588 15036 43594 15088
rect 39899 15011 39957 15017
rect 39899 15008 39911 15011
rect 39264 14980 39911 15008
rect 39264 14968 39270 14980
rect 39899 14977 39911 14980
rect 39945 14977 39957 15011
rect 39899 14971 39957 14977
rect 40312 15011 40370 15017
rect 40312 14977 40324 15011
rect 40358 14977 40370 15011
rect 40312 14971 40370 14977
rect 40402 14968 40408 15020
rect 40460 15008 40466 15020
rect 41322 15017 41328 15020
rect 41049 15011 41107 15017
rect 40460 14980 40505 15008
rect 40460 14968 40466 14980
rect 41049 14977 41061 15011
rect 41095 14977 41107 15011
rect 41318 15008 41328 15017
rect 41283 14980 41328 15008
rect 41049 14971 41107 14977
rect 41318 14971 41328 14980
rect 38565 14943 38623 14949
rect 38565 14909 38577 14943
rect 38611 14909 38623 14943
rect 38746 14940 38752 14952
rect 38707 14912 38752 14940
rect 38565 14903 38623 14909
rect 38746 14900 38752 14912
rect 38804 14900 38810 14952
rect 34333 14875 34391 14881
rect 34333 14872 34345 14875
rect 33152 14844 34345 14872
rect 29871 14841 29883 14844
rect 29825 14835 29883 14841
rect 34333 14841 34345 14844
rect 34379 14841 34391 14875
rect 34333 14835 34391 14841
rect 37553 14875 37611 14881
rect 37553 14841 37565 14875
rect 37599 14841 37611 14875
rect 37553 14835 37611 14841
rect 37737 14875 37795 14881
rect 37737 14841 37749 14875
rect 37783 14872 37795 14875
rect 41064 14872 41092 14971
rect 41322 14968 41328 14971
rect 41380 14968 41386 15020
rect 41506 15008 41512 15020
rect 41467 14980 41512 15008
rect 41506 14968 41512 14980
rect 41564 14968 41570 15020
rect 43073 15011 43131 15017
rect 43073 14977 43085 15011
rect 43119 15008 43131 15011
rect 43162 15008 43168 15020
rect 43119 14980 43168 15008
rect 43119 14977 43131 14980
rect 43073 14971 43131 14977
rect 43162 14968 43168 14980
rect 43220 14968 43226 15020
rect 43346 15008 43352 15020
rect 43307 14980 43352 15008
rect 43346 14968 43352 14980
rect 43404 14968 43410 15020
rect 44082 15017 44088 15020
rect 44076 14971 44088 15017
rect 44140 15008 44146 15020
rect 44140 14980 44176 15008
rect 44082 14968 44088 14971
rect 44140 14968 44146 14980
rect 42426 14900 42432 14952
rect 42484 14940 42490 14952
rect 43809 14943 43867 14949
rect 43809 14940 43821 14943
rect 42484 14912 43821 14940
rect 42484 14900 42490 14912
rect 43809 14909 43821 14912
rect 43855 14909 43867 14943
rect 43809 14903 43867 14909
rect 41138 14872 41144 14884
rect 37783 14844 41144 14872
rect 37783 14841 37795 14844
rect 37737 14835 37795 14841
rect 6641 14807 6699 14813
rect 6641 14804 6653 14807
rect 6604 14776 6653 14804
rect 6604 14764 6610 14776
rect 6641 14773 6653 14776
rect 6687 14773 6699 14807
rect 6641 14767 6699 14773
rect 7929 14807 7987 14813
rect 7929 14773 7941 14807
rect 7975 14804 7987 14807
rect 8570 14804 8576 14816
rect 7975 14776 8576 14804
rect 7975 14773 7987 14776
rect 7929 14767 7987 14773
rect 8570 14764 8576 14776
rect 8628 14804 8634 14816
rect 12526 14804 12532 14816
rect 8628 14776 12532 14804
rect 8628 14764 8634 14776
rect 12526 14764 12532 14776
rect 12584 14804 12590 14816
rect 15565 14807 15623 14813
rect 15565 14804 15577 14807
rect 12584 14776 15577 14804
rect 12584 14764 12590 14776
rect 15565 14773 15577 14776
rect 15611 14804 15623 14807
rect 19334 14804 19340 14816
rect 15611 14776 19340 14804
rect 15611 14773 15623 14776
rect 15565 14767 15623 14773
rect 19334 14764 19340 14776
rect 19392 14764 19398 14816
rect 19521 14807 19579 14813
rect 19521 14773 19533 14807
rect 19567 14804 19579 14807
rect 19610 14804 19616 14816
rect 19567 14776 19616 14804
rect 19567 14773 19579 14776
rect 19521 14767 19579 14773
rect 19610 14764 19616 14776
rect 19668 14764 19674 14816
rect 21726 14764 21732 14816
rect 21784 14804 21790 14816
rect 22005 14807 22063 14813
rect 22005 14804 22017 14807
rect 21784 14776 22017 14804
rect 21784 14764 21790 14776
rect 22005 14773 22017 14776
rect 22051 14773 22063 14807
rect 22005 14767 22063 14773
rect 24486 14764 24492 14816
rect 24544 14804 24550 14816
rect 27338 14804 27344 14816
rect 24544 14776 27344 14804
rect 24544 14764 24550 14776
rect 27338 14764 27344 14776
rect 27396 14764 27402 14816
rect 30745 14807 30803 14813
rect 30745 14773 30757 14807
rect 30791 14804 30803 14807
rect 31938 14804 31944 14816
rect 30791 14776 31944 14804
rect 30791 14773 30803 14776
rect 30745 14767 30803 14773
rect 31938 14764 31944 14776
rect 31996 14764 32002 14816
rect 36446 14764 36452 14816
rect 36504 14804 36510 14816
rect 36633 14807 36691 14813
rect 36633 14804 36645 14807
rect 36504 14776 36645 14804
rect 36504 14764 36510 14776
rect 36633 14773 36645 14776
rect 36679 14804 36691 14807
rect 37568 14804 37596 14835
rect 41138 14832 41144 14844
rect 41196 14832 41202 14884
rect 36679 14776 37596 14804
rect 36679 14773 36691 14776
rect 36633 14767 36691 14773
rect 39114 14764 39120 14816
rect 39172 14804 39178 14816
rect 39209 14807 39267 14813
rect 39209 14804 39221 14807
rect 39172 14776 39221 14804
rect 39172 14764 39178 14776
rect 39209 14773 39221 14776
rect 39255 14773 39267 14807
rect 45186 14804 45192 14816
rect 45147 14776 45192 14804
rect 39209 14767 39267 14773
rect 45186 14764 45192 14776
rect 45244 14764 45250 14816
rect 45462 14764 45468 14816
rect 45520 14804 45526 14816
rect 45649 14807 45707 14813
rect 45649 14804 45661 14807
rect 45520 14776 45661 14804
rect 45520 14764 45526 14776
rect 45649 14773 45661 14776
rect 45695 14773 45707 14807
rect 45649 14767 45707 14773
rect 1104 14714 68816 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 65654 14714
rect 65706 14662 65718 14714
rect 65770 14662 65782 14714
rect 65834 14662 65846 14714
rect 65898 14662 65910 14714
rect 65962 14662 68816 14714
rect 1104 14640 68816 14662
rect 6362 14600 6368 14612
rect 6323 14572 6368 14600
rect 6362 14560 6368 14572
rect 6420 14560 6426 14612
rect 9950 14600 9956 14612
rect 9911 14572 9956 14600
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 12437 14603 12495 14609
rect 12437 14569 12449 14603
rect 12483 14600 12495 14603
rect 12526 14600 12532 14612
rect 12483 14572 12532 14600
rect 12483 14569 12495 14572
rect 12437 14563 12495 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13446 14600 13452 14612
rect 13407 14572 13452 14600
rect 13446 14560 13452 14572
rect 13504 14560 13510 14612
rect 17037 14603 17095 14609
rect 17037 14569 17049 14603
rect 17083 14600 17095 14603
rect 18414 14600 18420 14612
rect 17083 14572 18420 14600
rect 17083 14569 17095 14572
rect 17037 14563 17095 14569
rect 18414 14560 18420 14572
rect 18472 14560 18478 14612
rect 20530 14600 20536 14612
rect 20491 14572 20536 14600
rect 20530 14560 20536 14572
rect 20588 14560 20594 14612
rect 22462 14560 22468 14612
rect 22520 14600 22526 14612
rect 22557 14603 22615 14609
rect 22557 14600 22569 14603
rect 22520 14572 22569 14600
rect 22520 14560 22526 14572
rect 22557 14569 22569 14572
rect 22603 14569 22615 14603
rect 22557 14563 22615 14569
rect 23293 14603 23351 14609
rect 23293 14569 23305 14603
rect 23339 14600 23351 14603
rect 24210 14600 24216 14612
rect 23339 14572 24216 14600
rect 23339 14569 23351 14572
rect 23293 14563 23351 14569
rect 24210 14560 24216 14572
rect 24268 14560 24274 14612
rect 26786 14560 26792 14612
rect 26844 14600 26850 14612
rect 26881 14603 26939 14609
rect 26881 14600 26893 14603
rect 26844 14572 26893 14600
rect 26844 14560 26850 14572
rect 26881 14569 26893 14572
rect 26927 14569 26939 14603
rect 26881 14563 26939 14569
rect 28350 14560 28356 14612
rect 28408 14600 28414 14612
rect 28537 14603 28595 14609
rect 28537 14600 28549 14603
rect 28408 14572 28549 14600
rect 28408 14560 28414 14572
rect 28537 14569 28549 14572
rect 28583 14569 28595 14603
rect 28537 14563 28595 14569
rect 29454 14560 29460 14612
rect 29512 14600 29518 14612
rect 29549 14603 29607 14609
rect 29549 14600 29561 14603
rect 29512 14572 29561 14600
rect 29512 14560 29518 14572
rect 29549 14569 29561 14572
rect 29595 14569 29607 14603
rect 32306 14600 32312 14612
rect 32267 14572 32312 14600
rect 29549 14563 29607 14569
rect 32306 14560 32312 14572
rect 32364 14560 32370 14612
rect 37274 14600 37280 14612
rect 37235 14572 37280 14600
rect 37274 14560 37280 14572
rect 37332 14560 37338 14612
rect 39206 14600 39212 14612
rect 39167 14572 39212 14600
rect 39206 14560 39212 14572
rect 39264 14560 39270 14612
rect 40310 14600 40316 14612
rect 40271 14572 40316 14600
rect 40310 14560 40316 14572
rect 40368 14560 40374 14612
rect 40402 14560 40408 14612
rect 40460 14600 40466 14612
rect 41325 14603 41383 14609
rect 41325 14600 41337 14603
rect 40460 14572 41337 14600
rect 40460 14560 40466 14572
rect 41325 14569 41337 14572
rect 41371 14569 41383 14603
rect 41325 14563 41383 14569
rect 16393 14535 16451 14541
rect 16393 14501 16405 14535
rect 16439 14532 16451 14535
rect 17218 14532 17224 14544
rect 16439 14504 17224 14532
rect 16439 14501 16451 14504
rect 16393 14495 16451 14501
rect 17218 14492 17224 14504
rect 17276 14492 17282 14544
rect 18322 14492 18328 14544
rect 18380 14492 18386 14544
rect 24670 14492 24676 14544
rect 24728 14532 24734 14544
rect 24728 14504 24900 14532
rect 24728 14492 24734 14504
rect 15746 14464 15752 14476
rect 15707 14436 15752 14464
rect 15746 14424 15752 14436
rect 15804 14424 15810 14476
rect 18233 14467 18291 14473
rect 18233 14433 18245 14467
rect 18279 14464 18291 14467
rect 18340 14464 18368 14492
rect 18279 14436 18368 14464
rect 18693 14467 18751 14473
rect 18279 14433 18291 14436
rect 18233 14427 18291 14433
rect 18693 14433 18705 14467
rect 18739 14464 18751 14467
rect 19426 14464 19432 14476
rect 18739 14436 19432 14464
rect 18739 14433 18751 14436
rect 18693 14427 18751 14433
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 19889 14467 19947 14473
rect 19889 14433 19901 14467
rect 19935 14464 19947 14467
rect 20530 14464 20536 14476
rect 19935 14436 20536 14464
rect 19935 14433 19947 14436
rect 19889 14427 19947 14433
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 24762 14464 24768 14476
rect 20640 14436 24768 14464
rect 6546 14396 6552 14408
rect 6507 14368 6552 14396
rect 6546 14356 6552 14368
rect 6604 14356 6610 14408
rect 8202 14396 8208 14408
rect 8163 14368 8208 14396
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 10134 14396 10140 14408
rect 10095 14368 10140 14396
rect 10134 14356 10140 14368
rect 10192 14356 10198 14408
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 16209 14399 16267 14405
rect 16209 14396 16221 14399
rect 14424 14368 16221 14396
rect 14424 14356 14430 14368
rect 16209 14365 16221 14368
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14396 16451 14399
rect 16758 14396 16764 14408
rect 16439 14368 16764 14396
rect 16439 14365 16451 14368
rect 16393 14359 16451 14365
rect 16758 14356 16764 14368
rect 16816 14356 16822 14408
rect 16853 14399 16911 14405
rect 16853 14365 16865 14399
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 15504 14331 15562 14337
rect 15504 14297 15516 14331
rect 15550 14328 15562 14331
rect 16114 14328 16120 14340
rect 15550 14300 16120 14328
rect 15550 14297 15562 14300
rect 15504 14291 15562 14297
rect 16114 14288 16120 14300
rect 16172 14288 16178 14340
rect 16868 14328 16896 14359
rect 16942 14356 16948 14408
rect 17000 14396 17006 14408
rect 17497 14399 17555 14405
rect 17497 14396 17509 14399
rect 17000 14368 17509 14396
rect 17000 14356 17006 14368
rect 17497 14365 17509 14368
rect 17543 14365 17555 14399
rect 17497 14359 17555 14365
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 18506 14396 18512 14408
rect 18371 14368 18512 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 18506 14356 18512 14368
rect 18564 14396 18570 14408
rect 19242 14396 19248 14408
rect 18564 14368 19248 14396
rect 18564 14356 18570 14368
rect 19242 14356 19248 14368
rect 19300 14356 19306 14408
rect 19610 14396 19616 14408
rect 19571 14368 19616 14396
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 19705 14399 19763 14405
rect 19705 14365 19717 14399
rect 19751 14396 19763 14399
rect 20640 14396 20668 14436
rect 24762 14424 24768 14436
rect 24820 14424 24826 14476
rect 24872 14464 24900 14504
rect 28166 14492 28172 14544
rect 28224 14532 28230 14544
rect 28629 14535 28687 14541
rect 28629 14532 28641 14535
rect 28224 14504 28641 14532
rect 28224 14492 28230 14504
rect 28629 14501 28641 14504
rect 28675 14501 28687 14535
rect 35526 14532 35532 14544
rect 28629 14495 28687 14501
rect 28736 14504 35532 14532
rect 28736 14464 28764 14504
rect 35526 14492 35532 14504
rect 35584 14492 35590 14544
rect 39224 14532 39252 14560
rect 40957 14535 41015 14541
rect 40957 14532 40969 14535
rect 39224 14504 40969 14532
rect 40957 14501 40969 14504
rect 41003 14501 41015 14535
rect 40957 14495 41015 14501
rect 48682 14492 48688 14544
rect 48740 14532 48746 14544
rect 56318 14532 56324 14544
rect 48740 14504 56324 14532
rect 48740 14492 48746 14504
rect 56318 14492 56324 14504
rect 56376 14492 56382 14544
rect 24872 14436 28764 14464
rect 28997 14467 29055 14473
rect 28997 14433 29009 14467
rect 29043 14464 29055 14467
rect 30098 14464 30104 14476
rect 29043 14436 30104 14464
rect 29043 14433 29055 14436
rect 28997 14427 29055 14433
rect 30098 14424 30104 14436
rect 30156 14424 30162 14476
rect 31938 14464 31944 14476
rect 31899 14436 31944 14464
rect 31938 14424 31944 14436
rect 31996 14424 32002 14476
rect 37182 14424 37188 14476
rect 37240 14464 37246 14476
rect 38289 14467 38347 14473
rect 38289 14464 38301 14467
rect 37240 14436 38301 14464
rect 37240 14424 37246 14436
rect 38289 14433 38301 14436
rect 38335 14464 38347 14467
rect 39945 14467 40003 14473
rect 38335 14436 38608 14464
rect 38335 14433 38347 14436
rect 38289 14427 38347 14433
rect 19751 14368 20668 14396
rect 20717 14399 20775 14405
rect 19751 14365 19763 14368
rect 19705 14359 19763 14365
rect 20717 14365 20729 14399
rect 20763 14396 20775 14399
rect 20898 14396 20904 14408
rect 20763 14368 20904 14396
rect 20763 14365 20775 14368
rect 20717 14359 20775 14365
rect 16868 14300 19288 14328
rect 7098 14260 7104 14272
rect 7059 14232 7104 14260
rect 7098 14220 7104 14232
rect 7156 14220 7162 14272
rect 7374 14220 7380 14272
rect 7432 14260 7438 14272
rect 8297 14263 8355 14269
rect 8297 14260 8309 14263
rect 7432 14232 8309 14260
rect 7432 14220 7438 14232
rect 8297 14229 8309 14232
rect 8343 14229 8355 14263
rect 8297 14223 8355 14229
rect 14369 14263 14427 14269
rect 14369 14229 14381 14263
rect 14415 14260 14427 14263
rect 15194 14260 15200 14272
rect 14415 14232 15200 14260
rect 14415 14229 14427 14232
rect 14369 14223 14427 14229
rect 15194 14220 15200 14232
rect 15252 14220 15258 14272
rect 17589 14263 17647 14269
rect 17589 14229 17601 14263
rect 17635 14260 17647 14263
rect 19150 14260 19156 14272
rect 17635 14232 19156 14260
rect 17635 14229 17647 14232
rect 17589 14223 17647 14229
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 19260 14269 19288 14300
rect 19245 14263 19303 14269
rect 19245 14229 19257 14263
rect 19291 14229 19303 14263
rect 19245 14223 19303 14229
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19720 14260 19748 14359
rect 20898 14356 20904 14368
rect 20956 14356 20962 14408
rect 21177 14399 21235 14405
rect 21177 14365 21189 14399
rect 21223 14365 21235 14399
rect 21177 14359 21235 14365
rect 19794 14288 19800 14340
rect 19852 14328 19858 14340
rect 21192 14328 21220 14359
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 22281 14399 22339 14405
rect 22281 14396 22293 14399
rect 22152 14368 22293 14396
rect 22152 14356 22158 14368
rect 22281 14365 22293 14368
rect 22327 14365 22339 14399
rect 22281 14359 22339 14365
rect 23109 14399 23167 14405
rect 23109 14365 23121 14399
rect 23155 14396 23167 14399
rect 23658 14396 23664 14408
rect 23155 14368 23664 14396
rect 23155 14365 23167 14368
rect 23109 14359 23167 14365
rect 23658 14356 23664 14368
rect 23716 14356 23722 14408
rect 29362 14356 29368 14408
rect 29420 14396 29426 14408
rect 29549 14399 29607 14405
rect 29549 14396 29561 14399
rect 29420 14368 29561 14396
rect 29420 14356 29426 14368
rect 29549 14365 29561 14368
rect 29595 14365 29607 14399
rect 29549 14359 29607 14365
rect 29825 14399 29883 14405
rect 29825 14365 29837 14399
rect 29871 14396 29883 14399
rect 30558 14396 30564 14408
rect 29871 14368 30564 14396
rect 29871 14365 29883 14368
rect 29825 14359 29883 14365
rect 30558 14356 30564 14368
rect 30616 14356 30622 14408
rect 32033 14399 32091 14405
rect 32033 14365 32045 14399
rect 32079 14396 32091 14399
rect 32766 14396 32772 14408
rect 32079 14368 32772 14396
rect 32079 14365 32091 14368
rect 32033 14359 32091 14365
rect 32766 14356 32772 14368
rect 32824 14356 32830 14408
rect 33134 14396 33140 14408
rect 33095 14368 33140 14396
rect 33134 14356 33140 14368
rect 33192 14356 33198 14408
rect 35897 14399 35955 14405
rect 35897 14365 35909 14399
rect 35943 14396 35955 14399
rect 38470 14396 38476 14408
rect 35943 14368 38476 14396
rect 35943 14365 35955 14368
rect 35897 14359 35955 14365
rect 38470 14356 38476 14368
rect 38528 14356 38534 14408
rect 19852 14300 21220 14328
rect 19852 14288 19858 14300
rect 21634 14288 21640 14340
rect 21692 14328 21698 14340
rect 22557 14331 22615 14337
rect 22557 14328 22569 14331
rect 21692 14300 22569 14328
rect 21692 14288 21698 14300
rect 22557 14297 22569 14300
rect 22603 14328 22615 14331
rect 23290 14328 23296 14340
rect 22603 14300 23296 14328
rect 22603 14297 22615 14300
rect 22557 14291 22615 14297
rect 23290 14288 23296 14300
rect 23348 14288 23354 14340
rect 26510 14328 26516 14340
rect 25240 14300 26516 14328
rect 19392 14232 19748 14260
rect 19392 14220 19398 14232
rect 20990 14220 20996 14272
rect 21048 14260 21054 14272
rect 21269 14263 21327 14269
rect 21269 14260 21281 14263
rect 21048 14232 21281 14260
rect 21048 14220 21054 14232
rect 21269 14229 21281 14232
rect 21315 14229 21327 14263
rect 21269 14223 21327 14229
rect 21726 14220 21732 14272
rect 21784 14260 21790 14272
rect 22373 14263 22431 14269
rect 22373 14260 22385 14263
rect 21784 14232 22385 14260
rect 21784 14220 21790 14232
rect 22373 14229 22385 14232
rect 22419 14260 22431 14263
rect 25240 14260 25268 14300
rect 26510 14288 26516 14300
rect 26568 14288 26574 14340
rect 36170 14337 36176 14340
rect 36164 14291 36176 14337
rect 36228 14328 36234 14340
rect 36228 14300 36264 14328
rect 36170 14288 36176 14291
rect 36228 14288 36234 14300
rect 37274 14288 37280 14340
rect 37332 14328 37338 14340
rect 38197 14331 38255 14337
rect 38197 14328 38209 14331
rect 37332 14300 38209 14328
rect 37332 14288 37338 14300
rect 38197 14297 38209 14300
rect 38243 14297 38255 14331
rect 38580 14328 38608 14436
rect 39945 14433 39957 14467
rect 39991 14433 40003 14467
rect 42705 14467 42763 14473
rect 42705 14464 42717 14467
rect 39945 14427 40003 14433
rect 41386 14436 42717 14464
rect 38746 14356 38752 14408
rect 38804 14396 38810 14408
rect 39117 14399 39175 14405
rect 39117 14396 39129 14399
rect 38804 14368 39129 14396
rect 38804 14356 38810 14368
rect 39117 14365 39129 14368
rect 39163 14396 39175 14399
rect 39850 14396 39856 14408
rect 39163 14368 39856 14396
rect 39163 14365 39175 14368
rect 39117 14359 39175 14365
rect 39850 14356 39856 14368
rect 39908 14396 39914 14408
rect 39960 14396 39988 14427
rect 39908 14368 39988 14396
rect 39908 14356 39914 14368
rect 40034 14356 40040 14408
rect 40092 14396 40098 14408
rect 40862 14396 40868 14408
rect 40092 14368 40137 14396
rect 40823 14368 40868 14396
rect 40092 14356 40098 14368
rect 40862 14356 40868 14368
rect 40920 14356 40926 14408
rect 41138 14396 41144 14408
rect 41099 14368 41144 14396
rect 41138 14356 41144 14368
rect 41196 14356 41202 14408
rect 41386 14328 41414 14436
rect 42705 14433 42717 14436
rect 42751 14464 42763 14467
rect 43441 14467 43499 14473
rect 43441 14464 43453 14467
rect 42751 14436 43453 14464
rect 42751 14433 42763 14436
rect 42705 14427 42763 14433
rect 43441 14433 43453 14436
rect 43487 14433 43499 14467
rect 43441 14427 43499 14433
rect 42521 14399 42579 14405
rect 42521 14365 42533 14399
rect 42567 14396 42579 14399
rect 42610 14396 42616 14408
rect 42567 14368 42616 14396
rect 42567 14365 42579 14368
rect 42521 14359 42579 14365
rect 42610 14356 42616 14368
rect 42668 14356 42674 14408
rect 43625 14399 43683 14405
rect 43625 14365 43637 14399
rect 43671 14396 43683 14399
rect 45186 14396 45192 14408
rect 43671 14368 45192 14396
rect 43671 14365 43683 14368
rect 43625 14359 43683 14365
rect 45186 14356 45192 14368
rect 45244 14396 45250 14408
rect 45373 14399 45431 14405
rect 45373 14396 45385 14399
rect 45244 14368 45385 14396
rect 45244 14356 45250 14368
rect 45373 14365 45385 14368
rect 45419 14365 45431 14399
rect 45373 14359 45431 14365
rect 45462 14356 45468 14408
rect 45520 14396 45526 14408
rect 45649 14399 45707 14405
rect 45649 14396 45661 14399
rect 45520 14368 45661 14396
rect 45520 14356 45526 14368
rect 45649 14365 45661 14368
rect 45695 14365 45707 14399
rect 45649 14359 45707 14365
rect 38580 14300 41414 14328
rect 38197 14291 38255 14297
rect 43346 14288 43352 14340
rect 43404 14328 43410 14340
rect 45005 14331 45063 14337
rect 45005 14328 45017 14331
rect 43404 14300 45017 14328
rect 43404 14288 43410 14300
rect 45005 14297 45017 14300
rect 45051 14297 45063 14331
rect 45005 14291 45063 14297
rect 26418 14260 26424 14272
rect 22419 14232 25268 14260
rect 26379 14232 26424 14260
rect 22419 14229 22431 14232
rect 22373 14223 22431 14229
rect 26418 14220 26424 14232
rect 26476 14220 26482 14272
rect 27430 14260 27436 14272
rect 27391 14232 27436 14260
rect 27430 14220 27436 14232
rect 27488 14220 27494 14272
rect 29730 14260 29736 14272
rect 29691 14232 29736 14260
rect 29730 14220 29736 14232
rect 29788 14220 29794 14272
rect 33321 14263 33379 14269
rect 33321 14229 33333 14263
rect 33367 14260 33379 14263
rect 33410 14260 33416 14272
rect 33367 14232 33416 14260
rect 33367 14229 33379 14232
rect 33321 14223 33379 14229
rect 33410 14220 33416 14232
rect 33468 14220 33474 14272
rect 37366 14220 37372 14272
rect 37424 14260 37430 14272
rect 37737 14263 37795 14269
rect 37737 14260 37749 14263
rect 37424 14232 37749 14260
rect 37424 14220 37430 14232
rect 37737 14229 37749 14232
rect 37783 14229 37795 14263
rect 38102 14260 38108 14272
rect 38063 14232 38108 14260
rect 37737 14223 37795 14229
rect 38102 14220 38108 14232
rect 38160 14220 38166 14272
rect 41690 14220 41696 14272
rect 41748 14260 41754 14272
rect 42153 14263 42211 14269
rect 42153 14260 42165 14263
rect 41748 14232 42165 14260
rect 41748 14220 41754 14232
rect 42153 14229 42165 14232
rect 42199 14229 42211 14263
rect 42153 14223 42211 14229
rect 42613 14263 42671 14269
rect 42613 14229 42625 14263
rect 42659 14260 42671 14263
rect 43070 14260 43076 14272
rect 42659 14232 43076 14260
rect 42659 14229 42671 14232
rect 42613 14223 42671 14229
rect 43070 14220 43076 14232
rect 43128 14220 43134 14272
rect 43622 14220 43628 14272
rect 43680 14260 43686 14272
rect 43717 14263 43775 14269
rect 43717 14260 43729 14263
rect 43680 14232 43729 14260
rect 43680 14220 43686 14232
rect 43717 14229 43729 14232
rect 43763 14229 43775 14263
rect 43717 14223 43775 14229
rect 44085 14263 44143 14269
rect 44085 14229 44097 14263
rect 44131 14260 44143 14263
rect 44174 14260 44180 14272
rect 44131 14232 44180 14260
rect 44131 14229 44143 14232
rect 44085 14223 44143 14229
rect 44174 14220 44180 14232
rect 44232 14220 44238 14272
rect 1104 14170 68816 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 68816 14170
rect 1104 14096 68816 14118
rect 11885 14059 11943 14065
rect 11885 14025 11897 14059
rect 11931 14056 11943 14059
rect 12066 14056 12072 14068
rect 11931 14028 12072 14056
rect 11931 14025 11943 14028
rect 11885 14019 11943 14025
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 15013 14059 15071 14065
rect 15013 14025 15025 14059
rect 15059 14056 15071 14059
rect 15194 14056 15200 14068
rect 15059 14028 15200 14056
rect 15059 14025 15071 14028
rect 15013 14019 15071 14025
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 16758 14056 16764 14068
rect 16719 14028 16764 14056
rect 16758 14016 16764 14028
rect 16816 14056 16822 14068
rect 17494 14056 17500 14068
rect 16816 14028 17500 14056
rect 16816 14016 16822 14028
rect 17494 14016 17500 14028
rect 17552 14016 17558 14068
rect 18877 14059 18935 14065
rect 18877 14025 18889 14059
rect 18923 14056 18935 14059
rect 19334 14056 19340 14068
rect 18923 14028 19340 14056
rect 18923 14025 18935 14028
rect 18877 14019 18935 14025
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 20533 14059 20591 14065
rect 19904 14028 20208 14056
rect 11977 13991 12035 13997
rect 11977 13957 11989 13991
rect 12023 13988 12035 13991
rect 12526 13988 12532 14000
rect 12023 13960 12532 13988
rect 12023 13957 12035 13960
rect 11977 13951 12035 13957
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 13814 13988 13820 14000
rect 13775 13960 13820 13988
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 16390 13988 16396 14000
rect 14016 13960 16396 13988
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13920 4767 13923
rect 4890 13920 4896 13932
rect 4755 13892 4896 13920
rect 4755 13889 4767 13892
rect 4709 13883 4767 13889
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 10778 13920 10784 13932
rect 10739 13892 10784 13920
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 14016 13929 14044 13960
rect 16390 13948 16396 13960
rect 16448 13948 16454 14000
rect 17218 13948 17224 14000
rect 17276 13988 17282 14000
rect 18141 13991 18199 13997
rect 18141 13988 18153 13991
rect 17276 13960 18153 13988
rect 17276 13948 17282 13960
rect 18141 13957 18153 13960
rect 18187 13957 18199 13991
rect 19904 13988 19932 14028
rect 20180 13997 20208 14028
rect 20272 14028 20484 14056
rect 20272 13997 20300 14028
rect 18141 13951 18199 13957
rect 19352 13960 19932 13988
rect 20165 13991 20223 13997
rect 12805 13923 12863 13929
rect 12805 13889 12817 13923
rect 12851 13920 12863 13923
rect 14001 13923 14059 13929
rect 14001 13920 14013 13923
rect 12851 13892 14013 13920
rect 12851 13889 12863 13892
rect 12805 13883 12863 13889
rect 14001 13889 14013 13892
rect 14047 13889 14059 13923
rect 14001 13883 14059 13889
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13920 14243 13923
rect 14366 13920 14372 13932
rect 14231 13892 14372 13920
rect 14231 13889 14243 13892
rect 14185 13883 14243 13889
rect 14366 13880 14372 13892
rect 14424 13880 14430 13932
rect 14918 13920 14924 13932
rect 14568 13892 14924 13920
rect 6730 13852 6736 13864
rect 6691 13824 6736 13852
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 10870 13852 10876 13864
rect 10551 13824 10876 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 10870 13812 10876 13824
rect 10928 13812 10934 13864
rect 12161 13855 12219 13861
rect 12161 13821 12173 13855
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 13357 13855 13415 13861
rect 13357 13821 13369 13855
rect 13403 13852 13415 13855
rect 14568 13852 14596 13892
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 19150 13880 19156 13932
rect 19208 13920 19214 13932
rect 19352 13929 19380 13960
rect 20165 13957 20177 13991
rect 20211 13957 20223 13991
rect 20165 13951 20223 13957
rect 20257 13991 20315 13997
rect 20257 13957 20269 13991
rect 20303 13957 20315 13991
rect 20456 13988 20484 14028
rect 20533 14025 20545 14059
rect 20579 14056 20591 14059
rect 20714 14056 20720 14068
rect 20579 14028 20720 14056
rect 20579 14025 20591 14028
rect 20533 14019 20591 14025
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 23290 14056 23296 14068
rect 23251 14028 23296 14056
rect 23290 14016 23296 14028
rect 23348 14016 23354 14068
rect 23658 14056 23664 14068
rect 23619 14028 23664 14056
rect 23658 14016 23664 14028
rect 23716 14016 23722 14068
rect 26418 14056 26424 14068
rect 26252 14028 26424 14056
rect 21634 13988 21640 14000
rect 20456 13960 21640 13988
rect 20257 13951 20315 13957
rect 19337 13923 19395 13929
rect 19337 13920 19349 13923
rect 19208 13892 19349 13920
rect 19208 13880 19214 13892
rect 19337 13889 19349 13892
rect 19383 13889 19395 13923
rect 19337 13883 19395 13889
rect 19521 13923 19579 13929
rect 19521 13889 19533 13923
rect 19567 13920 19579 13923
rect 19886 13920 19892 13932
rect 19567 13892 19892 13920
rect 19567 13889 19579 13892
rect 19521 13883 19579 13889
rect 19886 13880 19892 13892
rect 19944 13920 19950 13932
rect 19981 13923 20039 13929
rect 19981 13920 19993 13923
rect 19944 13892 19993 13920
rect 19944 13880 19950 13892
rect 19981 13889 19993 13892
rect 20027 13889 20039 13923
rect 19981 13883 20039 13889
rect 20349 13923 20407 13929
rect 20349 13889 20361 13923
rect 20395 13920 20407 13923
rect 20990 13920 20996 13932
rect 20395 13892 20996 13920
rect 20395 13889 20407 13892
rect 20349 13883 20407 13889
rect 20990 13880 20996 13892
rect 21048 13880 21054 13932
rect 21192 13929 21220 13960
rect 21634 13948 21640 13960
rect 21692 13948 21698 14000
rect 26252 13997 26280 14028
rect 26418 14016 26424 14028
rect 26476 14056 26482 14068
rect 35986 14056 35992 14068
rect 26476 14028 35992 14056
rect 26476 14016 26482 14028
rect 35986 14016 35992 14028
rect 36044 14016 36050 14068
rect 36170 14056 36176 14068
rect 36131 14028 36176 14056
rect 36170 14016 36176 14028
rect 36228 14016 36234 14068
rect 39850 14056 39856 14068
rect 39811 14028 39856 14056
rect 39850 14016 39856 14028
rect 39908 14016 39914 14068
rect 41877 14059 41935 14065
rect 41877 14025 41889 14059
rect 41923 14025 41935 14059
rect 41877 14019 41935 14025
rect 26237 13991 26295 13997
rect 26237 13957 26249 13991
rect 26283 13957 26295 13991
rect 26237 13951 26295 13957
rect 35618 13948 35624 14000
rect 35676 13988 35682 14000
rect 35713 13991 35771 13997
rect 35713 13988 35725 13991
rect 35676 13960 35725 13988
rect 35676 13948 35682 13960
rect 35713 13957 35725 13960
rect 35759 13988 35771 13991
rect 39666 13988 39672 14000
rect 35759 13960 37504 13988
rect 35759 13957 35771 13960
rect 35713 13951 35771 13957
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13889 21235 13923
rect 21177 13883 21235 13889
rect 22002 13880 22008 13932
rect 22060 13920 22066 13932
rect 23201 13923 23259 13929
rect 23201 13920 23213 13923
rect 22060 13892 22105 13920
rect 23032 13892 23213 13920
rect 22060 13880 22066 13892
rect 14734 13852 14740 13864
rect 13403 13824 14596 13852
rect 14695 13824 14740 13852
rect 13403 13821 13415 13824
rect 13357 13815 13415 13821
rect 7098 13784 7104 13796
rect 7011 13756 7104 13784
rect 7098 13744 7104 13756
rect 7156 13744 7162 13796
rect 7193 13787 7251 13793
rect 7193 13753 7205 13787
rect 7239 13784 7251 13787
rect 7742 13784 7748 13796
rect 7239 13756 7748 13784
rect 7239 13753 7251 13756
rect 7193 13747 7251 13753
rect 7742 13744 7748 13756
rect 7800 13744 7806 13796
rect 10229 13787 10287 13793
rect 10229 13753 10241 13787
rect 10275 13784 10287 13787
rect 10594 13784 10600 13796
rect 10275 13756 10600 13784
rect 10275 13753 10287 13756
rect 10229 13747 10287 13753
rect 10594 13744 10600 13756
rect 10652 13744 10658 13796
rect 12176 13784 12204 13815
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15470 13812 15476 13864
rect 15528 13852 15534 13864
rect 15933 13855 15991 13861
rect 15933 13852 15945 13855
rect 15528 13824 15945 13852
rect 15528 13812 15534 13824
rect 15933 13821 15945 13824
rect 15979 13852 15991 13855
rect 18325 13855 18383 13861
rect 15979 13824 18276 13852
rect 15979 13821 15991 13824
rect 15933 13815 15991 13821
rect 12618 13784 12624 13796
rect 12176 13756 12624 13784
rect 12618 13744 12624 13756
rect 12676 13744 12682 13796
rect 15381 13787 15439 13793
rect 15381 13753 15393 13787
rect 15427 13784 15439 13787
rect 16482 13784 16488 13796
rect 15427 13756 16488 13784
rect 15427 13753 15439 13756
rect 15381 13747 15439 13753
rect 16482 13744 16488 13756
rect 16540 13744 16546 13796
rect 18248 13784 18276 13824
rect 18325 13821 18337 13855
rect 18371 13852 18383 13855
rect 20530 13852 20536 13864
rect 18371 13824 20536 13852
rect 18371 13821 18383 13824
rect 18325 13815 18383 13821
rect 20530 13812 20536 13824
rect 20588 13812 20594 13864
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 21085 13855 21143 13861
rect 21085 13852 21097 13855
rect 20864 13824 21097 13852
rect 20864 13812 20870 13824
rect 21085 13821 21097 13824
rect 21131 13821 21143 13855
rect 21085 13815 21143 13821
rect 23032 13784 23060 13892
rect 23201 13889 23213 13892
rect 23247 13920 23259 13923
rect 23382 13920 23388 13932
rect 23247 13892 23388 13920
rect 23247 13889 23259 13892
rect 23201 13883 23259 13889
rect 23382 13880 23388 13892
rect 23440 13880 23446 13932
rect 25314 13880 25320 13932
rect 25372 13920 25378 13932
rect 25501 13923 25559 13929
rect 25501 13920 25513 13923
rect 25372 13892 25513 13920
rect 25372 13880 25378 13892
rect 25501 13889 25513 13892
rect 25547 13889 25559 13923
rect 25501 13883 25559 13889
rect 26421 13923 26479 13929
rect 26421 13889 26433 13923
rect 26467 13920 26479 13923
rect 26510 13920 26516 13932
rect 26467 13892 26516 13920
rect 26467 13889 26479 13892
rect 26421 13883 26479 13889
rect 26510 13880 26516 13892
rect 26568 13880 26574 13932
rect 33410 13929 33416 13932
rect 33404 13920 33416 13929
rect 33371 13892 33416 13920
rect 33404 13883 33416 13892
rect 33410 13880 33416 13883
rect 33468 13880 33474 13932
rect 36357 13923 36415 13929
rect 36357 13889 36369 13923
rect 36403 13920 36415 13923
rect 37366 13920 37372 13932
rect 36403 13892 37372 13920
rect 36403 13889 36415 13892
rect 36357 13883 36415 13889
rect 37366 13880 37372 13892
rect 37424 13880 37430 13932
rect 37476 13929 37504 13960
rect 37844 13960 39672 13988
rect 37461 13923 37519 13929
rect 37461 13889 37473 13923
rect 37507 13889 37519 13923
rect 37461 13883 37519 13889
rect 23109 13855 23167 13861
rect 23109 13821 23121 13855
rect 23155 13821 23167 13855
rect 25682 13852 25688 13864
rect 25643 13824 25688 13852
rect 23109 13815 23167 13821
rect 18248 13756 23060 13784
rect 23124 13784 23152 13815
rect 25682 13812 25688 13824
rect 25740 13812 25746 13864
rect 26326 13812 26332 13864
rect 26384 13852 26390 13864
rect 27430 13852 27436 13864
rect 26384 13824 27436 13852
rect 26384 13812 26390 13824
rect 27430 13812 27436 13824
rect 27488 13812 27494 13864
rect 27709 13855 27767 13861
rect 27709 13821 27721 13855
rect 27755 13852 27767 13855
rect 27755 13824 29224 13852
rect 27755 13821 27767 13824
rect 27709 13815 27767 13821
rect 27062 13784 27068 13796
rect 23124 13756 27068 13784
rect 27062 13744 27068 13756
rect 27120 13744 27126 13796
rect 29196 13784 29224 13824
rect 32858 13812 32864 13864
rect 32916 13852 32922 13864
rect 33137 13855 33195 13861
rect 33137 13852 33149 13855
rect 32916 13824 33149 13852
rect 32916 13812 32922 13824
rect 33137 13821 33149 13824
rect 33183 13821 33195 13855
rect 33137 13815 33195 13821
rect 37274 13812 37280 13864
rect 37332 13852 37338 13864
rect 37844 13861 37872 13960
rect 39666 13948 39672 13960
rect 39724 13948 39730 14000
rect 41892 13988 41920 14019
rect 43162 14016 43168 14068
rect 43220 14056 43226 14068
rect 44269 14059 44327 14065
rect 44269 14056 44281 14059
rect 43220 14028 44281 14056
rect 43220 14016 43226 14028
rect 44269 14025 44281 14028
rect 44315 14025 44327 14059
rect 44269 14019 44327 14025
rect 42674 13991 42732 13997
rect 42674 13988 42686 13991
rect 41892 13960 42686 13988
rect 42674 13957 42686 13960
rect 42720 13957 42732 13991
rect 42674 13951 42732 13957
rect 44729 13991 44787 13997
rect 44729 13957 44741 13991
rect 44775 13988 44787 13991
rect 45186 13988 45192 14000
rect 44775 13960 45192 13988
rect 44775 13957 44787 13960
rect 44729 13951 44787 13957
rect 45186 13948 45192 13960
rect 45244 13948 45250 14000
rect 38470 13920 38476 13932
rect 38431 13892 38476 13920
rect 38470 13880 38476 13892
rect 38528 13880 38534 13932
rect 38746 13929 38752 13932
rect 38740 13883 38752 13929
rect 38804 13920 38810 13932
rect 41690 13920 41696 13932
rect 38804 13892 38840 13920
rect 41651 13892 41696 13920
rect 38746 13880 38752 13883
rect 38804 13880 38810 13892
rect 41690 13880 41696 13892
rect 41748 13880 41754 13932
rect 37553 13855 37611 13861
rect 37553 13852 37565 13855
rect 37332 13824 37565 13852
rect 37332 13812 37338 13824
rect 37553 13821 37565 13824
rect 37599 13821 37611 13855
rect 37553 13815 37611 13821
rect 37829 13855 37887 13861
rect 37829 13821 37841 13855
rect 37875 13821 37887 13855
rect 37829 13815 37887 13821
rect 39850 13812 39856 13864
rect 39908 13852 39914 13864
rect 40681 13855 40739 13861
rect 40681 13852 40693 13855
rect 39908 13824 40693 13852
rect 39908 13812 39914 13824
rect 40681 13821 40693 13824
rect 40727 13852 40739 13855
rect 40862 13852 40868 13864
rect 40727 13824 40868 13852
rect 40727 13821 40739 13824
rect 40681 13815 40739 13821
rect 40862 13812 40868 13824
rect 40920 13812 40926 13864
rect 41598 13812 41604 13864
rect 41656 13852 41662 13864
rect 42426 13852 42432 13864
rect 41656 13824 42432 13852
rect 41656 13812 41662 13824
rect 42426 13812 42432 13824
rect 42484 13812 42490 13864
rect 29822 13784 29828 13796
rect 29196 13756 29828 13784
rect 29822 13744 29828 13756
rect 29880 13784 29886 13796
rect 32490 13784 32496 13796
rect 29880 13756 32496 13784
rect 29880 13744 29886 13756
rect 32490 13744 32496 13756
rect 32548 13744 32554 13796
rect 32582 13744 32588 13796
rect 32640 13784 32646 13796
rect 33042 13784 33048 13796
rect 32640 13756 33048 13784
rect 32640 13744 32646 13756
rect 33042 13744 33048 13756
rect 33100 13744 33106 13796
rect 44358 13784 44364 13796
rect 44319 13756 44364 13784
rect 44358 13744 44364 13756
rect 44416 13784 44422 13796
rect 45189 13787 45247 13793
rect 45189 13784 45201 13787
rect 44416 13756 45201 13784
rect 44416 13744 44422 13756
rect 45189 13753 45201 13756
rect 45235 13784 45247 13787
rect 45462 13784 45468 13796
rect 45235 13756 45468 13784
rect 45235 13753 45247 13756
rect 45189 13747 45247 13753
rect 45462 13744 45468 13756
rect 45520 13744 45526 13796
rect 4893 13719 4951 13725
rect 4893 13685 4905 13719
rect 4939 13716 4951 13719
rect 4982 13716 4988 13728
rect 4939 13688 4988 13716
rect 4939 13685 4951 13688
rect 4893 13679 4951 13685
rect 4982 13676 4988 13688
rect 5040 13676 5046 13728
rect 7116 13716 7144 13744
rect 7650 13716 7656 13728
rect 7116 13688 7656 13716
rect 7650 13676 7656 13688
rect 7708 13676 7714 13728
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 10413 13719 10471 13725
rect 10413 13716 10425 13719
rect 9824 13688 10425 13716
rect 9824 13676 9830 13688
rect 10413 13685 10425 13688
rect 10459 13685 10471 13719
rect 10413 13679 10471 13685
rect 11517 13719 11575 13725
rect 11517 13685 11529 13719
rect 11563 13716 11575 13719
rect 11698 13716 11704 13728
rect 11563 13688 11704 13716
rect 11563 13685 11575 13688
rect 11517 13679 11575 13685
rect 11698 13676 11704 13688
rect 11756 13676 11762 13728
rect 19334 13716 19340 13728
rect 19295 13688 19340 13716
rect 19334 13676 19340 13688
rect 19392 13676 19398 13728
rect 19886 13676 19892 13728
rect 19944 13716 19950 13728
rect 21082 13716 21088 13728
rect 19944 13688 21088 13716
rect 19944 13676 19950 13688
rect 21082 13676 21088 13688
rect 21140 13676 21146 13728
rect 21818 13716 21824 13728
rect 21779 13688 21824 13716
rect 21818 13676 21824 13688
rect 21876 13676 21882 13728
rect 34514 13716 34520 13728
rect 34475 13688 34520 13716
rect 34514 13676 34520 13688
rect 34572 13676 34578 13728
rect 43070 13676 43076 13728
rect 43128 13716 43134 13728
rect 43809 13719 43867 13725
rect 43809 13716 43821 13719
rect 43128 13688 43821 13716
rect 43128 13676 43134 13688
rect 43809 13685 43821 13688
rect 43855 13685 43867 13719
rect 43809 13679 43867 13685
rect 1104 13626 68816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 65654 13626
rect 65706 13574 65718 13626
rect 65770 13574 65782 13626
rect 65834 13574 65846 13626
rect 65898 13574 65910 13626
rect 65962 13574 68816 13626
rect 1104 13552 68816 13574
rect 6825 13515 6883 13521
rect 6825 13481 6837 13515
rect 6871 13512 6883 13515
rect 7650 13512 7656 13524
rect 6871 13484 7656 13512
rect 6871 13481 6883 13484
rect 6825 13475 6883 13481
rect 7650 13472 7656 13484
rect 7708 13472 7714 13524
rect 11885 13515 11943 13521
rect 11885 13481 11897 13515
rect 11931 13512 11943 13515
rect 12066 13512 12072 13524
rect 11931 13484 12072 13512
rect 11931 13481 11943 13484
rect 11885 13475 11943 13481
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 14553 13515 14611 13521
rect 14553 13481 14565 13515
rect 14599 13512 14611 13515
rect 14734 13512 14740 13524
rect 14599 13484 14740 13512
rect 14599 13481 14611 13484
rect 14553 13475 14611 13481
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 16114 13472 16120 13524
rect 16172 13512 16178 13524
rect 16301 13515 16359 13521
rect 16301 13512 16313 13515
rect 16172 13484 16313 13512
rect 16172 13472 16178 13484
rect 16301 13481 16313 13484
rect 16347 13481 16359 13515
rect 16301 13475 16359 13481
rect 16390 13472 16396 13524
rect 16448 13512 16454 13524
rect 16945 13515 17003 13521
rect 16945 13512 16957 13515
rect 16448 13484 16957 13512
rect 16448 13472 16454 13484
rect 16945 13481 16957 13484
rect 16991 13481 17003 13515
rect 18230 13512 18236 13524
rect 18191 13484 18236 13512
rect 16945 13475 17003 13481
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 19150 13472 19156 13524
rect 19208 13512 19214 13524
rect 19208 13484 20576 13512
rect 19208 13472 19214 13484
rect 15657 13447 15715 13453
rect 15657 13444 15669 13447
rect 14660 13416 15669 13444
rect 7009 13379 7067 13385
rect 7009 13345 7021 13379
rect 7055 13345 7067 13379
rect 7009 13339 7067 13345
rect 4706 13308 4712 13320
rect 4667 13280 4712 13308
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 4982 13317 4988 13320
rect 4976 13308 4988 13317
rect 4943 13280 4988 13308
rect 4976 13271 4988 13280
rect 4982 13268 4988 13271
rect 5040 13268 5046 13320
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 6104 13280 6561 13308
rect 6104 13184 6132 13280
rect 6549 13277 6561 13280
rect 6595 13308 6607 13311
rect 6730 13308 6736 13320
rect 6595 13280 6736 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 6730 13268 6736 13280
rect 6788 13268 6794 13320
rect 7024 13308 7052 13339
rect 7469 13311 7527 13317
rect 7469 13308 7481 13311
rect 7024 13280 7481 13308
rect 7469 13277 7481 13280
rect 7515 13277 7527 13311
rect 7742 13308 7748 13320
rect 7703 13280 7748 13308
rect 7469 13271 7527 13277
rect 7742 13268 7748 13280
rect 7800 13268 7806 13320
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13308 10563 13311
rect 11514 13308 11520 13320
rect 10551 13280 11520 13308
rect 10551 13277 10563 13280
rect 10505 13271 10563 13277
rect 11514 13268 11520 13280
rect 11572 13308 11578 13320
rect 13081 13311 13139 13317
rect 13081 13308 13093 13311
rect 11572 13280 13093 13308
rect 11572 13268 11578 13280
rect 13081 13277 13093 13280
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 14550 13268 14556 13320
rect 14608 13308 14614 13320
rect 14660 13317 14688 13416
rect 15657 13413 15669 13416
rect 15703 13413 15715 13447
rect 15657 13407 15715 13413
rect 16206 13376 16212 13388
rect 15672 13348 16212 13376
rect 15672 13317 15700 13348
rect 16206 13336 16212 13348
rect 16264 13376 16270 13388
rect 16408 13376 16436 13472
rect 20548 13444 20576 13484
rect 20898 13472 20904 13524
rect 20956 13512 20962 13524
rect 20993 13515 21051 13521
rect 20993 13512 21005 13515
rect 20956 13484 21005 13512
rect 20956 13472 20962 13484
rect 20993 13481 21005 13484
rect 21039 13481 21051 13515
rect 28997 13515 29055 13521
rect 28997 13512 29009 13515
rect 20993 13475 21051 13481
rect 21100 13484 29009 13512
rect 21100 13444 21128 13484
rect 28997 13481 29009 13484
rect 29043 13481 29055 13515
rect 30098 13512 30104 13524
rect 30059 13484 30104 13512
rect 28997 13475 29055 13481
rect 23382 13444 23388 13456
rect 20548 13416 21128 13444
rect 23343 13416 23388 13444
rect 23382 13404 23388 13416
rect 23440 13404 23446 13456
rect 25685 13447 25743 13453
rect 25685 13413 25697 13447
rect 25731 13444 25743 13447
rect 26418 13444 26424 13456
rect 25731 13416 26424 13444
rect 25731 13413 25743 13416
rect 25685 13407 25743 13413
rect 26418 13404 26424 13416
rect 26476 13404 26482 13456
rect 29012 13444 29040 13475
rect 30098 13472 30104 13484
rect 30156 13472 30162 13524
rect 32953 13515 33011 13521
rect 32953 13481 32965 13515
rect 32999 13512 33011 13515
rect 33134 13512 33140 13524
rect 32999 13484 33140 13512
rect 32999 13481 33011 13484
rect 32953 13475 33011 13481
rect 33134 13472 33140 13484
rect 33192 13472 33198 13524
rect 35986 13472 35992 13524
rect 36044 13512 36050 13524
rect 36633 13515 36691 13521
rect 36633 13512 36645 13515
rect 36044 13484 36645 13512
rect 36044 13472 36050 13484
rect 36633 13481 36645 13484
rect 36679 13481 36691 13515
rect 36633 13475 36691 13481
rect 37645 13515 37703 13521
rect 37645 13481 37657 13515
rect 37691 13512 37703 13515
rect 38102 13512 38108 13524
rect 37691 13484 38108 13512
rect 37691 13481 37703 13484
rect 37645 13475 37703 13481
rect 32493 13447 32551 13453
rect 29012 13416 29776 13444
rect 16264 13348 16436 13376
rect 16264 13336 16270 13348
rect 17862 13336 17868 13388
rect 17920 13376 17926 13388
rect 19245 13379 19303 13385
rect 19245 13376 19257 13379
rect 17920 13348 19257 13376
rect 17920 13336 17926 13348
rect 19245 13345 19257 13348
rect 19291 13376 19303 13379
rect 21545 13379 21603 13385
rect 21545 13376 21557 13379
rect 19291 13348 21557 13376
rect 19291 13345 19303 13348
rect 19245 13339 19303 13345
rect 21545 13345 21557 13348
rect 21591 13345 21603 13379
rect 27522 13376 27528 13388
rect 27483 13348 27528 13376
rect 21545 13339 21603 13345
rect 27522 13336 27528 13348
rect 27580 13336 27586 13388
rect 28074 13336 28080 13388
rect 28132 13376 28138 13388
rect 29641 13379 29699 13385
rect 29641 13376 29653 13379
rect 28132 13348 29653 13376
rect 28132 13336 28138 13348
rect 29641 13345 29653 13348
rect 29687 13345 29699 13379
rect 29641 13339 29699 13345
rect 14645 13311 14703 13317
rect 14645 13308 14657 13311
rect 14608 13280 14657 13308
rect 14608 13268 14614 13280
rect 14645 13277 14657 13280
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 15657 13311 15715 13317
rect 15657 13277 15669 13311
rect 15703 13277 15715 13311
rect 15657 13271 15715 13277
rect 15746 13268 15752 13320
rect 15804 13308 15810 13320
rect 15841 13311 15899 13317
rect 15841 13308 15853 13311
rect 15804 13280 15853 13308
rect 15804 13268 15810 13280
rect 15841 13277 15853 13280
rect 15887 13277 15899 13311
rect 16482 13308 16488 13320
rect 16443 13280 16488 13308
rect 15841 13271 15899 13277
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 21818 13317 21824 13320
rect 21812 13308 21824 13317
rect 21779 13280 21824 13308
rect 21812 13271 21824 13280
rect 21818 13268 21824 13271
rect 21876 13268 21882 13320
rect 27706 13268 27712 13320
rect 27764 13308 27770 13320
rect 29748 13317 29776 13416
rect 32493 13413 32505 13447
rect 32539 13444 32551 13447
rect 33226 13444 33232 13456
rect 32539 13416 33232 13444
rect 32539 13413 32551 13416
rect 32493 13407 32551 13413
rect 33226 13404 33232 13416
rect 33284 13404 33290 13456
rect 32217 13379 32275 13385
rect 32217 13345 32229 13379
rect 32263 13376 32275 13379
rect 32582 13376 32588 13388
rect 32263 13348 32588 13376
rect 32263 13345 32275 13348
rect 32217 13339 32275 13345
rect 32582 13336 32588 13348
rect 32640 13336 32646 13388
rect 33597 13379 33655 13385
rect 33597 13345 33609 13379
rect 33643 13376 33655 13379
rect 33870 13376 33876 13388
rect 33643 13348 33876 13376
rect 33643 13345 33655 13348
rect 33597 13339 33655 13345
rect 33870 13336 33876 13348
rect 33928 13336 33934 13388
rect 28169 13311 28227 13317
rect 28169 13308 28181 13311
rect 27764 13280 28181 13308
rect 27764 13268 27770 13280
rect 28169 13277 28181 13280
rect 28215 13277 28227 13311
rect 28169 13271 28227 13277
rect 29733 13311 29791 13317
rect 29733 13277 29745 13311
rect 29779 13308 29791 13311
rect 29779 13280 31754 13308
rect 29779 13277 29791 13280
rect 29733 13271 29791 13277
rect 7561 13243 7619 13249
rect 7561 13209 7573 13243
rect 7607 13240 7619 13243
rect 8386 13240 8392 13252
rect 7607 13212 8392 13240
rect 7607 13209 7619 13212
rect 7561 13203 7619 13209
rect 8386 13200 8392 13212
rect 8444 13200 8450 13252
rect 10772 13243 10830 13249
rect 10772 13209 10784 13243
rect 10818 13240 10830 13243
rect 11422 13240 11428 13252
rect 10818 13212 11428 13240
rect 10818 13209 10830 13212
rect 10772 13203 10830 13209
rect 11422 13200 11428 13212
rect 11480 13200 11486 13252
rect 12345 13243 12403 13249
rect 12345 13209 12357 13243
rect 12391 13240 12403 13243
rect 12802 13240 12808 13252
rect 12391 13212 12808 13240
rect 12391 13209 12403 13212
rect 12345 13203 12403 13209
rect 12802 13200 12808 13212
rect 12860 13200 12866 13252
rect 14090 13200 14096 13252
rect 14148 13240 14154 13252
rect 14148 13212 17080 13240
rect 14148 13200 14154 13212
rect 6086 13172 6092 13184
rect 6047 13144 6092 13172
rect 6086 13132 6092 13144
rect 6144 13132 6150 13184
rect 7834 13132 7840 13184
rect 7892 13172 7898 13184
rect 7929 13175 7987 13181
rect 7929 13172 7941 13175
rect 7892 13144 7941 13172
rect 7892 13132 7898 13144
rect 7929 13141 7941 13144
rect 7975 13141 7987 13175
rect 17052 13172 17080 13212
rect 19426 13200 19432 13252
rect 19484 13240 19490 13252
rect 19521 13243 19579 13249
rect 19521 13240 19533 13243
rect 19484 13212 19533 13240
rect 19484 13200 19490 13212
rect 19521 13209 19533 13212
rect 19567 13209 19579 13243
rect 20898 13240 20904 13252
rect 20746 13212 20904 13240
rect 19521 13203 19579 13209
rect 20898 13200 20904 13212
rect 20956 13200 20962 13252
rect 24946 13240 24952 13252
rect 22066 13212 24952 13240
rect 22066 13172 22094 13212
rect 24946 13200 24952 13212
rect 25004 13200 25010 13252
rect 27280 13243 27338 13249
rect 27280 13209 27292 13243
rect 27326 13209 27338 13243
rect 31726 13240 31754 13280
rect 31938 13268 31944 13320
rect 31996 13308 32002 13320
rect 32125 13311 32183 13317
rect 32125 13308 32137 13311
rect 31996 13280 32137 13308
rect 31996 13268 32002 13280
rect 32125 13277 32137 13280
rect 32171 13277 32183 13311
rect 33410 13308 33416 13320
rect 33323 13280 33416 13308
rect 32125 13271 32183 13277
rect 33410 13268 33416 13280
rect 33468 13308 33474 13320
rect 34514 13308 34520 13320
rect 33468 13280 34520 13308
rect 33468 13268 33474 13280
rect 34514 13268 34520 13280
rect 34572 13268 34578 13320
rect 36648 13308 36676 13475
rect 38102 13472 38108 13484
rect 38160 13472 38166 13524
rect 38378 13512 38384 13524
rect 38339 13484 38384 13512
rect 38378 13472 38384 13484
rect 38436 13472 38442 13524
rect 38746 13472 38752 13524
rect 38804 13512 38810 13524
rect 38933 13515 38991 13521
rect 38933 13512 38945 13515
rect 38804 13484 38945 13512
rect 38804 13472 38810 13484
rect 38933 13481 38945 13484
rect 38979 13481 38991 13515
rect 38933 13475 38991 13481
rect 42242 13472 42248 13524
rect 42300 13512 42306 13524
rect 42521 13515 42579 13521
rect 42521 13512 42533 13515
rect 42300 13484 42533 13512
rect 42300 13472 42306 13484
rect 42521 13481 42533 13484
rect 42567 13481 42579 13515
rect 43346 13512 43352 13524
rect 43307 13484 43352 13512
rect 42521 13475 42579 13481
rect 43346 13472 43352 13484
rect 43404 13472 43410 13524
rect 43530 13512 43536 13524
rect 43491 13484 43536 13512
rect 43530 13472 43536 13484
rect 43588 13472 43594 13524
rect 43993 13515 44051 13521
rect 43993 13481 44005 13515
rect 44039 13512 44051 13515
rect 44082 13512 44088 13524
rect 44039 13484 44088 13512
rect 44039 13481 44051 13484
rect 43993 13475 44051 13481
rect 44082 13472 44088 13484
rect 44140 13472 44146 13524
rect 39850 13376 39856 13388
rect 38304 13348 39856 13376
rect 38304 13317 38332 13348
rect 39850 13336 39856 13348
rect 39908 13336 39914 13388
rect 42337 13379 42395 13385
rect 42337 13345 42349 13379
rect 42383 13345 42395 13379
rect 42337 13339 42395 13345
rect 38289 13311 38347 13317
rect 38289 13308 38301 13311
rect 36648 13280 38301 13308
rect 38289 13277 38301 13280
rect 38335 13277 38347 13311
rect 39114 13308 39120 13320
rect 39075 13280 39120 13308
rect 38289 13271 38347 13277
rect 39114 13268 39120 13280
rect 39172 13268 39178 13320
rect 42245 13311 42303 13317
rect 42245 13308 42257 13311
rect 41524 13280 42257 13308
rect 36446 13240 36452 13252
rect 31726 13212 36452 13240
rect 27280 13203 27338 13209
rect 17052 13144 22094 13172
rect 7929 13135 7987 13141
rect 22462 13132 22468 13184
rect 22520 13172 22526 13184
rect 22925 13175 22983 13181
rect 22925 13172 22937 13175
rect 22520 13144 22937 13172
rect 22520 13132 22526 13144
rect 22925 13141 22937 13144
rect 22971 13141 22983 13175
rect 26142 13172 26148 13184
rect 26103 13144 26148 13172
rect 22925 13135 22983 13141
rect 26142 13132 26148 13144
rect 26200 13132 26206 13184
rect 27295 13172 27323 13203
rect 36446 13200 36452 13212
rect 36504 13200 36510 13252
rect 36538 13200 36544 13252
rect 36596 13240 36602 13252
rect 38838 13240 38844 13252
rect 36596 13212 36641 13240
rect 36740 13212 38844 13240
rect 36596 13200 36602 13212
rect 27985 13175 28043 13181
rect 27985 13172 27997 13175
rect 27295 13144 27997 13172
rect 27985 13141 27997 13144
rect 28031 13141 28043 13175
rect 27985 13135 28043 13141
rect 32490 13132 32496 13184
rect 32548 13172 32554 13184
rect 33321 13175 33379 13181
rect 33321 13172 33333 13175
rect 32548 13144 33333 13172
rect 32548 13132 32554 13144
rect 33321 13141 33333 13144
rect 33367 13172 33379 13175
rect 36740 13172 36768 13212
rect 38838 13200 38844 13212
rect 38896 13200 38902 13252
rect 33367 13144 36768 13172
rect 33367 13141 33379 13144
rect 33321 13135 33379 13141
rect 41414 13132 41420 13184
rect 41472 13172 41478 13184
rect 41524 13181 41552 13280
rect 42245 13277 42257 13280
rect 42291 13277 42303 13311
rect 42352 13308 42380 13339
rect 43070 13308 43076 13320
rect 42352 13280 43076 13308
rect 42245 13271 42303 13277
rect 43070 13268 43076 13280
rect 43128 13268 43134 13320
rect 44174 13308 44180 13320
rect 44135 13280 44180 13308
rect 44174 13268 44180 13280
rect 44232 13268 44238 13320
rect 41509 13175 41567 13181
rect 41509 13172 41521 13175
rect 41472 13144 41521 13172
rect 41472 13132 41478 13144
rect 41509 13141 41521 13144
rect 41555 13141 41567 13175
rect 41509 13135 41567 13141
rect 1104 13082 68816 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 68816 13082
rect 1104 13008 68816 13030
rect 4890 12928 4896 12980
rect 4948 12968 4954 12980
rect 4985 12971 5043 12977
rect 4985 12968 4997 12971
rect 4948 12940 4997 12968
rect 4948 12928 4954 12940
rect 4985 12937 4997 12940
rect 5031 12937 5043 12971
rect 4985 12931 5043 12937
rect 5353 12971 5411 12977
rect 5353 12937 5365 12971
rect 5399 12968 5411 12971
rect 6086 12968 6092 12980
rect 5399 12940 6092 12968
rect 5399 12937 5411 12940
rect 5353 12931 5411 12937
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 7650 12968 7656 12980
rect 6472 12940 7656 12968
rect 6472 12909 6500 12940
rect 7650 12928 7656 12940
rect 7708 12968 7714 12980
rect 7708 12940 9720 12968
rect 7708 12928 7714 12940
rect 6457 12903 6515 12909
rect 6457 12869 6469 12903
rect 6503 12869 6515 12903
rect 6457 12863 6515 12869
rect 7742 12860 7748 12912
rect 7800 12900 7806 12912
rect 7800 12872 8616 12900
rect 7800 12860 7806 12872
rect 7098 12792 7104 12844
rect 7156 12832 7162 12844
rect 8588 12841 8616 12872
rect 7561 12835 7619 12841
rect 7561 12832 7573 12835
rect 7156 12804 7573 12832
rect 7156 12792 7162 12804
rect 7561 12801 7573 12804
rect 7607 12801 7619 12835
rect 7561 12795 7619 12801
rect 8389 12835 8447 12841
rect 8389 12801 8401 12835
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 8573 12835 8631 12841
rect 8573 12801 8585 12835
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 4571 12736 5457 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 5445 12733 5457 12736
rect 5491 12733 5503 12767
rect 5445 12727 5503 12733
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12764 5595 12767
rect 6454 12764 6460 12776
rect 5583 12736 6460 12764
rect 5583 12733 5595 12736
rect 5537 12727 5595 12733
rect 5460 12696 5488 12727
rect 6454 12724 6460 12736
rect 6512 12724 6518 12776
rect 7653 12767 7711 12773
rect 7653 12733 7665 12767
rect 7699 12764 7711 12767
rect 8294 12764 8300 12776
rect 7699 12736 8300 12764
rect 7699 12733 7711 12736
rect 7653 12727 7711 12733
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 5626 12696 5632 12708
rect 5460 12668 5632 12696
rect 5626 12656 5632 12668
rect 5684 12656 5690 12708
rect 6086 12656 6092 12708
rect 6144 12696 6150 12708
rect 6733 12699 6791 12705
rect 6733 12696 6745 12699
rect 6144 12668 6745 12696
rect 6144 12656 6150 12668
rect 6733 12665 6745 12668
rect 6779 12665 6791 12699
rect 6733 12659 6791 12665
rect 6917 12699 6975 12705
rect 6917 12665 6929 12699
rect 6963 12696 6975 12699
rect 8404 12696 8432 12795
rect 8662 12724 8668 12776
rect 8720 12764 8726 12776
rect 9692 12773 9720 12940
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 11517 12971 11575 12977
rect 11517 12968 11529 12971
rect 11480 12940 11529 12968
rect 11480 12928 11486 12940
rect 11517 12937 11529 12940
rect 11563 12937 11575 12971
rect 11517 12931 11575 12937
rect 13722 12928 13728 12980
rect 13780 12968 13786 12980
rect 14185 12971 14243 12977
rect 14185 12968 14197 12971
rect 13780 12940 14197 12968
rect 13780 12928 13786 12940
rect 14185 12937 14197 12940
rect 14231 12937 14243 12971
rect 14185 12931 14243 12937
rect 20073 12971 20131 12977
rect 20073 12937 20085 12971
rect 20119 12968 20131 12971
rect 20162 12968 20168 12980
rect 20119 12940 20168 12968
rect 20119 12937 20131 12940
rect 20073 12931 20131 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 22002 12968 22008 12980
rect 21963 12940 22008 12968
rect 22002 12928 22008 12940
rect 22060 12928 22066 12980
rect 22462 12968 22468 12980
rect 22423 12940 22468 12968
rect 22462 12928 22468 12940
rect 22520 12968 22526 12980
rect 24854 12968 24860 12980
rect 22520 12940 24860 12968
rect 22520 12928 22526 12940
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 26326 12968 26332 12980
rect 26287 12940 26332 12968
rect 26326 12928 26332 12940
rect 26384 12968 26390 12980
rect 27249 12971 27307 12977
rect 27249 12968 27261 12971
rect 26384 12940 27261 12968
rect 26384 12928 26390 12940
rect 27249 12937 27261 12940
rect 27295 12937 27307 12971
rect 27706 12968 27712 12980
rect 27667 12940 27712 12968
rect 27249 12931 27307 12937
rect 27706 12928 27712 12940
rect 27764 12928 27770 12980
rect 36538 12968 36544 12980
rect 31726 12940 36544 12968
rect 12437 12903 12495 12909
rect 12437 12869 12449 12903
rect 12483 12900 12495 12903
rect 12710 12900 12716 12912
rect 12483 12872 12716 12900
rect 12483 12869 12495 12872
rect 12437 12863 12495 12869
rect 12710 12860 12716 12872
rect 12768 12900 12774 12912
rect 13814 12900 13820 12912
rect 12768 12872 13820 12900
rect 12768 12860 12774 12872
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 15746 12900 15752 12912
rect 14292 12872 15752 12900
rect 10410 12832 10416 12844
rect 10371 12804 10416 12832
rect 10410 12792 10416 12804
rect 10468 12792 10474 12844
rect 10594 12832 10600 12844
rect 10555 12804 10600 12832
rect 10594 12792 10600 12804
rect 10652 12792 10658 12844
rect 11698 12832 11704 12844
rect 11659 12804 11704 12832
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12832 13691 12835
rect 14090 12832 14096 12844
rect 13679 12804 14096 12832
rect 13679 12801 13691 12804
rect 13633 12795 13691 12801
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14292 12841 14320 12872
rect 15746 12860 15752 12872
rect 15804 12860 15810 12912
rect 17862 12860 17868 12912
rect 17920 12900 17926 12912
rect 17957 12903 18015 12909
rect 17957 12900 17969 12903
rect 17920 12872 17969 12900
rect 17920 12860 17926 12872
rect 17957 12869 17969 12872
rect 18003 12869 18015 12903
rect 17957 12863 18015 12869
rect 18598 12860 18604 12912
rect 18656 12900 18662 12912
rect 19061 12903 19119 12909
rect 19061 12900 19073 12903
rect 18656 12872 19073 12900
rect 18656 12860 18662 12872
rect 19061 12869 19073 12872
rect 19107 12900 19119 12903
rect 19150 12900 19156 12912
rect 19107 12872 19156 12900
rect 19107 12869 19119 12872
rect 19061 12863 19119 12869
rect 19150 12860 19156 12872
rect 19208 12860 19214 12912
rect 20625 12903 20683 12909
rect 20625 12900 20637 12903
rect 19812 12872 20637 12900
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12801 14335 12835
rect 15194 12832 15200 12844
rect 14277 12795 14335 12801
rect 14384 12804 15200 12832
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8720 12736 9045 12764
rect 8720 12724 8726 12736
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 14384 12764 14412 12804
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 15933 12835 15991 12841
rect 15933 12832 15945 12835
rect 15304 12804 15945 12832
rect 15304 12776 15332 12804
rect 15933 12801 15945 12804
rect 15979 12801 15991 12835
rect 15933 12795 15991 12801
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 18230 12832 18236 12844
rect 17267 12804 18236 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 18690 12792 18696 12844
rect 18748 12832 18754 12844
rect 18877 12835 18935 12841
rect 18877 12832 18889 12835
rect 18748 12804 18889 12832
rect 18748 12792 18754 12804
rect 18877 12801 18889 12804
rect 18923 12801 18935 12835
rect 18877 12795 18935 12801
rect 19334 12792 19340 12844
rect 19392 12832 19398 12844
rect 19521 12835 19579 12841
rect 19521 12832 19533 12835
rect 19392 12804 19533 12832
rect 19392 12792 19398 12804
rect 19521 12801 19533 12804
rect 19567 12801 19579 12835
rect 19521 12795 19579 12801
rect 15286 12764 15292 12776
rect 9723 12736 14412 12764
rect 15247 12736 15292 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 17770 12764 17776 12776
rect 15396 12736 17776 12764
rect 6963 12668 8432 12696
rect 10413 12699 10471 12705
rect 6963 12665 6975 12668
rect 6917 12659 6975 12665
rect 10413 12665 10425 12699
rect 10459 12696 10471 12699
rect 10459 12668 12434 12696
rect 10459 12665 10471 12668
rect 10413 12659 10471 12665
rect 7837 12631 7895 12637
rect 7837 12597 7849 12631
rect 7883 12628 7895 12631
rect 8478 12628 8484 12640
rect 7883 12600 8484 12628
rect 7883 12597 7895 12600
rect 7837 12591 7895 12597
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 8573 12631 8631 12637
rect 8573 12597 8585 12631
rect 8619 12628 8631 12631
rect 8662 12628 8668 12640
rect 8619 12600 8668 12628
rect 8619 12597 8631 12600
rect 8573 12591 8631 12597
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 12406 12628 12434 12668
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 13078 12696 13084 12708
rect 12676 12668 13084 12696
rect 12676 12656 12682 12668
rect 13078 12656 13084 12668
rect 13136 12656 13142 12708
rect 15396 12696 15424 12736
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 19536 12764 19564 12795
rect 19610 12792 19616 12844
rect 19668 12832 19674 12844
rect 19812 12841 19840 12872
rect 20625 12869 20637 12872
rect 20671 12869 20683 12903
rect 20625 12863 20683 12869
rect 25314 12860 25320 12912
rect 25372 12900 25378 12912
rect 26142 12900 26148 12912
rect 25372 12872 26148 12900
rect 25372 12860 25378 12872
rect 26142 12860 26148 12872
rect 26200 12900 26206 12912
rect 31726 12900 31754 12940
rect 36538 12928 36544 12940
rect 36596 12968 36602 12980
rect 40034 12968 40040 12980
rect 36596 12940 40040 12968
rect 36596 12928 36602 12940
rect 40034 12928 40040 12940
rect 40092 12928 40098 12980
rect 43346 12928 43352 12980
rect 43404 12968 43410 12980
rect 43714 12968 43720 12980
rect 43404 12940 43720 12968
rect 43404 12928 43410 12940
rect 43714 12928 43720 12940
rect 43772 12928 43778 12980
rect 48608 12940 49372 12968
rect 26200 12872 31754 12900
rect 32677 12903 32735 12909
rect 26200 12860 26206 12872
rect 32677 12869 32689 12903
rect 32723 12900 32735 12903
rect 33318 12900 33324 12912
rect 32723 12872 33324 12900
rect 32723 12869 32735 12872
rect 32677 12863 32735 12869
rect 33318 12860 33324 12872
rect 33376 12900 33382 12912
rect 33505 12903 33563 12909
rect 33505 12900 33517 12903
rect 33376 12872 33517 12900
rect 33376 12860 33382 12872
rect 33505 12869 33517 12872
rect 33551 12900 33563 12903
rect 33778 12900 33784 12912
rect 33551 12872 33784 12900
rect 33551 12869 33563 12872
rect 33505 12863 33563 12869
rect 33778 12860 33784 12872
rect 33836 12860 33842 12912
rect 35526 12860 35532 12912
rect 35584 12900 35590 12912
rect 35621 12903 35679 12909
rect 35621 12900 35633 12903
rect 35584 12872 35633 12900
rect 35584 12860 35590 12872
rect 35621 12869 35633 12872
rect 35667 12900 35679 12903
rect 36354 12900 36360 12912
rect 35667 12872 36360 12900
rect 35667 12869 35679 12872
rect 35621 12863 35679 12869
rect 36354 12860 36360 12872
rect 36412 12860 36418 12912
rect 38470 12860 38476 12912
rect 38528 12900 38534 12912
rect 39485 12903 39543 12909
rect 39485 12900 39497 12903
rect 38528 12872 39497 12900
rect 38528 12860 38534 12872
rect 39485 12869 39497 12872
rect 39531 12869 39543 12903
rect 39485 12863 39543 12869
rect 41230 12860 41236 12912
rect 41288 12900 41294 12912
rect 44358 12900 44364 12912
rect 41288 12872 44364 12900
rect 41288 12860 41294 12872
rect 44358 12860 44364 12872
rect 44416 12860 44422 12912
rect 48608 12844 48636 12940
rect 48777 12903 48835 12909
rect 48777 12869 48789 12903
rect 48823 12900 48835 12903
rect 48958 12900 48964 12912
rect 48823 12872 48964 12900
rect 48823 12869 48835 12872
rect 48777 12863 48835 12869
rect 48958 12860 48964 12872
rect 49016 12860 49022 12912
rect 19797 12835 19855 12841
rect 19668 12804 19713 12832
rect 19668 12792 19674 12804
rect 19797 12801 19809 12835
rect 19843 12801 19855 12835
rect 19797 12795 19855 12801
rect 19889 12835 19947 12841
rect 19889 12801 19901 12835
rect 19935 12832 19947 12835
rect 20346 12832 20352 12844
rect 19935 12804 20352 12832
rect 19935 12801 19947 12804
rect 19889 12795 19947 12801
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 20714 12832 20720 12844
rect 20675 12804 20720 12832
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 21910 12792 21916 12844
rect 21968 12832 21974 12844
rect 22373 12835 22431 12841
rect 22373 12832 22385 12835
rect 21968 12804 22385 12832
rect 21968 12792 21974 12804
rect 22373 12801 22385 12804
rect 22419 12801 22431 12835
rect 22373 12795 22431 12801
rect 25501 12835 25559 12841
rect 25501 12801 25513 12835
rect 25547 12832 25559 12835
rect 26234 12832 26240 12844
rect 25547 12804 26240 12832
rect 25547 12801 25559 12804
rect 25501 12795 25559 12801
rect 26234 12792 26240 12804
rect 26292 12832 26298 12844
rect 26418 12832 26424 12844
rect 26292 12804 26424 12832
rect 26292 12792 26298 12804
rect 26418 12792 26424 12804
rect 26476 12792 26482 12844
rect 26510 12792 26516 12844
rect 26568 12832 26574 12844
rect 27341 12835 27399 12841
rect 27341 12832 27353 12835
rect 26568 12804 27353 12832
rect 26568 12792 26574 12804
rect 27341 12801 27353 12804
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 28353 12835 28411 12841
rect 28353 12801 28365 12835
rect 28399 12832 28411 12835
rect 33410 12832 33416 12844
rect 28399 12804 33416 12832
rect 28399 12801 28411 12804
rect 28353 12795 28411 12801
rect 33410 12792 33416 12804
rect 33468 12792 33474 12844
rect 37829 12835 37887 12841
rect 37829 12801 37841 12835
rect 37875 12832 37887 12835
rect 38562 12832 38568 12844
rect 37875 12804 38568 12832
rect 37875 12801 37887 12804
rect 37829 12795 37887 12801
rect 38562 12792 38568 12804
rect 38620 12792 38626 12844
rect 38746 12832 38752 12844
rect 38707 12804 38752 12832
rect 38746 12792 38752 12804
rect 38804 12792 38810 12844
rect 40310 12832 40316 12844
rect 40271 12804 40316 12832
rect 40310 12792 40316 12804
rect 40368 12792 40374 12844
rect 43257 12835 43315 12841
rect 43257 12801 43269 12835
rect 43303 12832 43315 12835
rect 43622 12832 43628 12844
rect 43303 12804 43628 12832
rect 43303 12801 43315 12804
rect 43257 12795 43315 12801
rect 43622 12792 43628 12804
rect 43680 12792 43686 12844
rect 48590 12832 48596 12844
rect 48551 12804 48596 12832
rect 48590 12792 48596 12804
rect 48648 12792 48654 12844
rect 49344 12841 49372 12940
rect 48869 12835 48927 12841
rect 48869 12801 48881 12835
rect 48915 12832 48927 12835
rect 49329 12835 49387 12841
rect 48915 12804 49280 12832
rect 48915 12801 48927 12804
rect 48869 12795 48927 12801
rect 20162 12764 20168 12776
rect 19536 12736 20168 12764
rect 20162 12724 20168 12736
rect 20220 12724 20226 12776
rect 22646 12764 22652 12776
rect 22607 12736 22652 12764
rect 22646 12724 22652 12736
rect 22704 12764 22710 12776
rect 23106 12764 23112 12776
rect 22704 12736 23112 12764
rect 22704 12724 22710 12736
rect 23106 12724 23112 12736
rect 23164 12724 23170 12776
rect 24854 12724 24860 12776
rect 24912 12764 24918 12776
rect 25409 12767 25467 12773
rect 25409 12764 25421 12767
rect 24912 12736 25421 12764
rect 24912 12724 24918 12736
rect 25409 12733 25421 12736
rect 25455 12764 25467 12767
rect 25590 12764 25596 12776
rect 25455 12736 25596 12764
rect 25455 12733 25467 12736
rect 25409 12727 25467 12733
rect 25590 12724 25596 12736
rect 25648 12724 25654 12776
rect 27062 12764 27068 12776
rect 27023 12736 27068 12764
rect 27062 12724 27068 12736
rect 27120 12724 27126 12776
rect 28261 12767 28319 12773
rect 28261 12733 28273 12767
rect 28307 12733 28319 12767
rect 33594 12764 33600 12776
rect 33555 12736 33600 12764
rect 28261 12727 28319 12733
rect 13188 12668 15424 12696
rect 13188 12628 13216 12668
rect 16390 12656 16396 12708
rect 16448 12696 16454 12708
rect 25682 12696 25688 12708
rect 16448 12668 25688 12696
rect 16448 12656 16454 12668
rect 25682 12656 25688 12668
rect 25740 12656 25746 12708
rect 25869 12699 25927 12705
rect 25869 12665 25881 12699
rect 25915 12696 25927 12699
rect 27430 12696 27436 12708
rect 25915 12668 27436 12696
rect 25915 12665 25927 12668
rect 25869 12659 25927 12665
rect 27430 12656 27436 12668
rect 27488 12696 27494 12708
rect 28276 12696 28304 12727
rect 33594 12724 33600 12736
rect 33652 12724 33658 12776
rect 33686 12724 33692 12776
rect 33744 12764 33750 12776
rect 33781 12767 33839 12773
rect 33781 12764 33793 12767
rect 33744 12736 33793 12764
rect 33744 12724 33750 12736
rect 33781 12733 33793 12736
rect 33827 12764 33839 12767
rect 33870 12764 33876 12776
rect 33827 12736 33876 12764
rect 33827 12733 33839 12736
rect 33781 12727 33839 12733
rect 33870 12724 33876 12736
rect 33928 12724 33934 12776
rect 49252 12764 49280 12804
rect 49329 12801 49341 12835
rect 49375 12801 49387 12835
rect 49329 12795 49387 12801
rect 49418 12764 49424 12776
rect 49252 12736 49424 12764
rect 49418 12724 49424 12736
rect 49476 12724 49482 12776
rect 27488 12668 28304 12696
rect 28721 12699 28779 12705
rect 27488 12656 27494 12668
rect 28721 12665 28733 12699
rect 28767 12696 28779 12699
rect 28810 12696 28816 12708
rect 28767 12668 28816 12696
rect 28767 12665 28779 12668
rect 28721 12659 28779 12665
rect 28810 12656 28816 12668
rect 28868 12656 28874 12708
rect 14918 12628 14924 12640
rect 12406 12600 13216 12628
rect 14879 12600 14924 12628
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 16025 12631 16083 12637
rect 16025 12597 16037 12631
rect 16071 12628 16083 12631
rect 16298 12628 16304 12640
rect 16071 12600 16304 12628
rect 16071 12597 16083 12600
rect 16025 12591 16083 12597
rect 16298 12588 16304 12600
rect 16356 12588 16362 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 19610 12628 19616 12640
rect 19392 12600 19616 12628
rect 19392 12588 19398 12600
rect 19610 12588 19616 12600
rect 19668 12628 19674 12640
rect 20438 12628 20444 12640
rect 19668 12600 20444 12628
rect 19668 12588 19674 12600
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 21266 12628 21272 12640
rect 21227 12600 21272 12628
rect 21266 12588 21272 12600
rect 21324 12588 21330 12640
rect 24857 12631 24915 12637
rect 24857 12597 24869 12631
rect 24903 12628 24915 12631
rect 24946 12628 24952 12640
rect 24903 12600 24952 12628
rect 24903 12597 24915 12600
rect 24857 12591 24915 12597
rect 24946 12588 24952 12600
rect 25004 12588 25010 12640
rect 33134 12628 33140 12640
rect 33095 12600 33140 12628
rect 33134 12588 33140 12600
rect 33192 12588 33198 12640
rect 37734 12628 37740 12640
rect 37695 12600 37740 12628
rect 37734 12588 37740 12600
rect 37792 12588 37798 12640
rect 38194 12588 38200 12640
rect 38252 12628 38258 12640
rect 40129 12631 40187 12637
rect 40129 12628 40141 12631
rect 38252 12600 40141 12628
rect 38252 12588 38258 12600
rect 40129 12597 40141 12600
rect 40175 12597 40187 12631
rect 40129 12591 40187 12597
rect 48593 12631 48651 12637
rect 48593 12597 48605 12631
rect 48639 12628 48651 12631
rect 49050 12628 49056 12640
rect 48639 12600 49056 12628
rect 48639 12597 48651 12600
rect 48593 12591 48651 12597
rect 49050 12588 49056 12600
rect 49108 12588 49114 12640
rect 49421 12631 49479 12637
rect 49421 12597 49433 12631
rect 49467 12628 49479 12631
rect 50154 12628 50160 12640
rect 49467 12600 50160 12628
rect 49467 12597 49479 12600
rect 49421 12591 49479 12597
rect 50154 12588 50160 12600
rect 50212 12588 50218 12640
rect 1104 12538 68816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 65654 12538
rect 65706 12486 65718 12538
rect 65770 12486 65782 12538
rect 65834 12486 65846 12538
rect 65898 12486 65910 12538
rect 65962 12486 68816 12538
rect 1104 12464 68816 12486
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8662 12424 8668 12436
rect 8352 12396 8668 12424
rect 8352 12384 8358 12396
rect 8662 12384 8668 12396
rect 8720 12384 8726 12436
rect 9585 12427 9643 12433
rect 9585 12393 9597 12427
rect 9631 12424 9643 12427
rect 10410 12424 10416 12436
rect 9631 12396 10416 12424
rect 9631 12393 9643 12396
rect 9585 12387 9643 12393
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 12710 12424 12716 12436
rect 12671 12396 12716 12424
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 12802 12384 12808 12436
rect 12860 12424 12866 12436
rect 13357 12427 13415 12433
rect 13357 12424 13369 12427
rect 12860 12396 13369 12424
rect 12860 12384 12866 12396
rect 13357 12393 13369 12396
rect 13403 12393 13415 12427
rect 13357 12387 13415 12393
rect 16022 12384 16028 12436
rect 16080 12424 16086 12436
rect 16117 12427 16175 12433
rect 16117 12424 16129 12427
rect 16080 12396 16129 12424
rect 16080 12384 16086 12396
rect 16117 12393 16129 12396
rect 16163 12393 16175 12427
rect 19978 12424 19984 12436
rect 19939 12396 19984 12424
rect 16117 12387 16175 12393
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20162 12424 20168 12436
rect 20123 12396 20168 12424
rect 20162 12384 20168 12396
rect 20220 12384 20226 12436
rect 20898 12384 20904 12436
rect 20956 12424 20962 12436
rect 20993 12427 21051 12433
rect 20993 12424 21005 12427
rect 20956 12396 21005 12424
rect 20956 12384 20962 12396
rect 20993 12393 21005 12396
rect 21039 12393 21051 12427
rect 20993 12387 21051 12393
rect 21082 12384 21088 12436
rect 21140 12424 21146 12436
rect 21910 12424 21916 12436
rect 21140 12396 21916 12424
rect 21140 12384 21146 12396
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 26973 12427 27031 12433
rect 26973 12393 26985 12427
rect 27019 12424 27031 12427
rect 29270 12424 29276 12436
rect 27019 12396 29276 12424
rect 27019 12393 27031 12396
rect 26973 12387 27031 12393
rect 29270 12384 29276 12396
rect 29328 12384 29334 12436
rect 37734 12424 37740 12436
rect 36188 12396 37740 12424
rect 7926 12316 7932 12368
rect 7984 12356 7990 12368
rect 8205 12359 8263 12365
rect 8205 12356 8217 12359
rect 7984 12328 8217 12356
rect 7984 12316 7990 12328
rect 8205 12325 8217 12328
rect 8251 12325 8263 12359
rect 8205 12319 8263 12325
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 15565 12359 15623 12365
rect 15565 12356 15577 12359
rect 15252 12328 15577 12356
rect 15252 12316 15258 12328
rect 15565 12325 15577 12328
rect 15611 12356 15623 12359
rect 16390 12356 16396 12368
rect 15611 12328 16396 12356
rect 15611 12325 15623 12328
rect 15565 12319 15623 12325
rect 16390 12316 16396 12328
rect 16448 12316 16454 12368
rect 21726 12356 21732 12368
rect 17696 12328 21732 12356
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 4893 12291 4951 12297
rect 4893 12288 4905 12291
rect 4764 12260 4905 12288
rect 4764 12248 4770 12260
rect 4893 12257 4905 12260
rect 4939 12257 4951 12291
rect 7374 12288 7380 12300
rect 7335 12260 7380 12288
rect 4893 12251 4951 12257
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 9306 12288 9312 12300
rect 9267 12260 9312 12288
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 17696 12288 17724 12328
rect 21726 12316 21732 12328
rect 21784 12316 21790 12368
rect 16408 12260 17724 12288
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 5684 12192 7236 12220
rect 5684 12180 5690 12192
rect 5160 12155 5218 12161
rect 5160 12121 5172 12155
rect 5206 12152 5218 12155
rect 5258 12152 5264 12164
rect 5206 12124 5264 12152
rect 5206 12121 5218 12124
rect 5160 12115 5218 12121
rect 5258 12112 5264 12124
rect 5316 12112 5322 12164
rect 7098 12152 7104 12164
rect 6288 12124 7104 12152
rect 6288 12093 6316 12124
rect 7098 12112 7104 12124
rect 7156 12112 7162 12164
rect 6273 12087 6331 12093
rect 6273 12053 6285 12087
rect 6319 12053 6331 12087
rect 6730 12084 6736 12096
rect 6691 12056 6736 12084
rect 6273 12047 6331 12053
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 7208 12093 7236 12192
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 9585 12223 9643 12229
rect 9585 12220 9597 12223
rect 8720 12192 9597 12220
rect 8720 12180 8726 12192
rect 9585 12189 9597 12192
rect 9631 12189 9643 12223
rect 9585 12183 9643 12189
rect 9677 12223 9735 12229
rect 9677 12189 9689 12223
rect 9723 12220 9735 12223
rect 10410 12220 10416 12232
rect 9723 12192 10416 12220
rect 9723 12189 9735 12192
rect 9677 12183 9735 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12220 12219 12223
rect 12250 12220 12256 12232
rect 12207 12192 12256 12220
rect 12207 12189 12219 12192
rect 12161 12183 12219 12189
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 16298 12229 16304 12232
rect 16296 12220 16304 12229
rect 16259 12192 16304 12220
rect 16296 12183 16304 12192
rect 16298 12180 16304 12183
rect 16356 12180 16362 12232
rect 16408 12229 16436 12260
rect 17770 12248 17776 12300
rect 17828 12288 17834 12300
rect 35437 12291 35495 12297
rect 35437 12288 35449 12291
rect 17828 12260 35449 12288
rect 17828 12248 17834 12260
rect 35437 12257 35449 12260
rect 35483 12288 35495 12291
rect 36078 12288 36084 12300
rect 35483 12260 36084 12288
rect 35483 12257 35495 12260
rect 35437 12251 35495 12257
rect 36078 12248 36084 12260
rect 36136 12248 36142 12300
rect 36188 12297 36216 12396
rect 37734 12384 37740 12396
rect 37792 12384 37798 12436
rect 38746 12384 38752 12436
rect 38804 12424 38810 12436
rect 39853 12427 39911 12433
rect 39853 12424 39865 12427
rect 38804 12396 39865 12424
rect 38804 12384 38810 12396
rect 39853 12393 39865 12396
rect 39899 12393 39911 12427
rect 39853 12387 39911 12393
rect 48225 12427 48283 12433
rect 48225 12393 48237 12427
rect 48271 12424 48283 12427
rect 48271 12396 48820 12424
rect 48271 12393 48283 12396
rect 48225 12387 48283 12393
rect 38841 12359 38899 12365
rect 38841 12325 38853 12359
rect 38887 12356 38899 12359
rect 40310 12356 40316 12368
rect 38887 12328 40316 12356
rect 38887 12325 38899 12328
rect 38841 12319 38899 12325
rect 40310 12316 40316 12328
rect 40368 12316 40374 12368
rect 47946 12316 47952 12368
rect 48004 12356 48010 12368
rect 48685 12359 48743 12365
rect 48685 12356 48697 12359
rect 48004 12328 48697 12356
rect 48004 12316 48010 12328
rect 48685 12325 48697 12328
rect 48731 12325 48743 12359
rect 48792 12356 48820 12396
rect 48866 12384 48872 12436
rect 48924 12424 48930 12436
rect 48924 12396 48969 12424
rect 48924 12384 48930 12396
rect 48958 12356 48964 12368
rect 48792 12328 48964 12356
rect 48685 12319 48743 12325
rect 48958 12316 48964 12328
rect 49016 12316 49022 12368
rect 36173 12291 36231 12297
rect 36173 12257 36185 12291
rect 36219 12257 36231 12291
rect 36354 12288 36360 12300
rect 36315 12260 36360 12288
rect 36173 12251 36231 12257
rect 36354 12248 36360 12260
rect 36412 12248 36418 12300
rect 16393 12223 16451 12229
rect 16393 12189 16405 12223
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 16574 12180 16580 12232
rect 16632 12229 16638 12232
rect 16632 12223 16671 12229
rect 16659 12189 16671 12223
rect 16632 12183 16671 12189
rect 16632 12180 16638 12183
rect 16758 12180 16764 12232
rect 16816 12220 16822 12232
rect 19426 12220 19432 12232
rect 16816 12192 16861 12220
rect 19387 12192 19432 12220
rect 16816 12180 16822 12192
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12189 20223 12223
rect 20165 12183 20223 12189
rect 20257 12223 20315 12229
rect 20257 12189 20269 12223
rect 20303 12220 20315 12223
rect 20898 12220 20904 12232
rect 20303 12192 20904 12220
rect 20303 12189 20315 12192
rect 20257 12183 20315 12189
rect 7929 12155 7987 12161
rect 7929 12121 7941 12155
rect 7975 12152 7987 12155
rect 8570 12152 8576 12164
rect 7975 12124 8576 12152
rect 7975 12121 7987 12124
rect 7929 12115 7987 12121
rect 8570 12112 8576 12124
rect 8628 12112 8634 12164
rect 14553 12155 14611 12161
rect 14553 12121 14565 12155
rect 14599 12152 14611 12155
rect 15010 12152 15016 12164
rect 14599 12124 15016 12152
rect 14599 12121 14611 12124
rect 14553 12115 14611 12121
rect 15010 12112 15016 12124
rect 15068 12152 15074 12164
rect 15286 12152 15292 12164
rect 15068 12124 15292 12152
rect 15068 12112 15074 12124
rect 15286 12112 15292 12124
rect 15344 12112 15350 12164
rect 16485 12155 16543 12161
rect 16485 12121 16497 12155
rect 16531 12152 16543 12155
rect 20180 12152 20208 12183
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 21085 12223 21143 12229
rect 21085 12189 21097 12223
rect 21131 12220 21143 12223
rect 21266 12220 21272 12232
rect 21131 12192 21272 12220
rect 21131 12189 21143 12192
rect 21085 12183 21143 12189
rect 21266 12180 21272 12192
rect 21324 12220 21330 12232
rect 23474 12220 23480 12232
rect 21324 12192 23480 12220
rect 21324 12180 21330 12192
rect 23474 12180 23480 12192
rect 23532 12180 23538 12232
rect 23750 12180 23756 12232
rect 23808 12220 23814 12232
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 23808 12192 24593 12220
rect 23808 12180 23814 12192
rect 24581 12189 24593 12192
rect 24627 12220 24639 12223
rect 24670 12220 24676 12232
rect 24627 12192 24676 12220
rect 24627 12189 24639 12192
rect 24581 12183 24639 12189
rect 24670 12180 24676 12192
rect 24728 12180 24734 12232
rect 25222 12220 25228 12232
rect 25183 12192 25228 12220
rect 25222 12180 25228 12192
rect 25280 12180 25286 12232
rect 25590 12220 25596 12232
rect 25551 12192 25596 12220
rect 25590 12180 25596 12192
rect 25648 12180 25654 12232
rect 26142 12220 26148 12232
rect 26103 12192 26148 12220
rect 26142 12180 26148 12192
rect 26200 12180 26206 12232
rect 26602 12220 26608 12232
rect 26563 12192 26608 12220
rect 26602 12180 26608 12192
rect 26660 12180 26666 12232
rect 26786 12180 26792 12232
rect 26844 12220 26850 12232
rect 26844 12192 26889 12220
rect 26844 12180 26850 12192
rect 31294 12180 31300 12232
rect 31352 12220 31358 12232
rect 31481 12223 31539 12229
rect 31481 12220 31493 12223
rect 31352 12192 31493 12220
rect 31352 12180 31358 12192
rect 31481 12189 31493 12192
rect 31527 12189 31539 12223
rect 31481 12183 31539 12189
rect 36265 12223 36323 12229
rect 36265 12189 36277 12223
rect 36311 12220 36323 12223
rect 36906 12220 36912 12232
rect 36311 12192 36912 12220
rect 36311 12189 36323 12192
rect 36265 12183 36323 12189
rect 36906 12180 36912 12192
rect 36964 12180 36970 12232
rect 37001 12223 37059 12229
rect 37001 12189 37013 12223
rect 37047 12220 37059 12223
rect 37182 12220 37188 12232
rect 37047 12192 37188 12220
rect 37047 12189 37059 12192
rect 37001 12183 37059 12189
rect 37182 12180 37188 12192
rect 37240 12180 37246 12232
rect 37277 12223 37335 12229
rect 37277 12189 37289 12223
rect 37323 12189 37335 12223
rect 37277 12183 37335 12189
rect 20438 12152 20444 12164
rect 16531 12124 16712 12152
rect 20180 12124 20300 12152
rect 20399 12124 20444 12152
rect 16531 12121 16543 12124
rect 16485 12115 16543 12121
rect 16684 12096 16712 12124
rect 7193 12087 7251 12093
rect 7193 12053 7205 12087
rect 7239 12084 7251 12087
rect 7282 12084 7288 12096
rect 7239 12056 7288 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 8389 12087 8447 12093
rect 8389 12053 8401 12087
rect 8435 12084 8447 12087
rect 8754 12084 8760 12096
rect 8435 12056 8760 12084
rect 8435 12053 8447 12056
rect 8389 12047 8447 12053
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 9490 12084 9496 12096
rect 9451 12056 9496 12084
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 11054 12084 11060 12096
rect 11015 12056 11060 12084
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 11974 12084 11980 12096
rect 11935 12056 11980 12084
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 14645 12087 14703 12093
rect 14645 12053 14657 12087
rect 14691 12084 14703 12087
rect 14826 12084 14832 12096
rect 14691 12056 14832 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 16666 12044 16672 12096
rect 16724 12044 16730 12096
rect 18690 12084 18696 12096
rect 18651 12056 18696 12084
rect 18690 12044 18696 12056
rect 18748 12044 18754 12096
rect 19242 12084 19248 12096
rect 19203 12056 19248 12084
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 20272 12084 20300 12124
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 32030 12112 32036 12164
rect 32088 12152 32094 12164
rect 32125 12155 32183 12161
rect 32125 12152 32137 12155
rect 32088 12124 32137 12152
rect 32088 12112 32094 12124
rect 32125 12121 32137 12124
rect 32171 12121 32183 12155
rect 32125 12115 32183 12121
rect 20622 12084 20628 12096
rect 20272 12056 20628 12084
rect 20622 12044 20628 12056
rect 20680 12084 20686 12096
rect 20990 12084 20996 12096
rect 20680 12056 20996 12084
rect 20680 12044 20686 12056
rect 20990 12044 20996 12056
rect 21048 12044 21054 12096
rect 24394 12044 24400 12096
rect 24452 12084 24458 12096
rect 24489 12087 24547 12093
rect 24489 12084 24501 12087
rect 24452 12056 24501 12084
rect 24452 12044 24458 12056
rect 24489 12053 24501 12056
rect 24535 12053 24547 12087
rect 31662 12084 31668 12096
rect 31623 12056 31668 12084
rect 24489 12047 24547 12053
rect 31662 12044 31668 12056
rect 31720 12044 31726 12096
rect 32140 12084 32168 12115
rect 32858 12112 32864 12164
rect 32916 12152 32922 12164
rect 32953 12155 33011 12161
rect 32953 12152 32965 12155
rect 32916 12124 32965 12152
rect 32916 12112 32922 12124
rect 32953 12121 32965 12124
rect 32999 12152 33011 12155
rect 33042 12152 33048 12164
rect 32999 12124 33048 12152
rect 32999 12121 33011 12124
rect 32953 12115 33011 12121
rect 33042 12112 33048 12124
rect 33100 12112 33106 12164
rect 37292 12152 37320 12183
rect 37366 12180 37372 12232
rect 37424 12220 37430 12232
rect 38194 12220 38200 12232
rect 37424 12192 38200 12220
rect 37424 12180 37430 12192
rect 38194 12180 38200 12192
rect 38252 12180 38258 12232
rect 38562 12220 38568 12232
rect 38523 12192 38568 12220
rect 38562 12180 38568 12192
rect 38620 12180 38626 12232
rect 38657 12223 38715 12229
rect 38657 12189 38669 12223
rect 38703 12189 38715 12223
rect 38657 12183 38715 12189
rect 38672 12152 38700 12183
rect 40126 12180 40132 12232
rect 40184 12220 40190 12232
rect 40497 12223 40555 12229
rect 40497 12220 40509 12223
rect 40184 12192 40509 12220
rect 40184 12180 40190 12192
rect 40497 12189 40509 12192
rect 40543 12220 40555 12223
rect 40957 12223 41015 12229
rect 40957 12220 40969 12223
rect 40543 12192 40969 12220
rect 40543 12189 40555 12192
rect 40497 12183 40555 12189
rect 40957 12189 40969 12192
rect 41003 12220 41015 12223
rect 43714 12220 43720 12232
rect 41003 12192 43720 12220
rect 41003 12189 41015 12192
rect 40957 12183 41015 12189
rect 43714 12180 43720 12192
rect 43772 12180 43778 12232
rect 44266 12180 44272 12232
rect 44324 12220 44330 12232
rect 45189 12223 45247 12229
rect 45189 12220 45201 12223
rect 44324 12192 45201 12220
rect 44324 12180 44330 12192
rect 45189 12189 45201 12192
rect 45235 12220 45247 12223
rect 45462 12220 45468 12232
rect 45235 12192 45468 12220
rect 45235 12189 45247 12192
rect 45189 12183 45247 12189
rect 45462 12180 45468 12192
rect 45520 12180 45526 12232
rect 48038 12220 48044 12232
rect 47999 12192 48044 12220
rect 48038 12180 48044 12192
rect 48096 12180 48102 12232
rect 36556 12124 37320 12152
rect 37936 12124 38700 12152
rect 33597 12087 33655 12093
rect 33597 12084 33609 12087
rect 32140 12056 33609 12084
rect 33597 12053 33609 12056
rect 33643 12084 33655 12087
rect 33962 12084 33968 12096
rect 33643 12056 33968 12084
rect 33643 12053 33655 12056
rect 33597 12047 33655 12053
rect 33962 12044 33968 12056
rect 34020 12044 34026 12096
rect 36556 12093 36584 12124
rect 36541 12087 36599 12093
rect 36541 12053 36553 12087
rect 36587 12053 36599 12087
rect 36541 12047 36599 12053
rect 36906 12044 36912 12096
rect 36964 12084 36970 12096
rect 37936 12084 37964 12124
rect 48130 12112 48136 12164
rect 48188 12152 48194 12164
rect 48837 12155 48895 12161
rect 48837 12152 48849 12155
rect 48188 12124 48849 12152
rect 48188 12112 48194 12124
rect 48837 12121 48849 12124
rect 48883 12121 48895 12155
rect 49050 12152 49056 12164
rect 49011 12124 49056 12152
rect 48837 12115 48895 12121
rect 49050 12112 49056 12124
rect 49108 12112 49114 12164
rect 36964 12056 37964 12084
rect 38013 12087 38071 12093
rect 36964 12044 36970 12056
rect 38013 12053 38025 12087
rect 38059 12084 38071 12087
rect 38286 12084 38292 12096
rect 38059 12056 38292 12084
rect 38059 12053 38071 12056
rect 38013 12047 38071 12053
rect 38286 12044 38292 12056
rect 38344 12044 38350 12096
rect 40678 12044 40684 12096
rect 40736 12084 40742 12096
rect 41141 12087 41199 12093
rect 41141 12084 41153 12087
rect 40736 12056 41153 12084
rect 40736 12044 40742 12056
rect 41141 12053 41153 12056
rect 41187 12084 41199 12087
rect 41322 12084 41328 12096
rect 41187 12056 41328 12084
rect 41187 12053 41199 12056
rect 41141 12047 41199 12053
rect 41322 12044 41328 12056
rect 41380 12044 41386 12096
rect 45094 12084 45100 12096
rect 45055 12056 45100 12084
rect 45094 12044 45100 12056
rect 45152 12044 45158 12096
rect 45554 12044 45560 12096
rect 45612 12084 45618 12096
rect 46842 12084 46848 12096
rect 45612 12056 46848 12084
rect 45612 12044 45618 12056
rect 46842 12044 46848 12056
rect 46900 12084 46906 12096
rect 48314 12084 48320 12096
rect 46900 12056 48320 12084
rect 46900 12044 46906 12056
rect 48314 12044 48320 12056
rect 48372 12044 48378 12096
rect 1104 11994 68816 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 68816 11994
rect 1104 11920 68816 11942
rect 5258 11880 5264 11892
rect 5219 11852 5264 11880
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 8297 11883 8355 11889
rect 8297 11880 8309 11883
rect 8168 11852 8309 11880
rect 8168 11840 8174 11852
rect 8297 11849 8309 11852
rect 8343 11849 8355 11883
rect 10410 11880 10416 11892
rect 10371 11852 10416 11880
rect 8297 11843 8355 11849
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 16669 11883 16727 11889
rect 16669 11849 16681 11883
rect 16715 11880 16727 11883
rect 16758 11880 16764 11892
rect 16715 11852 16764 11880
rect 16715 11849 16727 11852
rect 16669 11843 16727 11849
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 17954 11880 17960 11892
rect 17788 11852 17960 11880
rect 8386 11772 8392 11824
rect 8444 11812 8450 11824
rect 11876 11815 11934 11821
rect 8444 11784 8984 11812
rect 8444 11772 8450 11784
rect 5445 11747 5503 11753
rect 5445 11713 5457 11747
rect 5491 11744 5503 11747
rect 6730 11744 6736 11756
rect 5491 11716 6736 11744
rect 5491 11713 5503 11716
rect 5445 11707 5503 11713
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 7834 11744 7840 11756
rect 7795 11716 7840 11744
rect 7834 11704 7840 11716
rect 7892 11704 7898 11756
rect 8021 11747 8079 11753
rect 8021 11713 8033 11747
rect 8067 11744 8079 11747
rect 8294 11744 8300 11756
rect 8067 11716 8300 11744
rect 8067 11713 8079 11716
rect 8021 11707 8079 11713
rect 8294 11704 8300 11716
rect 8352 11704 8358 11756
rect 8754 11744 8760 11756
rect 8715 11716 8760 11744
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 8956 11753 8984 11784
rect 11876 11781 11888 11815
rect 11922 11812 11934 11815
rect 11974 11812 11980 11824
rect 11922 11784 11980 11812
rect 11922 11781 11934 11784
rect 11876 11775 11934 11781
rect 11974 11772 11980 11784
rect 12032 11772 12038 11824
rect 17788 11812 17816 11852
rect 17954 11840 17960 11852
rect 18012 11880 18018 11892
rect 18506 11880 18512 11892
rect 18012 11852 18512 11880
rect 18012 11840 18018 11852
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 20438 11880 20444 11892
rect 20399 11852 20444 11880
rect 20438 11840 20444 11852
rect 20496 11840 20502 11892
rect 24765 11883 24823 11889
rect 24765 11849 24777 11883
rect 24811 11880 24823 11883
rect 25314 11880 25320 11892
rect 24811 11852 25320 11880
rect 24811 11849 24823 11852
rect 24765 11843 24823 11849
rect 25314 11840 25320 11852
rect 25372 11840 25378 11892
rect 25409 11883 25467 11889
rect 25409 11849 25421 11883
rect 25455 11880 25467 11883
rect 26878 11880 26884 11892
rect 25455 11852 26884 11880
rect 25455 11849 25467 11852
rect 25409 11843 25467 11849
rect 26878 11840 26884 11852
rect 26936 11840 26942 11892
rect 32769 11883 32827 11889
rect 32769 11849 32781 11883
rect 32815 11849 32827 11883
rect 32769 11843 32827 11849
rect 12406 11784 17816 11812
rect 8941 11747 8999 11753
rect 8941 11713 8953 11747
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11744 10655 11747
rect 11238 11744 11244 11756
rect 10643 11716 11244 11744
rect 10643 11713 10655 11716
rect 10597 11707 10655 11713
rect 11238 11704 11244 11716
rect 11296 11744 11302 11756
rect 12406 11744 12434 11784
rect 17862 11772 17868 11824
rect 17920 11812 17926 11824
rect 17920 11784 23060 11812
rect 17920 11772 17926 11784
rect 14185 11747 14243 11753
rect 14185 11744 14197 11747
rect 11296 11716 12434 11744
rect 13004 11716 14197 11744
rect 11296 11704 11302 11716
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11645 7987 11679
rect 8110 11676 8116 11688
rect 8071 11648 8116 11676
rect 7929 11639 7987 11645
rect 7944 11608 7972 11639
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 10686 11676 10692 11688
rect 10647 11648 10692 11676
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 10781 11679 10839 11685
rect 10781 11645 10793 11679
rect 10827 11676 10839 11679
rect 11054 11676 11060 11688
rect 10827 11648 11060 11676
rect 10827 11645 10839 11648
rect 10781 11639 10839 11645
rect 11054 11636 11060 11648
rect 11112 11636 11118 11688
rect 11514 11636 11520 11688
rect 11572 11676 11578 11688
rect 11609 11679 11667 11685
rect 11609 11676 11621 11679
rect 11572 11648 11621 11676
rect 11572 11636 11578 11648
rect 11609 11645 11621 11648
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 7944 11580 8156 11608
rect 8128 11552 8156 11580
rect 12618 11568 12624 11620
rect 12676 11608 12682 11620
rect 13004 11617 13032 11716
rect 14185 11713 14197 11716
rect 14231 11713 14243 11747
rect 16850 11744 16856 11756
rect 16811 11716 16856 11744
rect 14185 11707 14243 11713
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 18616 11753 18644 11784
rect 18601 11747 18659 11753
rect 18601 11713 18613 11747
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 18868 11747 18926 11753
rect 18868 11713 18880 11747
rect 18914 11744 18926 11747
rect 19242 11744 19248 11756
rect 18914 11716 19248 11744
rect 18914 11713 18926 11716
rect 18868 11707 18926 11713
rect 19242 11704 19248 11716
rect 19300 11704 19306 11756
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11744 20775 11747
rect 20806 11744 20812 11756
rect 20763 11716 20812 11744
rect 20763 11713 20775 11716
rect 20717 11707 20775 11713
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 20990 11744 20996 11756
rect 20951 11716 20996 11744
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 23032 11753 23060 11784
rect 25222 11772 25228 11824
rect 25280 11812 25286 11824
rect 26329 11815 26387 11821
rect 26329 11812 26341 11815
rect 25280 11784 26341 11812
rect 25280 11772 25286 11784
rect 26329 11781 26341 11784
rect 26375 11781 26387 11815
rect 26329 11775 26387 11781
rect 30561 11815 30619 11821
rect 30561 11781 30573 11815
rect 30607 11812 30619 11815
rect 32122 11812 32128 11824
rect 30607 11784 32128 11812
rect 30607 11781 30619 11784
rect 30561 11775 30619 11781
rect 32122 11772 32128 11784
rect 32180 11772 32186 11824
rect 32784 11812 32812 11843
rect 37274 11840 37280 11892
rect 37332 11880 37338 11892
rect 37461 11883 37519 11889
rect 37461 11880 37473 11883
rect 37332 11852 37473 11880
rect 37332 11840 37338 11852
rect 37461 11849 37473 11852
rect 37507 11880 37519 11883
rect 37734 11880 37740 11892
rect 37507 11852 37740 11880
rect 37507 11849 37519 11852
rect 37461 11843 37519 11849
rect 37734 11840 37740 11852
rect 37792 11840 37798 11892
rect 38470 11880 38476 11892
rect 38028 11852 38476 11880
rect 33474 11815 33532 11821
rect 33474 11812 33486 11815
rect 32784 11784 33486 11812
rect 33474 11781 33486 11784
rect 33520 11781 33532 11815
rect 38028 11812 38056 11852
rect 38470 11840 38476 11852
rect 38528 11880 38534 11892
rect 41598 11880 41604 11892
rect 38528 11852 41604 11880
rect 38528 11840 38534 11852
rect 41598 11840 41604 11852
rect 41656 11840 41662 11892
rect 42150 11840 42156 11892
rect 42208 11880 42214 11892
rect 42521 11883 42579 11889
rect 42521 11880 42533 11883
rect 42208 11852 42533 11880
rect 42208 11840 42214 11852
rect 42521 11849 42533 11852
rect 42567 11880 42579 11883
rect 45554 11880 45560 11892
rect 42567 11852 45560 11880
rect 42567 11849 42579 11852
rect 42521 11843 42579 11849
rect 45554 11840 45560 11852
rect 45612 11840 45618 11892
rect 45649 11883 45707 11889
rect 45649 11849 45661 11883
rect 45695 11880 45707 11883
rect 48038 11880 48044 11892
rect 45695 11852 48044 11880
rect 45695 11849 45707 11852
rect 45649 11843 45707 11849
rect 48038 11840 48044 11852
rect 48096 11880 48102 11892
rect 49234 11880 49240 11892
rect 48096 11852 49240 11880
rect 48096 11840 48102 11852
rect 49234 11840 49240 11852
rect 49292 11840 49298 11892
rect 49694 11840 49700 11892
rect 49752 11880 49758 11892
rect 50801 11883 50859 11889
rect 50801 11880 50813 11883
rect 49752 11852 50813 11880
rect 49752 11840 49758 11852
rect 38286 11812 38292 11824
rect 33474 11775 33532 11781
rect 36464 11784 38056 11812
rect 38247 11784 38292 11812
rect 23017 11747 23075 11753
rect 23017 11713 23029 11747
rect 23063 11713 23075 11747
rect 23017 11707 23075 11713
rect 24394 11704 24400 11756
rect 24452 11704 24458 11756
rect 24946 11704 24952 11756
rect 25004 11744 25010 11756
rect 25593 11747 25651 11753
rect 25593 11744 25605 11747
rect 25004 11716 25605 11744
rect 25004 11704 25010 11716
rect 25593 11713 25605 11716
rect 25639 11713 25651 11747
rect 25593 11707 25651 11713
rect 26234 11704 26240 11756
rect 26292 11744 26298 11756
rect 26970 11744 26976 11756
rect 26292 11716 26337 11744
rect 26931 11716 26976 11744
rect 26292 11704 26298 11716
rect 26970 11704 26976 11716
rect 27028 11704 27034 11756
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11744 27215 11747
rect 27430 11744 27436 11756
rect 27203 11716 27436 11744
rect 27203 11713 27215 11716
rect 27157 11707 27215 11713
rect 27430 11704 27436 11716
rect 27488 11704 27494 11756
rect 28902 11744 28908 11756
rect 28863 11716 28908 11744
rect 28902 11704 28908 11716
rect 28960 11704 28966 11756
rect 30469 11747 30527 11753
rect 30469 11744 30481 11747
rect 29288 11716 30481 11744
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11645 14335 11679
rect 15654 11676 15660 11688
rect 15615 11648 15660 11676
rect 14277 11639 14335 11645
rect 12989 11611 13047 11617
rect 12989 11608 13001 11611
rect 12676 11580 13001 11608
rect 12676 11568 12682 11580
rect 12989 11577 13001 11580
rect 13035 11577 13047 11611
rect 14292 11608 14320 11639
rect 15654 11636 15660 11648
rect 15712 11636 15718 11688
rect 16298 11636 16304 11688
rect 16356 11676 16362 11688
rect 17037 11679 17095 11685
rect 17037 11676 17049 11679
rect 16356 11648 17049 11676
rect 16356 11636 16362 11648
rect 17037 11645 17049 11648
rect 17083 11645 17095 11679
rect 17037 11639 17095 11645
rect 17129 11679 17187 11685
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 17589 11679 17647 11685
rect 17589 11676 17601 11679
rect 17175 11648 17601 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 17589 11645 17601 11648
rect 17635 11645 17647 11679
rect 23290 11676 23296 11688
rect 23251 11648 23296 11676
rect 17589 11639 17647 11645
rect 14918 11608 14924 11620
rect 14292 11580 14924 11608
rect 12989 11571 13047 11577
rect 14918 11568 14924 11580
rect 14976 11608 14982 11620
rect 15933 11611 15991 11617
rect 15933 11608 15945 11611
rect 14976 11580 15945 11608
rect 14976 11568 14982 11580
rect 15933 11577 15945 11580
rect 15979 11577 15991 11611
rect 15933 11571 15991 11577
rect 7282 11540 7288 11552
rect 7243 11512 7288 11540
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 8941 11543 8999 11549
rect 8941 11540 8953 11543
rect 8168 11512 8953 11540
rect 8168 11500 8174 11512
rect 8941 11509 8953 11512
rect 8987 11540 8999 11543
rect 9490 11540 9496 11552
rect 8987 11512 9496 11540
rect 8987 11509 8999 11512
rect 8941 11503 8999 11509
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 14461 11543 14519 11549
rect 14461 11509 14473 11543
rect 14507 11540 14519 11543
rect 14734 11540 14740 11552
rect 14507 11512 14740 11540
rect 14507 11509 14519 11512
rect 14461 11503 14519 11509
rect 14734 11500 14740 11512
rect 14792 11500 14798 11552
rect 15105 11543 15163 11549
rect 15105 11509 15117 11543
rect 15151 11540 15163 11543
rect 15286 11540 15292 11552
rect 15151 11512 15292 11540
rect 15151 11509 15163 11512
rect 15105 11503 15163 11509
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 16117 11543 16175 11549
rect 16117 11509 16129 11543
rect 16163 11540 16175 11543
rect 16666 11540 16672 11552
rect 16163 11512 16672 11540
rect 16163 11509 16175 11512
rect 16117 11503 16175 11509
rect 16666 11500 16672 11512
rect 16724 11500 16730 11552
rect 17604 11540 17632 11639
rect 23290 11636 23296 11648
rect 23348 11636 23354 11688
rect 25038 11636 25044 11688
rect 25096 11676 25102 11688
rect 25225 11679 25283 11685
rect 25225 11676 25237 11679
rect 25096 11648 25237 11676
rect 25096 11636 25102 11648
rect 25225 11645 25237 11648
rect 25271 11645 25283 11679
rect 28810 11676 28816 11688
rect 28771 11648 28816 11676
rect 25225 11639 25283 11645
rect 28810 11636 28816 11648
rect 28868 11636 28874 11688
rect 25792 11580 26234 11608
rect 19794 11540 19800 11552
rect 17604 11512 19800 11540
rect 19794 11500 19800 11512
rect 19852 11500 19858 11552
rect 19978 11540 19984 11552
rect 19939 11512 19984 11540
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 20714 11540 20720 11552
rect 20675 11512 20720 11540
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 25792 11549 25820 11580
rect 25777 11543 25835 11549
rect 25777 11509 25789 11543
rect 25823 11509 25835 11543
rect 26206 11540 26234 11580
rect 26602 11568 26608 11620
rect 26660 11608 26666 11620
rect 27065 11611 27123 11617
rect 27065 11608 27077 11611
rect 26660 11580 27077 11608
rect 26660 11568 26666 11580
rect 27065 11577 27077 11580
rect 27111 11608 27123 11611
rect 28994 11608 29000 11620
rect 27111 11580 29000 11608
rect 27111 11577 27123 11580
rect 27065 11571 27123 11577
rect 28994 11568 29000 11580
rect 29052 11568 29058 11620
rect 29288 11617 29316 11716
rect 30469 11713 30481 11716
rect 30515 11713 30527 11747
rect 30650 11744 30656 11756
rect 30611 11716 30656 11744
rect 30469 11707 30527 11713
rect 30650 11704 30656 11716
rect 30708 11704 30714 11756
rect 30926 11744 30932 11756
rect 30887 11716 30932 11744
rect 30926 11704 30932 11716
rect 30984 11704 30990 11756
rect 31110 11744 31116 11756
rect 31071 11716 31116 11744
rect 31110 11704 31116 11716
rect 31168 11704 31174 11756
rect 31386 11744 31392 11756
rect 31347 11716 31392 11744
rect 31386 11704 31392 11716
rect 31444 11704 31450 11756
rect 32585 11747 32643 11753
rect 32585 11713 32597 11747
rect 32631 11744 32643 11747
rect 33134 11744 33140 11756
rect 32631 11716 33140 11744
rect 32631 11713 32643 11716
rect 32585 11707 32643 11713
rect 33134 11704 33140 11716
rect 33192 11704 33198 11756
rect 33778 11704 33784 11756
rect 33836 11744 33842 11756
rect 36464 11753 36492 11784
rect 38028 11753 38056 11784
rect 38286 11772 38292 11784
rect 38344 11772 38350 11824
rect 40313 11815 40371 11821
rect 40313 11812 40325 11815
rect 39514 11784 40325 11812
rect 40313 11781 40325 11784
rect 40359 11781 40371 11815
rect 46201 11815 46259 11821
rect 46201 11812 46213 11815
rect 45402 11784 46213 11812
rect 40313 11775 40371 11781
rect 46201 11781 46213 11784
rect 46247 11781 46259 11815
rect 46201 11775 46259 11781
rect 48130 11772 48136 11824
rect 48188 11812 48194 11824
rect 50172 11821 50200 11852
rect 50801 11849 50813 11852
rect 50847 11849 50859 11883
rect 50801 11843 50859 11849
rect 49973 11815 50031 11821
rect 49973 11812 49985 11815
rect 48188 11784 49985 11812
rect 48188 11772 48194 11784
rect 49973 11781 49985 11784
rect 50019 11781 50031 11815
rect 49973 11775 50031 11781
rect 50157 11815 50215 11821
rect 50157 11781 50169 11815
rect 50203 11781 50215 11815
rect 50157 11775 50215 11781
rect 36182 11747 36240 11753
rect 36182 11744 36194 11747
rect 33836 11716 36194 11744
rect 33836 11704 33842 11716
rect 36182 11713 36194 11716
rect 36228 11713 36240 11747
rect 36182 11707 36240 11713
rect 36449 11747 36507 11753
rect 36449 11713 36461 11747
rect 36495 11713 36507 11747
rect 37277 11747 37335 11753
rect 37277 11744 37289 11747
rect 36449 11707 36507 11713
rect 36556 11716 37289 11744
rect 33042 11636 33048 11688
rect 33100 11676 33106 11688
rect 33229 11679 33287 11685
rect 33229 11676 33241 11679
rect 33100 11648 33241 11676
rect 33100 11636 33106 11648
rect 33229 11645 33241 11648
rect 33275 11645 33287 11679
rect 33229 11639 33287 11645
rect 29273 11611 29331 11617
rect 29273 11577 29285 11611
rect 29319 11577 29331 11611
rect 33134 11608 33140 11620
rect 29273 11571 29331 11577
rect 29932 11580 33140 11608
rect 27709 11543 27767 11549
rect 27709 11540 27721 11543
rect 26206 11512 27721 11540
rect 25777 11503 25835 11509
rect 27709 11509 27721 11512
rect 27755 11540 27767 11543
rect 29932 11540 29960 11580
rect 33134 11568 33140 11580
rect 33192 11568 33198 11620
rect 27755 11512 29960 11540
rect 27755 11509 27767 11512
rect 27709 11503 27767 11509
rect 31386 11500 31392 11552
rect 31444 11540 31450 11552
rect 33594 11540 33600 11552
rect 31444 11512 33600 11540
rect 31444 11500 31450 11512
rect 33594 11500 33600 11512
rect 33652 11540 33658 11552
rect 34609 11543 34667 11549
rect 34609 11540 34621 11543
rect 33652 11512 34621 11540
rect 33652 11500 33658 11512
rect 34609 11509 34621 11512
rect 34655 11509 34667 11543
rect 34609 11503 34667 11509
rect 34698 11500 34704 11552
rect 34756 11540 34762 11552
rect 35069 11543 35127 11549
rect 35069 11540 35081 11543
rect 34756 11512 35081 11540
rect 34756 11500 34762 11512
rect 35069 11509 35081 11512
rect 35115 11509 35127 11543
rect 35069 11503 35127 11509
rect 36078 11500 36084 11552
rect 36136 11540 36142 11552
rect 36556 11540 36584 11716
rect 37277 11713 37289 11716
rect 37323 11713 37335 11747
rect 37277 11707 37335 11713
rect 37553 11747 37611 11753
rect 37553 11713 37565 11747
rect 37599 11713 37611 11747
rect 37553 11707 37611 11713
rect 38013 11747 38071 11753
rect 38013 11713 38025 11747
rect 38059 11713 38071 11747
rect 38013 11707 38071 11713
rect 40405 11747 40463 11753
rect 40405 11713 40417 11747
rect 40451 11744 40463 11747
rect 41414 11744 41420 11756
rect 40451 11716 41420 11744
rect 40451 11713 40463 11716
rect 40405 11707 40463 11713
rect 36906 11636 36912 11688
rect 36964 11676 36970 11688
rect 37568 11676 37596 11707
rect 41414 11704 41420 11716
rect 41472 11744 41478 11756
rect 41874 11744 41880 11756
rect 41472 11716 41880 11744
rect 41472 11704 41478 11716
rect 41874 11704 41880 11716
rect 41932 11704 41938 11756
rect 45462 11704 45468 11756
rect 45520 11744 45526 11756
rect 46109 11747 46167 11753
rect 46109 11744 46121 11747
rect 45520 11716 46121 11744
rect 45520 11704 45526 11716
rect 46109 11713 46121 11716
rect 46155 11713 46167 11747
rect 46109 11707 46167 11713
rect 47946 11704 47952 11756
rect 48004 11744 48010 11756
rect 48317 11747 48375 11753
rect 48317 11744 48329 11747
rect 48004 11716 48329 11744
rect 48004 11704 48010 11716
rect 48317 11713 48329 11716
rect 48363 11713 48375 11747
rect 48498 11744 48504 11756
rect 48459 11716 48504 11744
rect 48317 11707 48375 11713
rect 48498 11704 48504 11716
rect 48556 11704 48562 11756
rect 48593 11747 48651 11753
rect 48593 11713 48605 11747
rect 48639 11744 48651 11747
rect 49142 11744 49148 11756
rect 48639 11716 49148 11744
rect 48639 11713 48651 11716
rect 48593 11707 48651 11713
rect 49142 11704 49148 11716
rect 49200 11704 49206 11756
rect 49234 11704 49240 11756
rect 49292 11744 49298 11756
rect 49292 11716 49337 11744
rect 49292 11704 49298 11716
rect 49418 11704 49424 11756
rect 49476 11744 49482 11756
rect 49878 11744 49884 11756
rect 49476 11716 49521 11744
rect 49839 11716 49884 11744
rect 49476 11704 49482 11716
rect 49878 11704 49884 11716
rect 49936 11704 49942 11756
rect 50617 11747 50675 11753
rect 50617 11713 50629 11747
rect 50663 11713 50675 11747
rect 67358 11744 67364 11756
rect 67319 11716 67364 11744
rect 50617 11707 50675 11713
rect 39761 11679 39819 11685
rect 39761 11676 39773 11679
rect 36964 11648 39773 11676
rect 36964 11636 36970 11648
rect 39761 11645 39773 11648
rect 39807 11645 39819 11679
rect 43898 11676 43904 11688
rect 43859 11648 43904 11676
rect 39761 11639 39819 11645
rect 43898 11636 43904 11648
rect 43956 11636 43962 11688
rect 44177 11679 44235 11685
rect 44177 11645 44189 11679
rect 44223 11676 44235 11679
rect 44223 11648 50200 11676
rect 44223 11645 44235 11648
rect 44177 11639 44235 11645
rect 46750 11568 46756 11620
rect 46808 11608 46814 11620
rect 48590 11608 48596 11620
rect 46808 11580 48596 11608
rect 46808 11568 46814 11580
rect 48590 11568 48596 11580
rect 48648 11608 48654 11620
rect 50172 11617 50200 11648
rect 50157 11611 50215 11617
rect 48648 11580 50108 11608
rect 48648 11568 48654 11580
rect 36136 11512 36584 11540
rect 37277 11543 37335 11549
rect 36136 11500 36142 11512
rect 37277 11509 37289 11543
rect 37323 11540 37335 11543
rect 37826 11540 37832 11552
rect 37323 11512 37832 11540
rect 37323 11509 37335 11512
rect 37277 11503 37335 11509
rect 37826 11500 37832 11512
rect 37884 11500 37890 11552
rect 42702 11500 42708 11552
rect 42760 11540 42766 11552
rect 42981 11543 43039 11549
rect 42981 11540 42993 11543
rect 42760 11512 42993 11540
rect 42760 11500 42766 11512
rect 42981 11509 42993 11512
rect 43027 11509 43039 11543
rect 42981 11503 43039 11509
rect 46934 11500 46940 11552
rect 46992 11540 46998 11552
rect 48133 11543 48191 11549
rect 48133 11540 48145 11543
rect 46992 11512 48145 11540
rect 46992 11500 46998 11512
rect 48133 11509 48145 11512
rect 48179 11509 48191 11543
rect 48133 11503 48191 11509
rect 48866 11500 48872 11552
rect 48924 11540 48930 11552
rect 49053 11543 49111 11549
rect 49053 11540 49065 11543
rect 48924 11512 49065 11540
rect 48924 11500 48930 11512
rect 49053 11509 49065 11512
rect 49099 11509 49111 11543
rect 50080 11540 50108 11580
rect 50157 11577 50169 11611
rect 50203 11577 50215 11611
rect 50157 11571 50215 11577
rect 50632 11540 50660 11707
rect 67358 11704 67364 11716
rect 67416 11704 67422 11756
rect 67542 11540 67548 11552
rect 50080 11512 50660 11540
rect 67503 11512 67548 11540
rect 49053 11503 49111 11509
rect 67542 11500 67548 11512
rect 67600 11500 67606 11552
rect 1104 11450 68816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 65654 11450
rect 65706 11398 65718 11450
rect 65770 11398 65782 11450
rect 65834 11398 65846 11450
rect 65898 11398 65910 11450
rect 65962 11398 68816 11450
rect 1104 11376 68816 11398
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 8297 11339 8355 11345
rect 7340 11308 8248 11336
rect 7340 11296 7346 11308
rect 6181 11271 6239 11277
rect 6181 11237 6193 11271
rect 6227 11268 6239 11271
rect 8113 11271 8171 11277
rect 6227 11240 6776 11268
rect 6227 11237 6239 11240
rect 6181 11231 6239 11237
rect 6748 11212 6776 11240
rect 8113 11237 8125 11271
rect 8159 11237 8171 11271
rect 8220 11268 8248 11308
rect 8297 11305 8309 11339
rect 8343 11336 8355 11339
rect 8386 11336 8392 11348
rect 8343 11308 8392 11336
rect 8343 11305 8355 11308
rect 8297 11299 8355 11305
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 11238 11336 11244 11348
rect 11199 11308 11244 11336
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 12250 11336 12256 11348
rect 12211 11308 12256 11336
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 13541 11339 13599 11345
rect 13541 11336 13553 11339
rect 12820 11308 13553 11336
rect 12820 11268 12848 11308
rect 13541 11305 13553 11308
rect 13587 11336 13599 11339
rect 14826 11336 14832 11348
rect 13587 11308 14832 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 14826 11296 14832 11308
rect 14884 11336 14890 11348
rect 19245 11339 19303 11345
rect 14884 11308 18736 11336
rect 14884 11296 14890 11308
rect 8220 11240 12848 11268
rect 8113 11231 8171 11237
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 4801 11203 4859 11209
rect 4801 11200 4813 11203
rect 4764 11172 4813 11200
rect 4764 11160 4770 11172
rect 4801 11169 4813 11172
rect 4847 11169 4859 11203
rect 4801 11163 4859 11169
rect 6730 11160 6736 11212
rect 6788 11200 6794 11212
rect 7837 11203 7895 11209
rect 7837 11200 7849 11203
rect 6788 11172 7849 11200
rect 6788 11160 6794 11172
rect 7837 11169 7849 11172
rect 7883 11200 7895 11203
rect 7926 11200 7932 11212
rect 7883 11172 7932 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 5068 11067 5126 11073
rect 5068 11033 5080 11067
rect 5114 11064 5126 11067
rect 5166 11064 5172 11076
rect 5114 11036 5172 11064
rect 5114 11033 5126 11036
rect 5068 11027 5126 11033
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 8128 11064 8156 11231
rect 8478 11160 8484 11212
rect 8536 11200 8542 11212
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 8536 11172 9045 11200
rect 8536 11160 8542 11172
rect 9033 11169 9045 11172
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11200 12771 11203
rect 12820 11200 12848 11240
rect 13446 11228 13452 11280
rect 13504 11268 13510 11280
rect 14461 11271 14519 11277
rect 14461 11268 14473 11271
rect 13504 11240 14473 11268
rect 13504 11228 13510 11240
rect 14461 11237 14473 11240
rect 14507 11237 14519 11271
rect 14461 11231 14519 11237
rect 16485 11271 16543 11277
rect 16485 11237 16497 11271
rect 16531 11268 16543 11271
rect 16758 11268 16764 11280
rect 16531 11240 16764 11268
rect 16531 11237 16543 11240
rect 16485 11231 16543 11237
rect 16758 11228 16764 11240
rect 16816 11268 16822 11280
rect 18598 11268 18604 11280
rect 16816 11240 18604 11268
rect 16816 11228 16822 11240
rect 18598 11228 18604 11240
rect 18656 11228 18662 11280
rect 18708 11277 18736 11308
rect 19245 11305 19257 11339
rect 19291 11336 19303 11339
rect 19426 11336 19432 11348
rect 19291 11308 19432 11336
rect 19291 11305 19303 11308
rect 19245 11299 19303 11305
rect 19426 11296 19432 11308
rect 19484 11296 19490 11348
rect 19794 11296 19800 11348
rect 19852 11336 19858 11348
rect 20809 11339 20867 11345
rect 20809 11336 20821 11339
rect 19852 11308 20821 11336
rect 19852 11296 19858 11308
rect 20809 11305 20821 11308
rect 20855 11336 20867 11339
rect 21174 11336 21180 11348
rect 20855 11308 21180 11336
rect 20855 11305 20867 11308
rect 20809 11299 20867 11305
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 21637 11339 21695 11345
rect 21637 11305 21649 11339
rect 21683 11305 21695 11339
rect 21637 11299 21695 11305
rect 23109 11339 23167 11345
rect 23109 11305 23121 11339
rect 23155 11336 23167 11339
rect 23290 11336 23296 11348
rect 23155 11308 23296 11336
rect 23155 11305 23167 11308
rect 23109 11299 23167 11305
rect 18693 11271 18751 11277
rect 18693 11237 18705 11271
rect 18739 11268 18751 11271
rect 21082 11268 21088 11280
rect 18739 11240 21088 11268
rect 18739 11237 18751 11240
rect 18693 11231 18751 11237
rect 12759 11172 12848 11200
rect 12897 11203 12955 11209
rect 12759 11169 12771 11172
rect 12713 11163 12771 11169
rect 12897 11169 12909 11203
rect 12943 11200 12955 11203
rect 13078 11200 13084 11212
rect 12943 11172 13084 11200
rect 12943 11169 12955 11172
rect 12897 11163 12955 11169
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 14734 11200 14740 11212
rect 14695 11172 14740 11200
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 16669 11203 16727 11209
rect 16669 11169 16681 11203
rect 16715 11200 16727 11203
rect 16850 11200 16856 11212
rect 16715 11172 16856 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 16850 11160 16856 11172
rect 16908 11200 16914 11212
rect 19720 11209 19748 11240
rect 21082 11228 21088 11240
rect 21140 11228 21146 11280
rect 19705 11203 19763 11209
rect 16908 11172 17632 11200
rect 16908 11160 16914 11172
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 8444 11104 9137 11132
rect 8444 11092 8450 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 12618 11132 12624 11144
rect 12579 11104 12624 11132
rect 9125 11095 9183 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 14829 11135 14887 11141
rect 14829 11101 14841 11135
rect 14875 11132 14887 11135
rect 17497 11135 17555 11141
rect 17497 11132 17509 11135
rect 14875 11104 17509 11132
rect 14875 11101 14887 11104
rect 14829 11095 14887 11101
rect 17497 11101 17509 11104
rect 17543 11101 17555 11135
rect 17497 11095 17555 11101
rect 8570 11064 8576 11076
rect 8128 11036 8576 11064
rect 8570 11024 8576 11036
rect 8628 11064 8634 11076
rect 16209 11067 16267 11073
rect 8628 11036 9628 11064
rect 8628 11024 8634 11036
rect 9600 11008 9628 11036
rect 12636 11036 12848 11064
rect 9490 10996 9496 11008
rect 9451 10968 9496 10996
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 9582 10956 9588 11008
rect 9640 10996 9646 11008
rect 12636 10996 12664 11036
rect 9640 10968 12664 10996
rect 12820 10996 12848 11036
rect 13372 11036 13584 11064
rect 13372 10996 13400 11036
rect 12820 10968 13400 10996
rect 13556 10996 13584 11036
rect 16209 11033 16221 11067
rect 16255 11064 16267 11067
rect 16942 11064 16948 11076
rect 16255 11036 16948 11064
rect 16255 11033 16267 11036
rect 16209 11027 16267 11033
rect 16942 11024 16948 11036
rect 17000 11024 17006 11076
rect 17126 11064 17132 11076
rect 17087 11036 17132 11064
rect 17126 11024 17132 11036
rect 17184 11024 17190 11076
rect 17313 11067 17371 11073
rect 17313 11033 17325 11067
rect 17359 11064 17371 11067
rect 17604 11064 17632 11172
rect 19705 11169 19717 11203
rect 19751 11169 19763 11203
rect 19705 11163 19763 11169
rect 19889 11203 19947 11209
rect 19889 11169 19901 11203
rect 19935 11200 19947 11203
rect 20070 11200 20076 11212
rect 19935 11172 20076 11200
rect 19935 11169 19947 11172
rect 19889 11163 19947 11169
rect 20070 11160 20076 11172
rect 20128 11200 20134 11212
rect 20530 11200 20536 11212
rect 20128 11172 20536 11200
rect 20128 11160 20134 11172
rect 20530 11160 20536 11172
rect 20588 11160 20594 11212
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11132 19671 11135
rect 19978 11132 19984 11144
rect 19659 11104 19984 11132
rect 19659 11101 19671 11104
rect 19613 11095 19671 11101
rect 19978 11092 19984 11104
rect 20036 11132 20042 11144
rect 20901 11135 20959 11141
rect 20901 11132 20913 11135
rect 20036 11104 20913 11132
rect 20036 11092 20042 11104
rect 20901 11101 20913 11104
rect 20947 11132 20959 11135
rect 21652 11132 21680 11299
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 26421 11339 26479 11345
rect 26421 11305 26433 11339
rect 26467 11336 26479 11339
rect 28902 11336 28908 11348
rect 26467 11308 28908 11336
rect 26467 11305 26479 11308
rect 26421 11299 26479 11305
rect 28902 11296 28908 11308
rect 28960 11296 28966 11348
rect 28994 11296 29000 11348
rect 29052 11336 29058 11348
rect 29549 11339 29607 11345
rect 29549 11336 29561 11339
rect 29052 11308 29561 11336
rect 29052 11296 29058 11308
rect 29549 11305 29561 11308
rect 29595 11305 29607 11339
rect 29549 11299 29607 11305
rect 30009 11339 30067 11345
rect 30009 11305 30021 11339
rect 30055 11336 30067 11339
rect 30190 11336 30196 11348
rect 30055 11308 30196 11336
rect 30055 11305 30067 11308
rect 30009 11299 30067 11305
rect 30190 11296 30196 11308
rect 30248 11296 30254 11348
rect 31294 11336 31300 11348
rect 31255 11308 31300 11336
rect 31294 11296 31300 11308
rect 31352 11296 31358 11348
rect 33778 11336 33784 11348
rect 33739 11308 33784 11336
rect 33778 11296 33784 11308
rect 33836 11296 33842 11348
rect 36078 11296 36084 11348
rect 36136 11336 36142 11348
rect 36725 11339 36783 11345
rect 36725 11336 36737 11339
rect 36136 11308 36737 11336
rect 36136 11296 36142 11308
rect 36725 11305 36737 11308
rect 36771 11305 36783 11339
rect 36725 11299 36783 11305
rect 38562 11296 38568 11348
rect 38620 11336 38626 11348
rect 39853 11339 39911 11345
rect 39853 11336 39865 11339
rect 38620 11308 39865 11336
rect 38620 11296 38626 11308
rect 39853 11305 39865 11308
rect 39899 11305 39911 11339
rect 39853 11299 39911 11305
rect 43717 11339 43775 11345
rect 43717 11305 43729 11339
rect 43763 11336 43775 11339
rect 43806 11336 43812 11348
rect 43763 11308 43812 11336
rect 43763 11305 43775 11308
rect 43717 11299 43775 11305
rect 43806 11296 43812 11308
rect 43864 11336 43870 11348
rect 44174 11336 44180 11348
rect 43864 11308 44180 11336
rect 43864 11296 43870 11308
rect 44174 11296 44180 11308
rect 44232 11296 44238 11348
rect 46750 11336 46756 11348
rect 46711 11308 46756 11336
rect 46750 11296 46756 11308
rect 46808 11296 46814 11348
rect 48130 11336 48136 11348
rect 48091 11308 48136 11336
rect 48130 11296 48136 11308
rect 48188 11296 48194 11348
rect 49053 11339 49111 11345
rect 49053 11305 49065 11339
rect 49099 11336 49111 11339
rect 49878 11336 49884 11348
rect 49099 11308 49884 11336
rect 49099 11305 49111 11308
rect 49053 11299 49111 11305
rect 49878 11296 49884 11308
rect 49936 11296 49942 11348
rect 50341 11339 50399 11345
rect 50341 11305 50353 11339
rect 50387 11305 50399 11339
rect 67358 11336 67364 11348
rect 67319 11308 67364 11336
rect 50341 11299 50399 11305
rect 21910 11228 21916 11280
rect 21968 11268 21974 11280
rect 22373 11271 22431 11277
rect 22373 11268 22385 11271
rect 21968 11240 22385 11268
rect 21968 11228 21974 11240
rect 22373 11237 22385 11240
rect 22419 11268 22431 11271
rect 23566 11268 23572 11280
rect 22419 11240 23572 11268
rect 22419 11237 22431 11240
rect 22373 11231 22431 11237
rect 23566 11228 23572 11240
rect 23624 11228 23630 11280
rect 25317 11271 25375 11277
rect 25317 11237 25329 11271
rect 25363 11268 25375 11271
rect 26786 11268 26792 11280
rect 25363 11240 26792 11268
rect 25363 11237 25375 11240
rect 25317 11231 25375 11237
rect 26786 11228 26792 11240
rect 26844 11228 26850 11280
rect 28258 11268 28264 11280
rect 28219 11240 28264 11268
rect 28258 11228 28264 11240
rect 28316 11228 28322 11280
rect 28445 11271 28503 11277
rect 28445 11237 28457 11271
rect 28491 11268 28503 11271
rect 29454 11268 29460 11280
rect 28491 11240 29460 11268
rect 28491 11237 28503 11240
rect 28445 11231 28503 11237
rect 29454 11228 29460 11240
rect 29512 11228 29518 11280
rect 33134 11228 33140 11280
rect 33192 11268 33198 11280
rect 47213 11271 47271 11277
rect 33192 11240 38056 11268
rect 33192 11228 33198 11240
rect 20947 11104 21680 11132
rect 21821 11135 21879 11141
rect 20947 11101 20959 11104
rect 20901 11095 20959 11101
rect 21821 11101 21833 11135
rect 21867 11132 21879 11135
rect 21928 11132 21956 11228
rect 22094 11160 22100 11212
rect 22152 11200 22158 11212
rect 22646 11200 22652 11212
rect 22152 11172 22652 11200
rect 22152 11160 22158 11172
rect 22646 11160 22652 11172
rect 22704 11200 22710 11212
rect 23293 11203 23351 11209
rect 23293 11200 23305 11203
rect 22704 11172 23305 11200
rect 22704 11160 22710 11172
rect 23293 11169 23305 11172
rect 23339 11169 23351 11203
rect 25222 11200 25228 11212
rect 23293 11163 23351 11169
rect 23400 11172 25228 11200
rect 23400 11141 23428 11172
rect 21867 11104 21956 11132
rect 23385 11135 23443 11141
rect 21867 11101 21879 11104
rect 21821 11095 21879 11101
rect 23385 11101 23397 11135
rect 23431 11101 23443 11135
rect 24854 11132 24860 11144
rect 24815 11104 24860 11132
rect 23385 11095 23443 11101
rect 17359 11036 17632 11064
rect 17359 11033 17371 11036
rect 17313 11027 17371 11033
rect 21174 11024 21180 11076
rect 21232 11064 21238 11076
rect 21836 11064 21864 11095
rect 24854 11092 24860 11104
rect 24912 11092 24918 11144
rect 24964 11141 24992 11172
rect 25222 11160 25228 11172
rect 25280 11160 25286 11212
rect 26326 11160 26332 11212
rect 26384 11200 26390 11212
rect 26881 11203 26939 11209
rect 26881 11200 26893 11203
rect 26384 11172 26893 11200
rect 26384 11160 26390 11172
rect 26881 11169 26893 11172
rect 26927 11169 26939 11203
rect 26881 11163 26939 11169
rect 27985 11203 28043 11209
rect 27985 11169 27997 11203
rect 28031 11200 28043 11203
rect 28074 11200 28080 11212
rect 28031 11172 28080 11200
rect 28031 11169 28043 11172
rect 27985 11163 28043 11169
rect 28074 11160 28080 11172
rect 28132 11160 28138 11212
rect 29086 11160 29092 11212
rect 29144 11200 29150 11212
rect 29641 11203 29699 11209
rect 29641 11200 29653 11203
rect 29144 11172 29653 11200
rect 29144 11160 29150 11172
rect 29641 11169 29653 11172
rect 29687 11169 29699 11203
rect 29641 11163 29699 11169
rect 30745 11203 30803 11209
rect 30745 11169 30757 11203
rect 30791 11200 30803 11203
rect 30791 11172 31616 11200
rect 30791 11169 30803 11172
rect 30745 11163 30803 11169
rect 24949 11135 25007 11141
rect 24949 11101 24961 11135
rect 24995 11101 25007 11135
rect 24949 11095 25007 11101
rect 25133 11135 25191 11141
rect 25133 11101 25145 11135
rect 25179 11132 25191 11135
rect 26053 11135 26111 11141
rect 26053 11132 26065 11135
rect 25179 11104 26065 11132
rect 25179 11101 25191 11104
rect 25133 11095 25191 11101
rect 26053 11101 26065 11104
rect 26099 11101 26111 11135
rect 26053 11095 26111 11101
rect 21232 11036 21864 11064
rect 21232 11024 21238 11036
rect 24486 11024 24492 11076
rect 24544 11064 24550 11076
rect 25148 11064 25176 11095
rect 26234 11092 26240 11144
rect 26292 11132 26298 11144
rect 29825 11135 29883 11141
rect 26292 11104 26337 11132
rect 26292 11092 26298 11104
rect 29825 11101 29837 11135
rect 29871 11132 29883 11135
rect 30466 11132 30472 11144
rect 29871 11104 30472 11132
rect 29871 11101 29883 11104
rect 29825 11095 29883 11101
rect 30466 11092 30472 11104
rect 30524 11092 30530 11144
rect 30929 11135 30987 11141
rect 30929 11101 30941 11135
rect 30975 11132 30987 11135
rect 31202 11132 31208 11144
rect 30975 11104 31208 11132
rect 30975 11101 30987 11104
rect 30929 11095 30987 11101
rect 31202 11092 31208 11104
rect 31260 11092 31266 11144
rect 24544 11036 25176 11064
rect 24544 11024 24550 11036
rect 29178 11024 29184 11076
rect 29236 11064 29242 11076
rect 29549 11067 29607 11073
rect 29549 11064 29561 11067
rect 29236 11036 29561 11064
rect 29236 11024 29242 11036
rect 29549 11033 29561 11036
rect 29595 11033 29607 11067
rect 29549 11027 29607 11033
rect 30742 11024 30748 11076
rect 30800 11064 30806 11076
rect 30837 11067 30895 11073
rect 30837 11064 30849 11067
rect 30800 11036 30849 11064
rect 30800 11024 30806 11036
rect 30837 11033 30849 11036
rect 30883 11064 30895 11067
rect 31588 11064 31616 11172
rect 36906 11160 36912 11212
rect 36964 11200 36970 11212
rect 36964 11172 37504 11200
rect 36964 11160 36970 11172
rect 31662 11092 31668 11144
rect 31720 11132 31726 11144
rect 32870 11135 32928 11141
rect 32870 11132 32882 11135
rect 31720 11104 32882 11132
rect 31720 11092 31726 11104
rect 32870 11101 32882 11104
rect 32916 11101 32928 11135
rect 32870 11095 32928 11101
rect 33042 11092 33048 11144
rect 33100 11132 33106 11144
rect 33137 11135 33195 11141
rect 33137 11132 33149 11135
rect 33100 11104 33149 11132
rect 33100 11092 33106 11104
rect 33137 11101 33149 11104
rect 33183 11101 33195 11135
rect 33594 11132 33600 11144
rect 33555 11104 33600 11132
rect 33137 11095 33195 11101
rect 33594 11092 33600 11104
rect 33652 11092 33658 11144
rect 37274 11132 37280 11144
rect 37235 11104 37280 11132
rect 37274 11092 37280 11104
rect 37332 11092 37338 11144
rect 37476 11141 37504 11172
rect 37461 11135 37519 11141
rect 37461 11101 37473 11135
rect 37507 11101 37519 11135
rect 38028 11132 38056 11240
rect 47213 11237 47225 11271
rect 47259 11237 47271 11271
rect 47213 11231 47271 11237
rect 38194 11200 38200 11212
rect 38155 11172 38200 11200
rect 38194 11160 38200 11172
rect 38252 11160 38258 11212
rect 38930 11160 38936 11212
rect 38988 11200 38994 11212
rect 41325 11203 41383 11209
rect 41325 11200 41337 11203
rect 38988 11172 41337 11200
rect 38988 11160 38994 11172
rect 41325 11169 41337 11172
rect 41371 11169 41383 11203
rect 41598 11200 41604 11212
rect 41511 11172 41604 11200
rect 41325 11163 41383 11169
rect 41598 11160 41604 11172
rect 41656 11200 41662 11212
rect 43898 11200 43904 11212
rect 41656 11172 43904 11200
rect 41656 11160 41662 11172
rect 43898 11160 43904 11172
rect 43956 11200 43962 11212
rect 45005 11203 45063 11209
rect 45005 11200 45017 11203
rect 43956 11172 45017 11200
rect 43956 11160 43962 11172
rect 45005 11169 45017 11172
rect 45051 11169 45063 11203
rect 45005 11163 45063 11169
rect 45281 11203 45339 11209
rect 45281 11169 45293 11203
rect 45327 11200 45339 11203
rect 47228 11200 47256 11231
rect 48038 11228 48044 11280
rect 48096 11228 48102 11280
rect 48958 11228 48964 11280
rect 49016 11268 49022 11280
rect 50356 11268 50384 11299
rect 67358 11296 67364 11308
rect 67416 11296 67422 11348
rect 50614 11268 50620 11280
rect 49016 11240 50620 11268
rect 49016 11228 49022 11240
rect 50614 11228 50620 11240
rect 50672 11228 50678 11280
rect 51046 11240 55214 11268
rect 45327 11172 47256 11200
rect 48056 11200 48084 11228
rect 48056 11172 48268 11200
rect 45327 11169 45339 11172
rect 45281 11163 45339 11169
rect 38378 11132 38384 11144
rect 38028 11104 38384 11132
rect 37461 11095 37519 11101
rect 38378 11092 38384 11104
rect 38436 11092 38442 11144
rect 38473 11135 38531 11141
rect 38473 11101 38485 11135
rect 38519 11101 38531 11135
rect 38473 11095 38531 11101
rect 39301 11135 39359 11141
rect 39301 11101 39313 11135
rect 39347 11132 39359 11135
rect 39850 11132 39856 11144
rect 39347 11104 39856 11132
rect 39347 11101 39359 11104
rect 39301 11095 39359 11101
rect 33686 11064 33692 11076
rect 30883 11036 31064 11064
rect 31588 11036 33692 11064
rect 30883 11033 30895 11036
rect 30837 11027 30895 11033
rect 16758 10996 16764 11008
rect 13556 10968 16764 10996
rect 9640 10956 9646 10968
rect 16758 10956 16764 10968
rect 16816 10956 16822 11008
rect 19978 10956 19984 11008
rect 20036 10996 20042 11008
rect 20441 10999 20499 11005
rect 20441 10996 20453 10999
rect 20036 10968 20453 10996
rect 20036 10956 20042 10968
rect 20441 10965 20453 10968
rect 20487 10965 20499 10999
rect 21358 10996 21364 11008
rect 21319 10968 21364 10996
rect 20441 10959 20499 10965
rect 21358 10956 21364 10968
rect 21416 10956 21422 11008
rect 31036 10996 31064 11036
rect 33686 11024 33692 11036
rect 33744 11024 33750 11076
rect 36170 11064 36176 11076
rect 36131 11036 36176 11064
rect 36170 11024 36176 11036
rect 36228 11064 36234 11076
rect 37369 11067 37427 11073
rect 37369 11064 37381 11067
rect 36228 11036 37381 11064
rect 36228 11024 36234 11036
rect 37369 11033 37381 11036
rect 37415 11064 37427 11067
rect 38488 11064 38516 11095
rect 39850 11092 39856 11104
rect 39908 11092 39914 11144
rect 42150 11132 42156 11144
rect 42111 11104 42156 11132
rect 42150 11092 42156 11104
rect 42208 11092 42214 11144
rect 42337 11135 42395 11141
rect 42337 11101 42349 11135
rect 42383 11132 42395 11135
rect 42702 11132 42708 11144
rect 42383 11104 42708 11132
rect 42383 11101 42395 11104
rect 42337 11095 42395 11101
rect 42702 11092 42708 11104
rect 42760 11132 42766 11144
rect 42889 11135 42947 11141
rect 42889 11132 42901 11135
rect 42760 11104 42901 11132
rect 42760 11092 42766 11104
rect 42889 11101 42901 11104
rect 42935 11101 42947 11135
rect 42889 11095 42947 11101
rect 43073 11135 43131 11141
rect 43073 11101 43085 11135
rect 43119 11132 43131 11135
rect 43533 11135 43591 11141
rect 43533 11132 43545 11135
rect 43119 11104 43545 11132
rect 43119 11101 43131 11104
rect 43073 11095 43131 11101
rect 43533 11101 43545 11104
rect 43579 11132 43591 11135
rect 44266 11132 44272 11144
rect 43579 11104 44272 11132
rect 43579 11101 43591 11104
rect 43533 11095 43591 11101
rect 44266 11092 44272 11104
rect 44324 11092 44330 11144
rect 47394 11132 47400 11144
rect 47355 11104 47400 11132
rect 47394 11092 47400 11104
rect 47452 11092 47458 11144
rect 48240 11141 48268 11172
rect 48314 11160 48320 11212
rect 48372 11200 48378 11212
rect 51046 11200 51074 11240
rect 48372 11172 51074 11200
rect 48372 11160 48378 11172
rect 48041 11135 48099 11141
rect 48041 11101 48053 11135
rect 48087 11101 48099 11135
rect 48041 11095 48099 11101
rect 48225 11135 48283 11141
rect 48225 11101 48237 11135
rect 48271 11101 48283 11135
rect 48225 11095 48283 11101
rect 37415 11036 38516 11064
rect 37415 11033 37427 11036
rect 37369 11027 37427 11033
rect 40770 11024 40776 11076
rect 40828 11024 40834 11076
rect 44361 11067 44419 11073
rect 44361 11033 44373 11067
rect 44407 11064 44419 11067
rect 44407 11036 45232 11064
rect 44407 11033 44419 11036
rect 44361 11027 44419 11033
rect 31757 10999 31815 11005
rect 31757 10996 31769 10999
rect 31036 10968 31769 10996
rect 31757 10965 31769 10968
rect 31803 10965 31815 10999
rect 45204 10996 45232 11036
rect 45388 11036 45770 11064
rect 45388 10996 45416 11036
rect 47026 11024 47032 11076
rect 47084 11064 47090 11076
rect 48056 11064 48084 11095
rect 48498 11092 48504 11144
rect 48556 11132 48562 11144
rect 48685 11135 48743 11141
rect 48685 11132 48697 11135
rect 48556 11104 48697 11132
rect 48556 11092 48562 11104
rect 48685 11101 48697 11104
rect 48731 11101 48743 11135
rect 48685 11095 48743 11101
rect 48869 11135 48927 11141
rect 48869 11101 48881 11135
rect 48915 11132 48927 11135
rect 48958 11132 48964 11144
rect 48915 11104 48964 11132
rect 48915 11101 48927 11104
rect 48869 11095 48927 11101
rect 48958 11092 48964 11104
rect 49016 11092 49022 11144
rect 49142 11092 49148 11144
rect 49200 11132 49206 11144
rect 49970 11132 49976 11144
rect 49200 11104 49976 11132
rect 49200 11092 49206 11104
rect 49970 11092 49976 11104
rect 50028 11132 50034 11144
rect 55186 11132 55214 11240
rect 67177 11135 67235 11141
rect 67177 11132 67189 11135
rect 50028 11104 50568 11132
rect 55186 11104 67189 11132
rect 50028 11092 50034 11104
rect 48516 11064 48544 11092
rect 50154 11064 50160 11076
rect 47084 11036 48544 11064
rect 50115 11036 50160 11064
rect 47084 11024 47090 11036
rect 50154 11024 50160 11036
rect 50212 11024 50218 11076
rect 45204 10968 45416 10996
rect 31757 10959 31815 10965
rect 49418 10956 49424 11008
rect 49476 10996 49482 11008
rect 50540 11005 50568 11104
rect 67177 11101 67189 11104
rect 67223 11132 67235 11135
rect 67821 11135 67879 11141
rect 67821 11132 67833 11135
rect 67223 11104 67833 11132
rect 67223 11101 67235 11104
rect 67177 11095 67235 11101
rect 67821 11101 67833 11104
rect 67867 11101 67879 11135
rect 67821 11095 67879 11101
rect 50357 10999 50415 11005
rect 50357 10996 50369 10999
rect 49476 10968 50369 10996
rect 49476 10956 49482 10968
rect 50357 10965 50369 10968
rect 50403 10965 50415 10999
rect 50357 10959 50415 10965
rect 50525 10999 50583 11005
rect 50525 10965 50537 10999
rect 50571 10965 50583 10999
rect 50525 10959 50583 10965
rect 1104 10906 68816 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 68816 10906
rect 1104 10832 68816 10854
rect 5166 10792 5172 10804
rect 5127 10764 5172 10792
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 6365 10795 6423 10801
rect 6365 10761 6377 10795
rect 6411 10761 6423 10795
rect 6730 10792 6736 10804
rect 6691 10764 6736 10792
rect 6365 10755 6423 10761
rect 5353 10659 5411 10665
rect 5353 10625 5365 10659
rect 5399 10656 5411 10659
rect 6380 10656 6408 10755
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 8941 10795 8999 10801
rect 8941 10761 8953 10795
rect 8987 10792 8999 10795
rect 9582 10792 9588 10804
rect 8987 10764 9588 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 13265 10795 13323 10801
rect 13265 10761 13277 10795
rect 13311 10761 13323 10795
rect 13722 10792 13728 10804
rect 13683 10764 13728 10792
rect 13265 10755 13323 10761
rect 8294 10684 8300 10736
rect 8352 10724 8358 10736
rect 8389 10727 8447 10733
rect 8389 10724 8401 10727
rect 8352 10696 8401 10724
rect 8352 10684 8358 10696
rect 8389 10693 8401 10696
rect 8435 10693 8447 10727
rect 8389 10687 8447 10693
rect 12894 10684 12900 10736
rect 12952 10724 12958 10736
rect 13280 10724 13308 10755
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 16758 10792 16764 10804
rect 16719 10764 16764 10792
rect 16758 10752 16764 10764
rect 16816 10752 16822 10804
rect 20346 10792 20352 10804
rect 20307 10764 20352 10792
rect 20346 10752 20352 10764
rect 20404 10752 20410 10804
rect 21910 10792 21916 10804
rect 21871 10764 21916 10792
rect 21910 10752 21916 10764
rect 21968 10752 21974 10804
rect 22002 10752 22008 10804
rect 22060 10792 22066 10804
rect 22922 10792 22928 10804
rect 22060 10764 22928 10792
rect 22060 10752 22066 10764
rect 22922 10752 22928 10764
rect 22980 10752 22986 10804
rect 30561 10795 30619 10801
rect 30561 10761 30573 10795
rect 30607 10792 30619 10795
rect 30650 10792 30656 10804
rect 30607 10764 30656 10792
rect 30607 10761 30619 10764
rect 30561 10755 30619 10761
rect 30650 10752 30656 10764
rect 30708 10752 30714 10804
rect 31938 10752 31944 10804
rect 31996 10792 32002 10804
rect 32493 10795 32551 10801
rect 32493 10792 32505 10795
rect 31996 10764 32505 10792
rect 31996 10752 32002 10764
rect 32493 10761 32505 10764
rect 32539 10761 32551 10795
rect 33502 10792 33508 10804
rect 33463 10764 33508 10792
rect 32493 10755 32551 10761
rect 33502 10752 33508 10764
rect 33560 10752 33566 10804
rect 33594 10752 33600 10804
rect 33652 10792 33658 10804
rect 33873 10795 33931 10801
rect 33873 10792 33885 10795
rect 33652 10764 33885 10792
rect 33652 10752 33658 10764
rect 33873 10761 33885 10764
rect 33919 10761 33931 10795
rect 33873 10755 33931 10761
rect 38565 10795 38623 10801
rect 38565 10761 38577 10795
rect 38611 10792 38623 10795
rect 38930 10792 38936 10804
rect 38611 10764 38936 10792
rect 38611 10761 38623 10764
rect 38565 10755 38623 10761
rect 38930 10752 38936 10764
rect 38988 10752 38994 10804
rect 40770 10792 40776 10804
rect 40731 10764 40776 10792
rect 40770 10752 40776 10764
rect 40828 10752 40834 10804
rect 42702 10752 42708 10804
rect 42760 10792 42766 10804
rect 43165 10795 43223 10801
rect 43165 10792 43177 10795
rect 42760 10764 43177 10792
rect 42760 10752 42766 10764
rect 43165 10761 43177 10764
rect 43211 10761 43223 10795
rect 46934 10792 46940 10804
rect 43165 10755 43223 10761
rect 44100 10764 46940 10792
rect 12952 10696 14136 10724
rect 12952 10684 12958 10696
rect 5399 10628 6408 10656
rect 5399 10625 5411 10628
rect 5353 10619 5411 10625
rect 6454 10616 6460 10668
rect 6512 10656 6518 10668
rect 8110 10656 8116 10668
rect 6512 10628 6960 10656
rect 8071 10628 8116 10656
rect 6512 10616 6518 10628
rect 6932 10597 6960 10628
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 8202 10616 8208 10668
rect 8260 10656 8266 10668
rect 12158 10665 12164 10668
rect 8260 10628 8305 10656
rect 8260 10616 8266 10628
rect 12152 10619 12164 10665
rect 12216 10656 12222 10668
rect 14108 10665 14136 10696
rect 23474 10684 23480 10736
rect 23532 10724 23538 10736
rect 30834 10724 30840 10736
rect 23532 10696 30840 10724
rect 23532 10684 23538 10696
rect 30834 10684 30840 10696
rect 30892 10684 30898 10736
rect 33413 10727 33471 10733
rect 33413 10724 33425 10727
rect 31404 10696 33425 10724
rect 14093 10659 14151 10665
rect 12216 10628 12252 10656
rect 12158 10616 12164 10619
rect 12216 10616 12222 10628
rect 14093 10625 14105 10659
rect 14139 10625 14151 10659
rect 14093 10619 14151 10625
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10656 15623 10659
rect 15654 10656 15660 10668
rect 15611 10628 15660 10656
rect 15611 10625 15623 10628
rect 15565 10619 15623 10625
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 20806 10656 20812 10668
rect 20767 10628 20812 10656
rect 20806 10616 20812 10628
rect 20864 10616 20870 10668
rect 25869 10659 25927 10665
rect 25869 10625 25881 10659
rect 25915 10656 25927 10659
rect 26418 10656 26424 10668
rect 25915 10628 26424 10656
rect 25915 10625 25927 10628
rect 25869 10619 25927 10625
rect 26418 10616 26424 10628
rect 26476 10656 26482 10668
rect 26970 10656 26976 10668
rect 26476 10628 26976 10656
rect 26476 10616 26482 10628
rect 26970 10616 26976 10628
rect 27028 10616 27034 10668
rect 29273 10659 29331 10665
rect 29273 10625 29285 10659
rect 29319 10656 29331 10659
rect 30742 10656 30748 10668
rect 29319 10628 30748 10656
rect 29319 10625 29331 10628
rect 29273 10619 29331 10625
rect 30742 10616 30748 10628
rect 30800 10616 30806 10668
rect 30929 10659 30987 10665
rect 30929 10625 30941 10659
rect 30975 10656 30987 10659
rect 31404 10656 31432 10696
rect 33413 10693 33425 10696
rect 33459 10724 33471 10727
rect 34698 10724 34704 10736
rect 33459 10696 34704 10724
rect 33459 10693 33471 10696
rect 33413 10687 33471 10693
rect 34698 10684 34704 10696
rect 34756 10684 34762 10736
rect 38194 10724 38200 10736
rect 37568 10696 38200 10724
rect 30975 10628 31432 10656
rect 30975 10625 30987 10628
rect 30929 10619 30987 10625
rect 31478 10616 31484 10668
rect 31536 10656 31542 10668
rect 32125 10659 32183 10665
rect 32125 10656 32137 10659
rect 31536 10628 32137 10656
rect 31536 10616 31542 10628
rect 32125 10625 32137 10628
rect 32171 10625 32183 10659
rect 32306 10656 32312 10668
rect 32267 10628 32312 10656
rect 32125 10619 32183 10625
rect 32306 10616 32312 10628
rect 32364 10616 32370 10668
rect 32582 10616 32588 10668
rect 32640 10656 32646 10668
rect 37568 10665 37596 10696
rect 38194 10684 38200 10696
rect 38252 10684 38258 10736
rect 38378 10684 38384 10736
rect 38436 10724 38442 10736
rect 39117 10727 39175 10733
rect 39117 10724 39129 10727
rect 38436 10696 39129 10724
rect 38436 10684 38442 10696
rect 39117 10693 39129 10696
rect 39163 10693 39175 10727
rect 41325 10727 41383 10733
rect 41325 10724 41337 10727
rect 39117 10687 39175 10693
rect 40512 10696 41337 10724
rect 37553 10659 37611 10665
rect 32640 10628 32685 10656
rect 32640 10616 32646 10628
rect 37553 10625 37565 10659
rect 37599 10625 37611 10659
rect 37826 10656 37832 10668
rect 37787 10628 37832 10656
rect 37553 10619 37611 10625
rect 37826 10616 37832 10628
rect 37884 10616 37890 10668
rect 39132 10656 39160 10687
rect 40512 10668 40540 10696
rect 41325 10693 41337 10696
rect 41371 10724 41383 10727
rect 41371 10696 42472 10724
rect 41371 10693 41383 10696
rect 41325 10687 41383 10693
rect 40221 10659 40279 10665
rect 40221 10656 40233 10659
rect 39132 10628 40233 10656
rect 40221 10625 40233 10628
rect 40267 10656 40279 10659
rect 40494 10656 40500 10668
rect 40267 10628 40500 10656
rect 40267 10625 40279 10628
rect 40221 10619 40279 10625
rect 40494 10616 40500 10628
rect 40552 10616 40558 10668
rect 40865 10659 40923 10665
rect 40865 10625 40877 10659
rect 40911 10656 40923 10659
rect 41414 10656 41420 10668
rect 40911 10628 41420 10656
rect 40911 10625 40923 10628
rect 40865 10619 40923 10625
rect 41414 10616 41420 10628
rect 41472 10616 41478 10668
rect 42444 10665 42472 10696
rect 42429 10659 42487 10665
rect 42429 10625 42441 10659
rect 42475 10656 42487 10659
rect 42720 10656 42748 10752
rect 44100 10733 44128 10764
rect 46934 10752 46940 10764
rect 46992 10752 46998 10804
rect 47026 10752 47032 10804
rect 47084 10792 47090 10804
rect 47084 10764 47129 10792
rect 47084 10752 47090 10764
rect 47394 10752 47400 10804
rect 47452 10792 47458 10804
rect 47581 10795 47639 10801
rect 47581 10792 47593 10795
rect 47452 10764 47593 10792
rect 47452 10752 47458 10764
rect 47581 10761 47593 10764
rect 47627 10761 47639 10795
rect 47581 10755 47639 10761
rect 49418 10752 49424 10804
rect 49476 10792 49482 10804
rect 49476 10764 50844 10792
rect 49476 10752 49482 10764
rect 44085 10727 44143 10733
rect 44085 10693 44097 10727
rect 44131 10693 44143 10727
rect 44085 10687 44143 10693
rect 45094 10684 45100 10736
rect 45152 10684 45158 10736
rect 47765 10727 47823 10733
rect 47765 10693 47777 10727
rect 47811 10724 47823 10727
rect 48777 10727 48835 10733
rect 47811 10696 48636 10724
rect 47811 10693 47823 10696
rect 47765 10687 47823 10693
rect 48608 10668 48636 10696
rect 48777 10693 48789 10727
rect 48823 10724 48835 10727
rect 50062 10724 50068 10736
rect 48823 10696 50068 10724
rect 48823 10693 48835 10696
rect 48777 10687 48835 10693
rect 50062 10684 50068 10696
rect 50120 10684 50126 10736
rect 50816 10668 50844 10764
rect 46842 10656 46848 10668
rect 42475 10628 42748 10656
rect 46803 10628 46848 10656
rect 42475 10625 42487 10628
rect 42429 10619 42487 10625
rect 46842 10616 46848 10628
rect 46900 10616 46906 10668
rect 47029 10659 47087 10665
rect 47029 10625 47041 10659
rect 47075 10625 47087 10659
rect 47029 10619 47087 10625
rect 47949 10659 48007 10665
rect 47949 10625 47961 10659
rect 47995 10625 48007 10659
rect 48590 10656 48596 10668
rect 48551 10628 48596 10656
rect 47949 10619 48007 10625
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10557 6975 10591
rect 6917 10551 6975 10557
rect 6840 10464 6868 10551
rect 11514 10548 11520 10600
rect 11572 10588 11578 10600
rect 11885 10591 11943 10597
rect 11885 10588 11897 10591
rect 11572 10560 11897 10588
rect 11572 10548 11578 10560
rect 11885 10557 11897 10560
rect 11931 10557 11943 10591
rect 11885 10551 11943 10557
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10588 14243 10591
rect 15197 10591 15255 10597
rect 15197 10588 15209 10591
rect 14231 10560 15209 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 15197 10557 15209 10560
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 15473 10591 15531 10597
rect 15473 10557 15485 10591
rect 15519 10588 15531 10591
rect 16574 10588 16580 10600
rect 15519 10560 16580 10588
rect 15519 10557 15531 10560
rect 15473 10551 15531 10557
rect 16574 10548 16580 10560
rect 16632 10548 16638 10600
rect 20530 10588 20536 10600
rect 20491 10560 20536 10588
rect 20530 10548 20536 10560
rect 20588 10548 20594 10600
rect 20625 10591 20683 10597
rect 20625 10557 20637 10591
rect 20671 10557 20683 10591
rect 20625 10551 20683 10557
rect 20717 10591 20775 10597
rect 20717 10557 20729 10591
rect 20763 10588 20775 10591
rect 21358 10588 21364 10600
rect 20763 10560 21364 10588
rect 20763 10557 20775 10560
rect 20717 10551 20775 10557
rect 8386 10520 8392 10532
rect 8347 10492 8392 10520
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 20254 10520 20260 10532
rect 13188 10492 20260 10520
rect 6822 10452 6828 10464
rect 6735 10424 6828 10452
rect 6822 10412 6828 10424
rect 6880 10452 6886 10464
rect 7650 10452 7656 10464
rect 6880 10424 7656 10452
rect 6880 10412 6886 10424
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 13188 10452 13216 10492
rect 20254 10480 20260 10492
rect 20312 10480 20318 10532
rect 20640 10464 20668 10551
rect 21358 10548 21364 10560
rect 21416 10548 21422 10600
rect 25958 10588 25964 10600
rect 25871 10560 25964 10588
rect 25958 10548 25964 10560
rect 26016 10588 26022 10600
rect 26142 10588 26148 10600
rect 26016 10560 26148 10588
rect 26016 10548 26022 10560
rect 26142 10548 26148 10560
rect 26200 10548 26206 10600
rect 29178 10588 29184 10600
rect 29139 10560 29184 10588
rect 29178 10548 29184 10560
rect 29236 10548 29242 10600
rect 30837 10591 30895 10597
rect 30837 10557 30849 10591
rect 30883 10557 30895 10591
rect 30837 10551 30895 10557
rect 33321 10591 33379 10597
rect 33321 10557 33333 10591
rect 33367 10588 33379 10591
rect 33686 10588 33692 10600
rect 33367 10560 33692 10588
rect 33367 10557 33379 10560
rect 33321 10551 33379 10557
rect 20990 10480 20996 10532
rect 21048 10520 21054 10532
rect 26237 10523 26295 10529
rect 21048 10492 25176 10520
rect 21048 10480 21054 10492
rect 11848 10424 13216 10452
rect 11848 10412 11854 10424
rect 20622 10412 20628 10464
rect 20680 10412 20686 10464
rect 25038 10452 25044 10464
rect 24999 10424 25044 10452
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 25148 10452 25176 10492
rect 26237 10489 26249 10523
rect 26283 10520 26295 10523
rect 30852 10520 30880 10551
rect 33686 10548 33692 10560
rect 33744 10548 33750 10600
rect 43622 10548 43628 10600
rect 43680 10588 43686 10600
rect 43809 10591 43867 10597
rect 43809 10588 43821 10591
rect 43680 10560 43821 10588
rect 43680 10548 43686 10560
rect 43809 10557 43821 10560
rect 43855 10557 43867 10591
rect 43809 10551 43867 10557
rect 46750 10548 46756 10600
rect 46808 10588 46814 10600
rect 47044 10588 47072 10619
rect 46808 10560 47072 10588
rect 47964 10588 47992 10619
rect 48590 10616 48596 10628
rect 48648 10616 48654 10668
rect 48869 10659 48927 10665
rect 48869 10625 48881 10659
rect 48915 10656 48927 10659
rect 50154 10656 50160 10668
rect 48915 10628 50016 10656
rect 50115 10628 50160 10656
rect 48915 10625 48927 10628
rect 48869 10619 48927 10625
rect 49786 10588 49792 10600
rect 47964 10560 49792 10588
rect 46808 10548 46814 10560
rect 49786 10548 49792 10560
rect 49844 10548 49850 10600
rect 49881 10591 49939 10597
rect 49881 10557 49893 10591
rect 49927 10557 49939 10591
rect 49988 10588 50016 10628
rect 50154 10616 50160 10628
rect 50212 10616 50218 10668
rect 50614 10656 50620 10668
rect 50575 10628 50620 10656
rect 50614 10616 50620 10628
rect 50672 10616 50678 10668
rect 50798 10616 50804 10668
rect 50856 10656 50862 10668
rect 50856 10628 50949 10656
rect 50856 10616 50862 10628
rect 50706 10588 50712 10600
rect 49988 10560 50712 10588
rect 49881 10551 49939 10557
rect 26283 10492 30880 10520
rect 40037 10523 40095 10529
rect 26283 10489 26295 10492
rect 26237 10483 26295 10489
rect 40037 10489 40049 10523
rect 40083 10520 40095 10523
rect 40586 10520 40592 10532
rect 40083 10492 40592 10520
rect 40083 10489 40095 10492
rect 40037 10483 40095 10489
rect 40586 10480 40592 10492
rect 40644 10520 40650 10532
rect 43530 10520 43536 10532
rect 40644 10492 43536 10520
rect 40644 10480 40650 10492
rect 43530 10480 43536 10492
rect 43588 10480 43594 10532
rect 45557 10523 45615 10529
rect 45557 10489 45569 10523
rect 45603 10520 45615 10523
rect 49418 10520 49424 10532
rect 45603 10492 49424 10520
rect 45603 10489 45615 10492
rect 45557 10483 45615 10489
rect 49418 10480 49424 10492
rect 49476 10480 49482 10532
rect 49602 10480 49608 10532
rect 49660 10520 49666 10532
rect 49896 10520 49924 10551
rect 50706 10548 50712 10560
rect 50764 10548 50770 10600
rect 49660 10492 49924 10520
rect 49660 10480 49666 10492
rect 29546 10452 29552 10464
rect 25148 10424 29552 10452
rect 29546 10412 29552 10424
rect 29604 10412 29610 10464
rect 29641 10455 29699 10461
rect 29641 10421 29653 10455
rect 29687 10452 29699 10455
rect 30374 10452 30380 10464
rect 29687 10424 30380 10452
rect 29687 10421 29699 10424
rect 29641 10415 29699 10421
rect 30374 10412 30380 10424
rect 30432 10412 30438 10464
rect 30834 10412 30840 10464
rect 30892 10452 30898 10464
rect 31846 10452 31852 10464
rect 30892 10424 31852 10452
rect 30892 10412 30898 10424
rect 31846 10412 31852 10424
rect 31904 10452 31910 10464
rect 39022 10452 39028 10464
rect 31904 10424 39028 10452
rect 31904 10412 31910 10424
rect 39022 10412 39028 10424
rect 39080 10452 39086 10464
rect 39209 10455 39267 10461
rect 39209 10452 39221 10455
rect 39080 10424 39221 10452
rect 39080 10412 39086 10424
rect 39209 10421 39221 10424
rect 39255 10421 39267 10455
rect 42610 10452 42616 10464
rect 42571 10424 42616 10452
rect 39209 10415 39267 10421
rect 42610 10412 42616 10424
rect 42668 10412 42674 10464
rect 48406 10452 48412 10464
rect 48367 10424 48412 10452
rect 48406 10412 48412 10424
rect 48464 10412 48470 10464
rect 50801 10455 50859 10461
rect 50801 10421 50813 10455
rect 50847 10452 50859 10455
rect 50890 10452 50896 10464
rect 50847 10424 50896 10452
rect 50847 10421 50859 10424
rect 50801 10415 50859 10421
rect 50890 10412 50896 10424
rect 50948 10412 50954 10464
rect 1104 10362 68816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 65654 10362
rect 65706 10310 65718 10362
rect 65770 10310 65782 10362
rect 65834 10310 65846 10362
rect 65898 10310 65910 10362
rect 65962 10310 68816 10362
rect 1104 10288 68816 10310
rect 7650 10208 7656 10260
rect 7708 10248 7714 10260
rect 12069 10251 12127 10257
rect 7708 10220 9352 10248
rect 7708 10208 7714 10220
rect 9122 10140 9128 10192
rect 9180 10180 9186 10192
rect 9217 10183 9275 10189
rect 9217 10180 9229 10183
rect 9180 10152 9229 10180
rect 9180 10140 9186 10152
rect 9217 10149 9229 10152
rect 9263 10149 9275 10183
rect 9324 10180 9352 10220
rect 12069 10217 12081 10251
rect 12115 10248 12127 10251
rect 12158 10248 12164 10260
rect 12115 10220 12164 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 12158 10208 12164 10220
rect 12216 10208 12222 10260
rect 16209 10251 16267 10257
rect 16209 10217 16221 10251
rect 16255 10248 16267 10251
rect 17126 10248 17132 10260
rect 16255 10220 17132 10248
rect 16255 10217 16267 10220
rect 16209 10211 16267 10217
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 20530 10208 20536 10260
rect 20588 10248 20594 10260
rect 20809 10251 20867 10257
rect 20809 10248 20821 10251
rect 20588 10220 20821 10248
rect 20588 10208 20594 10220
rect 20809 10217 20821 10220
rect 20855 10217 20867 10251
rect 20809 10211 20867 10217
rect 21177 10251 21235 10257
rect 21177 10217 21189 10251
rect 21223 10248 21235 10251
rect 21542 10248 21548 10260
rect 21223 10220 21548 10248
rect 21223 10217 21235 10220
rect 21177 10211 21235 10217
rect 21542 10208 21548 10220
rect 21600 10208 21606 10260
rect 25958 10248 25964 10260
rect 25919 10220 25964 10248
rect 25958 10208 25964 10220
rect 26016 10208 26022 10260
rect 26145 10251 26203 10257
rect 26145 10217 26157 10251
rect 26191 10248 26203 10251
rect 26234 10248 26240 10260
rect 26191 10220 26240 10248
rect 26191 10217 26203 10220
rect 26145 10211 26203 10217
rect 26234 10208 26240 10220
rect 26292 10208 26298 10260
rect 28353 10251 28411 10257
rect 28353 10217 28365 10251
rect 28399 10248 28411 10251
rect 29178 10248 29184 10260
rect 28399 10220 29184 10248
rect 28399 10217 28411 10220
rect 28353 10211 28411 10217
rect 29178 10208 29184 10220
rect 29236 10208 29242 10260
rect 30377 10251 30435 10257
rect 30377 10217 30389 10251
rect 30423 10248 30435 10251
rect 30926 10248 30932 10260
rect 30423 10220 30932 10248
rect 30423 10217 30435 10220
rect 30377 10211 30435 10217
rect 30926 10208 30932 10220
rect 30984 10208 30990 10260
rect 31202 10248 31208 10260
rect 31163 10220 31208 10248
rect 31202 10208 31208 10220
rect 31260 10208 31266 10260
rect 33413 10251 33471 10257
rect 33413 10217 33425 10251
rect 33459 10248 33471 10251
rect 33502 10248 33508 10260
rect 33459 10220 33508 10248
rect 33459 10217 33471 10220
rect 33413 10211 33471 10217
rect 33502 10208 33508 10220
rect 33560 10208 33566 10260
rect 40494 10248 40500 10260
rect 40455 10220 40500 10248
rect 40494 10208 40500 10220
rect 40552 10208 40558 10260
rect 44453 10251 44511 10257
rect 44453 10217 44465 10251
rect 44499 10248 44511 10251
rect 46842 10248 46848 10260
rect 44499 10220 46848 10248
rect 44499 10217 44511 10220
rect 44453 10211 44511 10217
rect 46842 10208 46848 10220
rect 46900 10208 46906 10260
rect 47397 10251 47455 10257
rect 47397 10217 47409 10251
rect 47443 10248 47455 10251
rect 48498 10248 48504 10260
rect 47443 10220 48504 10248
rect 47443 10217 47455 10220
rect 47397 10211 47455 10217
rect 48498 10208 48504 10220
rect 48556 10208 48562 10260
rect 48590 10208 48596 10260
rect 48648 10248 48654 10260
rect 49421 10251 49479 10257
rect 49421 10248 49433 10251
rect 48648 10220 49433 10248
rect 48648 10208 48654 10220
rect 49421 10217 49433 10220
rect 49467 10217 49479 10251
rect 49421 10211 49479 10217
rect 49786 10208 49792 10260
rect 49844 10248 49850 10260
rect 50157 10251 50215 10257
rect 50157 10248 50169 10251
rect 49844 10220 50169 10248
rect 49844 10208 49850 10220
rect 50157 10217 50169 10220
rect 50203 10217 50215 10251
rect 50157 10211 50215 10217
rect 50246 10208 50252 10260
rect 50304 10248 50310 10260
rect 50304 10220 50752 10248
rect 50304 10208 50310 10220
rect 16114 10180 16120 10192
rect 9324 10152 12434 10180
rect 16027 10152 16120 10180
rect 9217 10143 9275 10149
rect 6546 10112 6552 10124
rect 6507 10084 6552 10112
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10112 7067 10115
rect 8110 10112 8116 10124
rect 7055 10084 8116 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 8110 10072 8116 10084
rect 8168 10072 8174 10124
rect 8938 10112 8944 10124
rect 8899 10084 8944 10112
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10112 9367 10115
rect 9490 10112 9496 10124
rect 9355 10084 9496 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 12406 10112 12434 10152
rect 16114 10140 16120 10152
rect 16172 10180 16178 10192
rect 16574 10180 16580 10192
rect 16172 10152 16580 10180
rect 16172 10140 16178 10152
rect 16574 10140 16580 10152
rect 16632 10140 16638 10192
rect 17957 10183 18015 10189
rect 17957 10149 17969 10183
rect 18003 10180 18015 10183
rect 18690 10180 18696 10192
rect 18003 10152 18696 10180
rect 18003 10149 18015 10152
rect 17957 10143 18015 10149
rect 13078 10112 13084 10124
rect 12406 10084 12756 10112
rect 13039 10084 13084 10112
rect 6917 10047 6975 10053
rect 6917 10013 6929 10047
rect 6963 10044 6975 10047
rect 8202 10044 8208 10056
rect 6963 10016 8208 10044
rect 6963 10013 6975 10016
rect 6917 10007 6975 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9030 10044 9036 10056
rect 8991 10016 9036 10044
rect 9030 10004 9036 10016
rect 9088 10004 9094 10056
rect 9122 10004 9128 10056
rect 9180 10044 9186 10056
rect 9217 10047 9275 10053
rect 9217 10044 9229 10047
rect 9180 10016 9229 10044
rect 9180 10004 9186 10016
rect 9217 10013 9229 10016
rect 9263 10013 9275 10047
rect 9217 10007 9275 10013
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9401 10007 9459 10013
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10044 11943 10047
rect 11931 10016 12434 10044
rect 11931 10013 11943 10016
rect 11885 10007 11943 10013
rect 8294 9936 8300 9988
rect 8352 9976 8358 9988
rect 9416 9976 9444 10007
rect 8352 9948 9444 9976
rect 8352 9936 8358 9948
rect 12406 9908 12434 10016
rect 12728 9976 12756 10084
rect 13078 10072 13084 10084
rect 13136 10072 13142 10124
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 15749 10115 15807 10121
rect 15749 10112 15761 10115
rect 15712 10084 15761 10112
rect 15712 10072 15718 10084
rect 15749 10081 15761 10084
rect 15795 10112 15807 10115
rect 16853 10115 16911 10121
rect 16853 10112 16865 10115
rect 15795 10084 16865 10112
rect 15795 10081 15807 10084
rect 15749 10075 15807 10081
rect 16853 10081 16865 10084
rect 16899 10081 16911 10115
rect 16853 10075 16911 10081
rect 16942 10072 16948 10124
rect 17000 10112 17006 10124
rect 17129 10115 17187 10121
rect 17129 10112 17141 10115
rect 17000 10084 17141 10112
rect 17000 10072 17006 10084
rect 17129 10081 17141 10084
rect 17175 10112 17187 10115
rect 18046 10112 18052 10124
rect 17175 10084 18052 10112
rect 17175 10081 17187 10084
rect 17129 10075 17187 10081
rect 18046 10072 18052 10084
rect 18104 10072 18110 10124
rect 12894 10044 12900 10056
rect 12855 10016 12900 10044
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 17221 10047 17279 10053
rect 17221 10013 17233 10047
rect 17267 10044 17279 10047
rect 18156 10044 18184 10152
rect 18690 10140 18696 10152
rect 18748 10180 18754 10192
rect 24949 10183 25007 10189
rect 18748 10152 22140 10180
rect 18748 10140 18754 10152
rect 19981 10115 20039 10121
rect 19981 10081 19993 10115
rect 20027 10112 20039 10115
rect 21542 10112 21548 10124
rect 20027 10084 21548 10112
rect 20027 10081 20039 10084
rect 19981 10075 20039 10081
rect 21542 10072 21548 10084
rect 21600 10072 21606 10124
rect 17267 10016 18184 10044
rect 20349 10047 20407 10053
rect 17267 10013 17279 10016
rect 17221 10007 17279 10013
rect 20349 10013 20361 10047
rect 20395 10044 20407 10047
rect 21174 10044 21180 10056
rect 20395 10016 21180 10044
rect 20395 10013 20407 10016
rect 20349 10007 20407 10013
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 22112 10053 22140 10152
rect 24949 10149 24961 10183
rect 24995 10149 25007 10183
rect 24949 10143 25007 10149
rect 24118 10072 24124 10124
rect 24176 10112 24182 10124
rect 24489 10115 24547 10121
rect 24489 10112 24501 10115
rect 24176 10084 24501 10112
rect 24176 10072 24182 10084
rect 24489 10081 24501 10084
rect 24535 10081 24547 10115
rect 24489 10075 24547 10081
rect 21269 10047 21327 10053
rect 21269 10013 21281 10047
rect 21315 10013 21327 10047
rect 21269 10007 21327 10013
rect 22097 10047 22155 10053
rect 22097 10013 22109 10047
rect 22143 10013 22155 10047
rect 22097 10007 22155 10013
rect 22373 10047 22431 10053
rect 22373 10013 22385 10047
rect 22419 10044 22431 10047
rect 24578 10044 24584 10056
rect 22419 10016 24584 10044
rect 22419 10013 22431 10016
rect 22373 10007 22431 10013
rect 12728 9948 13032 9976
rect 13004 9917 13032 9948
rect 19886 9936 19892 9988
rect 19944 9976 19950 9988
rect 20257 9979 20315 9985
rect 20257 9976 20269 9979
rect 19944 9948 20269 9976
rect 19944 9936 19950 9948
rect 20257 9945 20269 9948
rect 20303 9976 20315 9979
rect 21284 9976 21312 10007
rect 20303 9948 21312 9976
rect 22112 9976 22140 10007
rect 24578 10004 24584 10016
rect 24636 10004 24642 10056
rect 24964 10044 24992 10143
rect 29546 10140 29552 10192
rect 29604 10180 29610 10192
rect 34422 10180 34428 10192
rect 29604 10152 34428 10180
rect 29604 10140 29610 10152
rect 34422 10140 34428 10152
rect 34480 10140 34486 10192
rect 41230 10180 41236 10192
rect 34992 10152 41236 10180
rect 29178 10072 29184 10124
rect 29236 10112 29242 10124
rect 29917 10115 29975 10121
rect 29917 10112 29929 10115
rect 29236 10084 29929 10112
rect 29236 10072 29242 10084
rect 29917 10081 29929 10084
rect 29963 10112 29975 10115
rect 32122 10112 32128 10124
rect 29963 10084 31248 10112
rect 32083 10084 32128 10112
rect 29963 10081 29975 10084
rect 29917 10075 29975 10081
rect 25685 10047 25743 10053
rect 25685 10044 25697 10047
rect 24964 10016 25697 10044
rect 25685 10013 25697 10016
rect 25731 10044 25743 10047
rect 26418 10044 26424 10056
rect 25731 10016 26424 10044
rect 25731 10013 25743 10016
rect 25685 10007 25743 10013
rect 26418 10004 26424 10016
rect 26476 10004 26482 10056
rect 30374 10044 30380 10056
rect 30335 10016 30380 10044
rect 30374 10004 30380 10016
rect 30432 10004 30438 10056
rect 30650 10044 30656 10056
rect 30611 10016 30656 10044
rect 30650 10004 30656 10016
rect 30708 10044 30714 10056
rect 31110 10044 31116 10056
rect 30708 10016 31116 10044
rect 30708 10004 30714 10016
rect 31110 10004 31116 10016
rect 31168 10004 31174 10056
rect 31220 10044 31248 10084
rect 32122 10072 32128 10084
rect 32180 10072 32186 10124
rect 32582 10072 32588 10124
rect 32640 10112 32646 10124
rect 32769 10115 32827 10121
rect 32769 10112 32781 10115
rect 32640 10084 32781 10112
rect 32640 10072 32646 10084
rect 32769 10081 32781 10084
rect 32815 10081 32827 10115
rect 32769 10075 32827 10081
rect 32217 10047 32275 10053
rect 32217 10044 32229 10047
rect 31220 10016 32229 10044
rect 32217 10013 32229 10016
rect 32263 10044 32275 10047
rect 34992 10044 35020 10152
rect 41230 10140 41236 10152
rect 41288 10140 41294 10192
rect 46860 10180 46888 10208
rect 49142 10180 49148 10192
rect 46860 10152 49148 10180
rect 49142 10140 49148 10152
rect 49200 10140 49206 10192
rect 49510 10180 49516 10192
rect 49471 10152 49516 10180
rect 49510 10140 49516 10152
rect 49568 10140 49574 10192
rect 41414 10112 41420 10124
rect 37292 10084 41420 10112
rect 37292 10053 37320 10084
rect 41414 10072 41420 10084
rect 41472 10072 41478 10124
rect 43530 10072 43536 10124
rect 43588 10112 43594 10124
rect 43588 10084 45692 10112
rect 43588 10072 43594 10084
rect 32263 10016 35020 10044
rect 37277 10047 37335 10053
rect 32263 10013 32275 10016
rect 32217 10007 32275 10013
rect 37277 10013 37289 10047
rect 37323 10013 37335 10047
rect 37277 10007 37335 10013
rect 38102 10004 38108 10056
rect 38160 10044 38166 10056
rect 38197 10047 38255 10053
rect 38197 10044 38209 10047
rect 38160 10016 38209 10044
rect 38160 10004 38166 10016
rect 38197 10013 38209 10016
rect 38243 10044 38255 10047
rect 38746 10044 38752 10056
rect 38243 10016 38752 10044
rect 38243 10013 38255 10016
rect 38197 10007 38255 10013
rect 38746 10004 38752 10016
rect 38804 10004 38810 10056
rect 40034 10044 40040 10056
rect 39995 10016 40040 10044
rect 40034 10004 40040 10016
rect 40092 10004 40098 10056
rect 42705 10047 42763 10053
rect 40328 10016 41414 10044
rect 40328 9988 40356 10016
rect 22112 9948 23520 9976
rect 20303 9945 20315 9948
rect 20257 9939 20315 9945
rect 12529 9911 12587 9917
rect 12529 9908 12541 9911
rect 12406 9880 12541 9908
rect 12529 9877 12541 9880
rect 12575 9877 12587 9911
rect 12529 9871 12587 9877
rect 12989 9911 13047 9917
rect 12989 9877 13001 9911
rect 13035 9908 13047 9911
rect 14185 9911 14243 9917
rect 14185 9908 14197 9911
rect 13035 9880 14197 9908
rect 13035 9877 13047 9880
rect 12989 9871 13047 9877
rect 14185 9877 14197 9880
rect 14231 9908 14243 9911
rect 14550 9908 14556 9920
rect 14231 9880 14556 9908
rect 14231 9877 14243 9880
rect 14185 9871 14243 9877
rect 14550 9868 14556 9880
rect 14608 9868 14614 9920
rect 20070 9908 20076 9920
rect 20031 9880 20076 9908
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 20165 9911 20223 9917
rect 20165 9877 20177 9911
rect 20211 9908 20223 9911
rect 21358 9908 21364 9920
rect 20211 9880 21364 9908
rect 20211 9877 20223 9880
rect 20165 9871 20223 9877
rect 21358 9868 21364 9880
rect 21416 9868 21422 9920
rect 23492 9917 23520 9948
rect 26326 9936 26332 9988
rect 26384 9976 26390 9988
rect 27985 9979 28043 9985
rect 27985 9976 27997 9979
rect 26384 9948 27997 9976
rect 26384 9936 26390 9948
rect 27985 9945 27997 9948
rect 28031 9945 28043 9979
rect 28166 9976 28172 9988
rect 28127 9948 28172 9976
rect 27985 9939 28043 9945
rect 28166 9936 28172 9948
rect 28224 9936 28230 9988
rect 30561 9979 30619 9985
rect 30561 9945 30573 9979
rect 30607 9976 30619 9979
rect 31386 9976 31392 9988
rect 30607 9948 31392 9976
rect 30607 9945 30619 9948
rect 30561 9939 30619 9945
rect 31386 9936 31392 9948
rect 31444 9936 31450 9988
rect 39025 9979 39083 9985
rect 39025 9945 39037 9979
rect 39071 9976 39083 9979
rect 40310 9976 40316 9988
rect 39071 9948 40316 9976
rect 39071 9945 39083 9948
rect 39025 9939 39083 9945
rect 40310 9936 40316 9948
rect 40368 9936 40374 9988
rect 23477 9911 23535 9917
rect 23477 9877 23489 9911
rect 23523 9908 23535 9911
rect 24762 9908 24768 9920
rect 23523 9880 24768 9908
rect 23523 9877 23535 9880
rect 23477 9871 23535 9877
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 28626 9868 28632 9920
rect 28684 9908 28690 9920
rect 33502 9908 33508 9920
rect 28684 9880 33508 9908
rect 28684 9868 28690 9880
rect 33502 9868 33508 9880
rect 33560 9868 33566 9920
rect 33962 9908 33968 9920
rect 33923 9880 33968 9908
rect 33962 9868 33968 9880
rect 34020 9868 34026 9920
rect 36446 9868 36452 9920
rect 36504 9908 36510 9920
rect 37185 9911 37243 9917
rect 37185 9908 37197 9911
rect 36504 9880 37197 9908
rect 36504 9868 36510 9880
rect 37185 9877 37197 9880
rect 37231 9877 37243 9911
rect 39942 9908 39948 9920
rect 39903 9880 39948 9908
rect 37185 9871 37243 9877
rect 39942 9868 39948 9880
rect 40000 9868 40006 9920
rect 41386 9908 41414 10016
rect 42705 10013 42717 10047
rect 42751 10013 42763 10047
rect 42705 10007 42763 10013
rect 45189 10047 45247 10053
rect 45189 10013 45201 10047
rect 45235 10044 45247 10047
rect 45462 10044 45468 10056
rect 45235 10016 45468 10044
rect 45235 10013 45247 10016
rect 45189 10007 45247 10013
rect 42720 9908 42748 10007
rect 45462 10004 45468 10016
rect 45520 10004 45526 10056
rect 45664 10053 45692 10084
rect 46750 10072 46756 10124
rect 46808 10112 46814 10124
rect 48041 10115 48099 10121
rect 48041 10112 48053 10115
rect 46808 10084 48053 10112
rect 46808 10072 46814 10084
rect 48041 10081 48053 10084
rect 48087 10081 48099 10115
rect 49326 10112 49332 10124
rect 49287 10084 49332 10112
rect 48041 10075 48099 10081
rect 49326 10072 49332 10084
rect 49384 10072 49390 10124
rect 49786 10072 49792 10124
rect 49844 10112 49850 10124
rect 49970 10112 49976 10124
rect 49844 10084 49976 10112
rect 49844 10072 49850 10084
rect 49970 10072 49976 10084
rect 50028 10072 50034 10124
rect 50430 10072 50436 10124
rect 50488 10112 50494 10124
rect 50617 10115 50675 10121
rect 50488 10084 50533 10112
rect 50488 10072 50494 10084
rect 50617 10081 50629 10115
rect 50663 10112 50675 10115
rect 50724 10112 50752 10220
rect 50663 10084 50752 10112
rect 50663 10081 50675 10084
rect 50617 10075 50675 10081
rect 45649 10047 45707 10053
rect 45649 10013 45661 10047
rect 45695 10013 45707 10047
rect 45649 10007 45707 10013
rect 47026 10004 47032 10056
rect 47084 10044 47090 10056
rect 47213 10047 47271 10053
rect 47213 10044 47225 10047
rect 47084 10016 47225 10044
rect 47084 10004 47090 10016
rect 47213 10013 47225 10016
rect 47259 10013 47271 10047
rect 47213 10007 47271 10013
rect 47397 10047 47455 10053
rect 47397 10013 47409 10047
rect 47443 10044 47455 10047
rect 48222 10044 48228 10056
rect 47443 10016 48228 10044
rect 47443 10013 47455 10016
rect 47397 10007 47455 10013
rect 48222 10004 48228 10016
rect 48280 10004 48286 10056
rect 48317 10047 48375 10053
rect 48317 10013 48329 10047
rect 48363 10044 48375 10047
rect 49234 10044 49240 10056
rect 48363 10016 49240 10044
rect 48363 10013 48375 10016
rect 48317 10007 48375 10013
rect 49234 10004 49240 10016
rect 49292 10004 49298 10056
rect 49605 10047 49663 10053
rect 49605 10013 49617 10047
rect 49651 10013 49663 10047
rect 49988 10044 50016 10072
rect 50315 10047 50373 10053
rect 50315 10044 50327 10047
rect 49988 10016 50327 10044
rect 49605 10007 49663 10013
rect 50315 10013 50327 10016
rect 50361 10013 50373 10047
rect 50315 10007 50373 10013
rect 50525 10047 50583 10053
rect 50525 10013 50537 10047
rect 50571 10013 50583 10047
rect 50525 10007 50583 10013
rect 51169 10047 51227 10053
rect 51169 10013 51181 10047
rect 51215 10013 51227 10047
rect 51169 10007 51227 10013
rect 42978 9976 42984 9988
rect 42939 9948 42984 9976
rect 42978 9936 42984 9948
rect 43036 9936 43042 9988
rect 45741 9979 45799 9985
rect 45741 9976 45753 9979
rect 44206 9948 45753 9976
rect 45741 9945 45753 9948
rect 45787 9945 45799 9979
rect 45741 9939 45799 9945
rect 48590 9936 48596 9988
rect 48648 9976 48654 9988
rect 49620 9976 49648 10007
rect 48648 9948 49648 9976
rect 48648 9936 48654 9948
rect 49970 9936 49976 9988
rect 50028 9976 50034 9988
rect 50541 9976 50569 10007
rect 51184 9976 51212 10007
rect 50028 9948 50569 9976
rect 51046 9948 51212 9976
rect 50028 9936 50034 9948
rect 43622 9908 43628 9920
rect 41386 9880 43628 9908
rect 43622 9868 43628 9880
rect 43680 9868 43686 9920
rect 45002 9868 45008 9920
rect 45060 9908 45066 9920
rect 45097 9911 45155 9917
rect 45097 9908 45109 9911
rect 45060 9880 45109 9908
rect 45060 9868 45066 9880
rect 45097 9877 45109 9880
rect 45143 9877 45155 9911
rect 47578 9908 47584 9920
rect 47539 9880 47584 9908
rect 45097 9871 45155 9877
rect 47578 9868 47584 9880
rect 47636 9868 47642 9920
rect 49142 9868 49148 9920
rect 49200 9908 49206 9920
rect 51046 9908 51074 9948
rect 51258 9908 51264 9920
rect 49200 9880 51074 9908
rect 51219 9880 51264 9908
rect 49200 9868 49206 9880
rect 51258 9868 51264 9880
rect 51316 9868 51322 9920
rect 1104 9818 68816 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 68816 9818
rect 1104 9744 68816 9766
rect 8297 9707 8355 9713
rect 8297 9673 8309 9707
rect 8343 9704 8355 9707
rect 8386 9704 8392 9716
rect 8343 9676 8392 9704
rect 8343 9673 8355 9676
rect 8297 9667 8355 9673
rect 8386 9664 8392 9676
rect 8444 9704 8450 9716
rect 8938 9704 8944 9716
rect 8444 9676 8944 9704
rect 8444 9664 8450 9676
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 16114 9704 16120 9716
rect 16075 9676 16120 9704
rect 16114 9664 16120 9676
rect 16172 9664 16178 9716
rect 20349 9707 20407 9713
rect 20349 9673 20361 9707
rect 20395 9704 20407 9707
rect 20622 9704 20628 9716
rect 20395 9676 20628 9704
rect 20395 9673 20407 9676
rect 20349 9667 20407 9673
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 25958 9704 25964 9716
rect 25919 9676 25964 9704
rect 25958 9664 25964 9676
rect 26016 9664 26022 9716
rect 32306 9664 32312 9716
rect 32364 9704 32370 9716
rect 32585 9707 32643 9713
rect 32585 9704 32597 9707
rect 32364 9676 32597 9704
rect 32364 9664 32370 9676
rect 32585 9673 32597 9676
rect 32631 9673 32643 9707
rect 32585 9667 32643 9673
rect 33962 9664 33968 9716
rect 34020 9704 34026 9716
rect 38102 9704 38108 9716
rect 34020 9676 38108 9704
rect 34020 9664 34026 9676
rect 9030 9636 9036 9648
rect 8220 9608 9036 9636
rect 6638 9568 6644 9580
rect 6599 9540 6644 9568
rect 6638 9528 6644 9540
rect 6696 9528 6702 9580
rect 8220 9577 8248 9608
rect 9030 9596 9036 9608
rect 9088 9596 9094 9648
rect 15378 9596 15384 9648
rect 15436 9636 15442 9648
rect 15749 9639 15807 9645
rect 15749 9636 15761 9639
rect 15436 9608 15761 9636
rect 15436 9596 15442 9608
rect 15749 9605 15761 9608
rect 15795 9636 15807 9639
rect 16666 9636 16672 9648
rect 15795 9608 16068 9636
rect 16627 9608 16672 9636
rect 15795 9605 15807 9608
rect 15749 9599 15807 9605
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 9306 9568 9312 9580
rect 8527 9540 8984 9568
rect 9267 9540 9312 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 6546 9500 6552 9512
rect 6507 9472 6552 9500
rect 6546 9460 6552 9472
rect 6604 9460 6610 9512
rect 8956 9509 8984 9540
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 13173 9571 13231 9577
rect 13173 9568 13185 9571
rect 12768 9540 13185 9568
rect 12768 9528 12774 9540
rect 13173 9537 13185 9540
rect 13219 9537 13231 9571
rect 13446 9568 13452 9580
rect 13407 9540 13452 9568
rect 13173 9531 13231 9537
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 15654 9568 15660 9580
rect 15615 9540 15660 9568
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 15930 9568 15936 9580
rect 15891 9540 15936 9568
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 16040 9568 16068 9608
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 17221 9639 17279 9645
rect 17221 9605 17233 9639
rect 17267 9636 17279 9639
rect 17678 9636 17684 9648
rect 17267 9608 17684 9636
rect 17267 9605 17279 9608
rect 17221 9599 17279 9605
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 24578 9636 24584 9648
rect 24044 9608 24584 9636
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16040 9540 16865 9568
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 16945 9571 17003 9577
rect 16945 9537 16957 9571
rect 16991 9537 17003 9571
rect 16945 9531 17003 9537
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9537 17095 9571
rect 17037 9531 17095 9537
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9469 8999 9503
rect 8941 9463 8999 9469
rect 9401 9503 9459 9509
rect 9401 9469 9413 9503
rect 9447 9500 9459 9503
rect 10686 9500 10692 9512
rect 9447 9472 10692 9500
rect 9447 9469 9459 9472
rect 9401 9463 9459 9469
rect 10686 9460 10692 9472
rect 10744 9500 10750 9512
rect 10962 9500 10968 9512
rect 10744 9472 10968 9500
rect 10744 9460 10750 9472
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 13262 9500 13268 9512
rect 13223 9472 13268 9500
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 15672 9500 15700 9528
rect 16960 9500 16988 9531
rect 15672 9472 16988 9500
rect 7009 9435 7067 9441
rect 7009 9401 7021 9435
rect 7055 9432 7067 9435
rect 8294 9432 8300 9444
rect 7055 9404 8300 9432
rect 7055 9401 7067 9404
rect 7009 9395 7067 9401
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 8481 9435 8539 9441
rect 8481 9401 8493 9435
rect 8527 9432 8539 9435
rect 9122 9432 9128 9444
rect 8527 9404 9128 9432
rect 8527 9401 8539 9404
rect 8481 9395 8539 9401
rect 9122 9392 9128 9404
rect 9180 9392 9186 9444
rect 13630 9432 13636 9444
rect 13591 9404 13636 9432
rect 13630 9392 13636 9404
rect 13688 9392 13694 9444
rect 14734 9392 14740 9444
rect 14792 9432 14798 9444
rect 17052 9432 17080 9531
rect 20070 9528 20076 9580
rect 20128 9568 20134 9580
rect 20533 9571 20591 9577
rect 20533 9568 20545 9571
rect 20128 9540 20545 9568
rect 20128 9528 20134 9540
rect 20533 9537 20545 9540
rect 20579 9568 20591 9571
rect 20622 9568 20628 9580
rect 20579 9540 20628 9568
rect 20579 9537 20591 9540
rect 20533 9531 20591 9537
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 20717 9571 20775 9577
rect 20717 9537 20729 9571
rect 20763 9537 20775 9571
rect 20717 9531 20775 9537
rect 20809 9571 20867 9577
rect 20809 9537 20821 9571
rect 20855 9568 20867 9571
rect 20898 9568 20904 9580
rect 20855 9540 20904 9568
rect 20855 9537 20867 9540
rect 20809 9531 20867 9537
rect 20732 9500 20760 9531
rect 20898 9528 20904 9540
rect 20956 9528 20962 9580
rect 21910 9528 21916 9580
rect 21968 9568 21974 9580
rect 24044 9577 24072 9608
rect 24578 9596 24584 9608
rect 24636 9636 24642 9648
rect 30837 9639 30895 9645
rect 24636 9608 27752 9636
rect 24636 9596 24642 9608
rect 22281 9571 22339 9577
rect 22281 9568 22293 9571
rect 21968 9540 22293 9568
rect 21968 9528 21974 9540
rect 22281 9537 22293 9540
rect 22327 9537 22339 9571
rect 22281 9531 22339 9537
rect 24029 9571 24087 9577
rect 24029 9537 24041 9571
rect 24075 9537 24087 9571
rect 24029 9531 24087 9537
rect 20548 9472 20760 9500
rect 20548 9444 20576 9472
rect 21174 9460 21180 9512
rect 21232 9500 21238 9512
rect 21821 9503 21879 9509
rect 21821 9500 21833 9503
rect 21232 9472 21833 9500
rect 21232 9460 21238 9472
rect 21821 9469 21833 9472
rect 21867 9469 21879 9503
rect 21821 9463 21879 9469
rect 14792 9404 17080 9432
rect 14792 9392 14798 9404
rect 20530 9392 20536 9444
rect 20588 9392 20594 9444
rect 24044 9432 24072 9531
rect 25774 9528 25780 9580
rect 25832 9568 25838 9580
rect 27724 9577 27752 9608
rect 30837 9605 30849 9639
rect 30883 9636 30895 9639
rect 32122 9636 32128 9648
rect 30883 9608 32128 9636
rect 30883 9605 30895 9608
rect 30837 9599 30895 9605
rect 32122 9596 32128 9608
rect 32180 9596 32186 9648
rect 34256 9645 34284 9676
rect 38102 9664 38108 9676
rect 38160 9664 38166 9716
rect 40034 9664 40040 9716
rect 40092 9704 40098 9716
rect 40092 9676 42932 9704
rect 40092 9664 40098 9676
rect 34241 9639 34299 9645
rect 34241 9605 34253 9639
rect 34287 9605 34299 9639
rect 39942 9636 39948 9648
rect 39790 9608 39948 9636
rect 34241 9599 34299 9605
rect 39942 9596 39948 9608
rect 40000 9596 40006 9648
rect 40310 9596 40316 9648
rect 40368 9636 40374 9648
rect 40368 9608 40540 9636
rect 40368 9596 40374 9608
rect 26145 9571 26203 9577
rect 26145 9568 26157 9571
rect 25832 9540 26157 9568
rect 25832 9528 25838 9540
rect 26145 9537 26157 9540
rect 26191 9537 26203 9571
rect 26145 9531 26203 9537
rect 27709 9571 27767 9577
rect 27709 9537 27721 9571
rect 27755 9568 27767 9571
rect 28258 9568 28264 9580
rect 27755 9540 28264 9568
rect 27755 9537 27767 9540
rect 27709 9531 27767 9537
rect 28258 9528 28264 9540
rect 28316 9528 28322 9580
rect 29365 9571 29423 9577
rect 29365 9537 29377 9571
rect 29411 9568 29423 9571
rect 29822 9568 29828 9580
rect 29411 9540 29828 9568
rect 29411 9537 29423 9540
rect 29365 9531 29423 9537
rect 29822 9528 29828 9540
rect 29880 9568 29886 9580
rect 30745 9571 30803 9577
rect 30745 9568 30757 9571
rect 29880 9540 30757 9568
rect 29880 9528 29886 9540
rect 30745 9537 30757 9540
rect 30791 9568 30803 9571
rect 33318 9568 33324 9580
rect 30791 9540 33324 9568
rect 30791 9537 30803 9540
rect 30745 9531 30803 9537
rect 33318 9528 33324 9540
rect 33376 9528 33382 9580
rect 35253 9571 35311 9577
rect 35253 9537 35265 9571
rect 35299 9568 35311 9571
rect 35342 9568 35348 9580
rect 35299 9540 35348 9568
rect 35299 9537 35311 9540
rect 35253 9531 35311 9537
rect 35342 9528 35348 9540
rect 35400 9528 35406 9580
rect 40512 9577 40540 9608
rect 40972 9577 41000 9676
rect 42904 9636 42932 9676
rect 42978 9664 42984 9716
rect 43036 9704 43042 9716
rect 43036 9676 45416 9704
rect 43036 9664 43042 9676
rect 44174 9636 44180 9648
rect 42904 9608 44180 9636
rect 44174 9596 44180 9608
rect 44232 9596 44238 9648
rect 45388 9636 45416 9676
rect 49234 9664 49240 9716
rect 49292 9704 49298 9716
rect 49970 9704 49976 9716
rect 49292 9676 49976 9704
rect 49292 9664 49298 9676
rect 49970 9664 49976 9676
rect 50028 9664 50034 9716
rect 50157 9707 50215 9713
rect 50157 9673 50169 9707
rect 50203 9704 50215 9707
rect 50614 9704 50620 9716
rect 50203 9676 50620 9704
rect 50203 9673 50215 9676
rect 50157 9667 50215 9673
rect 50614 9664 50620 9676
rect 50672 9664 50678 9716
rect 47581 9639 47639 9645
rect 47581 9636 47593 9639
rect 45388 9608 47593 9636
rect 47581 9605 47593 9608
rect 47627 9605 47639 9639
rect 49418 9636 49424 9648
rect 47581 9599 47639 9605
rect 48884 9608 49424 9636
rect 35989 9571 36047 9577
rect 35989 9568 36001 9571
rect 35452 9540 36001 9568
rect 24486 9500 24492 9512
rect 24447 9472 24492 9500
rect 24486 9460 24492 9472
rect 24544 9460 24550 9512
rect 26234 9460 26240 9512
rect 26292 9500 26298 9512
rect 26421 9503 26479 9509
rect 26421 9500 26433 9503
rect 26292 9472 26433 9500
rect 26292 9460 26298 9472
rect 26421 9469 26433 9472
rect 26467 9500 26479 9503
rect 27982 9500 27988 9512
rect 26467 9472 26924 9500
rect 27895 9472 27988 9500
rect 26467 9469 26479 9472
rect 26421 9463 26479 9469
rect 22204 9404 24072 9432
rect 13449 9367 13507 9373
rect 13449 9333 13461 9367
rect 13495 9364 13507 9367
rect 13722 9364 13728 9376
rect 13495 9336 13728 9364
rect 13495 9333 13507 9336
rect 13449 9327 13507 9333
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 22204 9373 22232 9404
rect 22189 9367 22247 9373
rect 22189 9333 22201 9367
rect 22235 9333 22247 9367
rect 24118 9364 24124 9376
rect 24079 9336 24124 9364
rect 22189 9327 22247 9333
rect 24118 9324 24124 9336
rect 24176 9324 24182 9376
rect 26329 9367 26387 9373
rect 26329 9333 26341 9367
rect 26375 9364 26387 9367
rect 26418 9364 26424 9376
rect 26375 9336 26424 9364
rect 26375 9333 26387 9336
rect 26329 9327 26387 9333
rect 26418 9324 26424 9336
rect 26476 9324 26482 9376
rect 26896 9364 26924 9472
rect 27982 9460 27988 9472
rect 28040 9500 28046 9512
rect 29638 9500 29644 9512
rect 28040 9472 29644 9500
rect 28040 9460 28046 9472
rect 29638 9460 29644 9472
rect 29696 9460 29702 9512
rect 30926 9500 30932 9512
rect 30887 9472 30932 9500
rect 30926 9460 30932 9472
rect 30984 9460 30990 9512
rect 32582 9460 32588 9512
rect 32640 9500 32646 9512
rect 33413 9503 33471 9509
rect 33413 9500 33425 9503
rect 32640 9472 33425 9500
rect 32640 9460 32646 9472
rect 33413 9469 33425 9472
rect 33459 9469 33471 9503
rect 35452 9500 35480 9540
rect 35989 9537 36001 9540
rect 36035 9537 36047 9571
rect 35989 9531 36047 9537
rect 40497 9571 40555 9577
rect 40497 9537 40509 9571
rect 40543 9537 40555 9571
rect 40497 9531 40555 9537
rect 40957 9571 41015 9577
rect 40957 9537 40969 9571
rect 41003 9537 41015 9571
rect 40957 9531 41015 9537
rect 45002 9528 45008 9580
rect 45060 9528 45066 9580
rect 47857 9571 47915 9577
rect 47857 9537 47869 9571
rect 47903 9568 47915 9571
rect 48590 9568 48596 9580
rect 47903 9540 48596 9568
rect 47903 9537 47915 9540
rect 47857 9531 47915 9537
rect 48590 9528 48596 9540
rect 48648 9528 48654 9580
rect 48884 9577 48912 9608
rect 49418 9596 49424 9608
rect 49476 9636 49482 9648
rect 49878 9636 49884 9648
rect 49476 9608 49884 9636
rect 49476 9596 49482 9608
rect 49878 9596 49884 9608
rect 49936 9596 49942 9648
rect 48869 9571 48927 9577
rect 48869 9537 48881 9571
rect 48915 9537 48927 9571
rect 49142 9568 49148 9580
rect 49103 9540 49148 9568
rect 48869 9531 48927 9537
rect 49142 9528 49148 9540
rect 49200 9528 49206 9580
rect 49694 9528 49700 9580
rect 49752 9568 49758 9580
rect 49789 9571 49847 9577
rect 49789 9568 49801 9571
rect 49752 9540 49801 9568
rect 49752 9528 49758 9540
rect 49789 9537 49801 9540
rect 49835 9537 49847 9571
rect 49988 9568 50016 9664
rect 50246 9596 50252 9648
rect 50304 9636 50310 9648
rect 51258 9636 51264 9648
rect 50304 9608 51264 9636
rect 50304 9596 50310 9608
rect 51258 9596 51264 9608
rect 51316 9596 51322 9648
rect 50065 9571 50123 9577
rect 50065 9568 50077 9571
rect 49988 9540 50077 9568
rect 49789 9531 49847 9537
rect 50065 9537 50077 9540
rect 50111 9568 50123 9571
rect 50893 9571 50951 9577
rect 50893 9568 50905 9571
rect 50111 9540 50905 9568
rect 50111 9537 50123 9540
rect 50065 9531 50123 9537
rect 50893 9537 50905 9540
rect 50939 9568 50951 9571
rect 51721 9571 51779 9577
rect 51721 9568 51733 9571
rect 50939 9540 51733 9568
rect 50939 9537 50951 9540
rect 50893 9531 50951 9537
rect 51721 9537 51733 9540
rect 51767 9537 51779 9571
rect 51721 9531 51779 9537
rect 35710 9500 35716 9512
rect 33413 9463 33471 9469
rect 35084 9472 35480 9500
rect 35671 9472 35716 9500
rect 27062 9432 27068 9444
rect 26975 9404 27068 9432
rect 27062 9392 27068 9404
rect 27120 9432 27126 9444
rect 29917 9435 29975 9441
rect 29917 9432 29929 9435
rect 27120 9404 29929 9432
rect 27120 9392 27126 9404
rect 29917 9401 29929 9404
rect 29963 9432 29975 9435
rect 32401 9435 32459 9441
rect 32401 9432 32413 9435
rect 29963 9404 32413 9432
rect 29963 9401 29975 9404
rect 29917 9395 29975 9401
rect 32401 9401 32413 9404
rect 32447 9401 32459 9435
rect 32401 9395 32459 9401
rect 34422 9392 34428 9444
rect 34480 9432 34486 9444
rect 35084 9441 35112 9472
rect 35710 9460 35716 9472
rect 35768 9460 35774 9512
rect 40218 9500 40224 9512
rect 40179 9472 40224 9500
rect 40218 9460 40224 9472
rect 40276 9460 40282 9512
rect 43622 9500 43628 9512
rect 43583 9472 43628 9500
rect 43622 9460 43628 9472
rect 43680 9460 43686 9512
rect 43901 9503 43959 9509
rect 43901 9469 43913 9503
rect 43947 9500 43959 9503
rect 45373 9503 45431 9509
rect 43947 9472 45324 9500
rect 43947 9469 43959 9472
rect 43901 9463 43959 9469
rect 35069 9435 35127 9441
rect 35069 9432 35081 9435
rect 34480 9404 35081 9432
rect 34480 9392 34486 9404
rect 35069 9401 35081 9404
rect 35115 9401 35127 9435
rect 45296 9432 45324 9472
rect 45373 9469 45385 9503
rect 45419 9500 45431 9503
rect 46750 9500 46756 9512
rect 45419 9472 46756 9500
rect 45419 9469 45431 9472
rect 45373 9463 45431 9469
rect 46750 9460 46756 9472
rect 46808 9460 46814 9512
rect 47578 9500 47584 9512
rect 47539 9472 47584 9500
rect 47578 9460 47584 9472
rect 47636 9460 47642 9512
rect 49605 9503 49663 9509
rect 49605 9469 49617 9503
rect 49651 9500 49663 9503
rect 49878 9500 49884 9512
rect 49651 9472 49884 9500
rect 49651 9469 49663 9472
rect 49605 9463 49663 9469
rect 49878 9460 49884 9472
rect 49936 9460 49942 9512
rect 49973 9503 50031 9509
rect 49973 9469 49985 9503
rect 50019 9500 50031 9503
rect 50798 9500 50804 9512
rect 50019 9472 50804 9500
rect 50019 9469 50031 9472
rect 49973 9463 50031 9469
rect 50798 9460 50804 9472
rect 50856 9460 50862 9512
rect 50982 9500 50988 9512
rect 50943 9472 50988 9500
rect 50982 9460 50988 9472
rect 51040 9460 51046 9512
rect 48406 9432 48412 9444
rect 45296 9404 48412 9432
rect 35069 9395 35127 9401
rect 48406 9392 48412 9404
rect 48464 9392 48470 9444
rect 50246 9432 50252 9444
rect 49896 9404 50252 9432
rect 29086 9364 29092 9376
rect 26896 9336 29092 9364
rect 29086 9324 29092 9336
rect 29144 9324 29150 9376
rect 30374 9364 30380 9376
rect 30335 9336 30380 9364
rect 30374 9324 30380 9336
rect 30432 9324 30438 9376
rect 36722 9364 36728 9376
rect 36683 9336 36728 9364
rect 36722 9324 36728 9336
rect 36780 9324 36786 9376
rect 38749 9367 38807 9373
rect 38749 9333 38761 9367
rect 38795 9364 38807 9367
rect 39206 9364 39212 9376
rect 38795 9336 39212 9364
rect 38795 9333 38807 9336
rect 38749 9327 38807 9333
rect 39206 9324 39212 9336
rect 39264 9324 39270 9376
rect 40954 9324 40960 9376
rect 41012 9364 41018 9376
rect 41049 9367 41107 9373
rect 41049 9364 41061 9367
rect 41012 9336 41061 9364
rect 41012 9324 41018 9336
rect 41049 9333 41061 9336
rect 41095 9333 41107 9367
rect 47762 9364 47768 9376
rect 47723 9336 47768 9364
rect 41049 9327 41107 9333
rect 47762 9324 47768 9336
rect 47820 9324 47826 9376
rect 48774 9324 48780 9376
rect 48832 9364 48838 9376
rect 49896 9373 49924 9404
rect 50246 9392 50252 9404
rect 50304 9392 50310 9444
rect 50522 9392 50528 9444
rect 50580 9432 50586 9444
rect 51813 9435 51871 9441
rect 51813 9432 51825 9435
rect 50580 9404 51825 9432
rect 50580 9392 50586 9404
rect 51813 9401 51825 9404
rect 51859 9401 51871 9435
rect 51813 9395 51871 9401
rect 49881 9367 49939 9373
rect 49881 9364 49893 9367
rect 48832 9336 49893 9364
rect 48832 9324 48838 9336
rect 49881 9333 49893 9336
rect 49927 9333 49939 9367
rect 49881 9327 49939 9333
rect 50706 9324 50712 9376
rect 50764 9364 50770 9376
rect 50982 9364 50988 9376
rect 50764 9336 50988 9364
rect 50764 9324 50770 9336
rect 50982 9324 50988 9336
rect 51040 9364 51046 9376
rect 51261 9367 51319 9373
rect 51261 9364 51273 9367
rect 51040 9336 51273 9364
rect 51040 9324 51046 9336
rect 51261 9333 51273 9336
rect 51307 9333 51319 9367
rect 51261 9327 51319 9333
rect 1104 9274 68816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 65654 9274
rect 65706 9222 65718 9274
rect 65770 9222 65782 9274
rect 65834 9222 65846 9274
rect 65898 9222 65910 9274
rect 65962 9222 68816 9274
rect 1104 9200 68816 9222
rect 15749 9163 15807 9169
rect 15749 9129 15761 9163
rect 15795 9160 15807 9163
rect 15930 9160 15936 9172
rect 15795 9132 15936 9160
rect 15795 9129 15807 9132
rect 15749 9123 15807 9129
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 19334 9120 19340 9172
rect 19392 9160 19398 9172
rect 20349 9163 20407 9169
rect 20349 9160 20361 9163
rect 19392 9132 20361 9160
rect 19392 9120 19398 9132
rect 20349 9129 20361 9132
rect 20395 9129 20407 9163
rect 21542 9160 21548 9172
rect 21503 9132 21548 9160
rect 20349 9123 20407 9129
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 21910 9160 21916 9172
rect 21871 9132 21916 9160
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 26973 9163 27031 9169
rect 26973 9129 26985 9163
rect 27019 9160 27031 9163
rect 28074 9160 28080 9172
rect 27019 9132 28080 9160
rect 27019 9129 27031 9132
rect 26973 9123 27031 9129
rect 28074 9120 28080 9132
rect 28132 9160 28138 9172
rect 29638 9160 29644 9172
rect 28132 9132 29132 9160
rect 29599 9132 29644 9160
rect 28132 9120 28138 9132
rect 8110 9052 8116 9104
rect 8168 9092 8174 9104
rect 9585 9095 9643 9101
rect 9585 9092 9597 9095
rect 8168 9064 9597 9092
rect 8168 9052 8174 9064
rect 9585 9061 9597 9064
rect 9631 9061 9643 9095
rect 9585 9055 9643 9061
rect 14090 9052 14096 9104
rect 14148 9092 14154 9104
rect 15841 9095 15899 9101
rect 15841 9092 15853 9095
rect 14148 9064 15853 9092
rect 14148 9052 14154 9064
rect 15841 9061 15853 9064
rect 15887 9092 15899 9095
rect 16114 9092 16120 9104
rect 15887 9064 16120 9092
rect 15887 9061 15899 9064
rect 15841 9055 15899 9061
rect 16114 9052 16120 9064
rect 16172 9092 16178 9104
rect 27062 9092 27068 9104
rect 16172 9064 27068 9092
rect 16172 9052 16178 9064
rect 25332 9036 25360 9064
rect 27062 9052 27068 9064
rect 27120 9052 27126 9104
rect 9766 9024 9772 9036
rect 9727 8996 9772 9024
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 15378 9024 15384 9036
rect 14568 8996 15384 9024
rect 9585 8959 9643 8965
rect 9585 8925 9597 8959
rect 9631 8956 9643 8959
rect 9674 8956 9680 8968
rect 9631 8928 9680 8956
rect 9631 8925 9643 8928
rect 9585 8919 9643 8925
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 14568 8965 14596 8996
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 16482 8984 16488 9036
rect 16540 9024 16546 9036
rect 16945 9027 17003 9033
rect 16945 9024 16957 9027
rect 16540 8996 16957 9024
rect 16540 8984 16546 8996
rect 16945 8993 16957 8996
rect 16991 8993 17003 9027
rect 16945 8987 17003 8993
rect 20533 9027 20591 9033
rect 20533 8993 20545 9027
rect 20579 9024 20591 9027
rect 21818 9024 21824 9036
rect 20579 8996 21824 9024
rect 20579 8993 20591 8996
rect 20533 8987 20591 8993
rect 21818 8984 21824 8996
rect 21876 8984 21882 9036
rect 25314 9024 25320 9036
rect 25227 8996 25320 9024
rect 25314 8984 25320 8996
rect 25372 8984 25378 9036
rect 26145 9027 26203 9033
rect 26145 8993 26157 9027
rect 26191 9024 26203 9027
rect 26234 9024 26240 9036
rect 26191 8996 26240 9024
rect 26191 8993 26203 8996
rect 26145 8987 26203 8993
rect 26234 8984 26240 8996
rect 26292 8984 26298 9036
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14734 8956 14740 8968
rect 14695 8928 14740 8956
rect 14553 8919 14611 8925
rect 14734 8916 14740 8928
rect 14792 8916 14798 8968
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 14976 8928 15301 8956
rect 14976 8916 14982 8928
rect 15289 8925 15301 8928
rect 15335 8956 15347 8959
rect 17037 8959 17095 8965
rect 15335 8928 16804 8956
rect 15335 8925 15347 8928
rect 15289 8919 15347 8925
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 10008 8860 10053 8888
rect 10008 8848 10014 8860
rect 15470 8848 15476 8900
rect 15528 8888 15534 8900
rect 16209 8891 16267 8897
rect 16209 8888 16221 8891
rect 15528 8860 16221 8888
rect 15528 8848 15534 8860
rect 16209 8857 16221 8860
rect 16255 8888 16267 8891
rect 16482 8888 16488 8900
rect 16255 8860 16488 8888
rect 16255 8857 16267 8860
rect 16209 8851 16267 8857
rect 16482 8848 16488 8860
rect 16540 8848 16546 8900
rect 12250 8780 12256 8832
rect 12308 8820 12314 8832
rect 14553 8823 14611 8829
rect 14553 8820 14565 8823
rect 12308 8792 14565 8820
rect 12308 8780 12314 8792
rect 14553 8789 14565 8792
rect 14599 8789 14611 8823
rect 14553 8783 14611 8789
rect 15654 8780 15660 8832
rect 15712 8820 15718 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 15712 8792 16681 8820
rect 15712 8780 15718 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16776 8820 16804 8928
rect 17037 8925 17049 8959
rect 17083 8958 17095 8959
rect 17083 8956 17172 8958
rect 18230 8956 18236 8968
rect 17083 8930 18236 8956
rect 17083 8925 17095 8930
rect 17144 8928 18236 8930
rect 17037 8919 17095 8925
rect 18230 8916 18236 8928
rect 18288 8916 18294 8968
rect 20162 8916 20168 8968
rect 20220 8956 20226 8968
rect 20349 8959 20407 8965
rect 20349 8956 20361 8959
rect 20220 8928 20361 8956
rect 20220 8916 20226 8928
rect 20349 8925 20361 8928
rect 20395 8925 20407 8959
rect 20622 8956 20628 8968
rect 20583 8928 20628 8956
rect 20349 8919 20407 8925
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 22005 8959 22063 8965
rect 22005 8925 22017 8959
rect 22051 8925 22063 8959
rect 22005 8919 22063 8925
rect 22020 8888 22048 8919
rect 25406 8916 25412 8968
rect 25464 8916 25470 8968
rect 28353 8959 28411 8965
rect 28353 8925 28365 8959
rect 28399 8956 28411 8959
rect 28442 8956 28448 8968
rect 28399 8928 28448 8956
rect 28399 8925 28411 8928
rect 28353 8919 28411 8925
rect 28442 8916 28448 8928
rect 28500 8916 28506 8968
rect 28994 8956 29000 8968
rect 28955 8928 29000 8956
rect 28994 8916 29000 8928
rect 29052 8916 29058 8968
rect 29104 8956 29132 9132
rect 29638 9120 29644 9132
rect 29696 9120 29702 9172
rect 29730 9120 29736 9172
rect 29788 9160 29794 9172
rect 30009 9163 30067 9169
rect 30009 9160 30021 9163
rect 29788 9132 30021 9160
rect 29788 9120 29794 9132
rect 30009 9129 30021 9132
rect 30055 9129 30067 9163
rect 30009 9123 30067 9129
rect 31849 9163 31907 9169
rect 31849 9129 31861 9163
rect 31895 9160 31907 9163
rect 32122 9160 32128 9172
rect 31895 9132 32128 9160
rect 31895 9129 31907 9132
rect 31849 9123 31907 9129
rect 32122 9120 32128 9132
rect 32180 9120 32186 9172
rect 33413 9163 33471 9169
rect 33413 9129 33425 9163
rect 33459 9160 33471 9163
rect 34606 9160 34612 9172
rect 33459 9132 34612 9160
rect 33459 9129 33471 9132
rect 33413 9123 33471 9129
rect 34606 9120 34612 9132
rect 34664 9120 34670 9172
rect 36722 9120 36728 9172
rect 36780 9160 36786 9172
rect 46934 9160 46940 9172
rect 36780 9132 46940 9160
rect 36780 9120 36786 9132
rect 46934 9120 46940 9132
rect 46992 9120 46998 9172
rect 48866 9160 48872 9172
rect 48827 9132 48872 9160
rect 48866 9120 48872 9132
rect 48924 9120 48930 9172
rect 49326 9160 49332 9172
rect 49287 9132 49332 9160
rect 49326 9120 49332 9132
rect 49384 9120 49390 9172
rect 50062 9120 50068 9172
rect 50120 9160 50126 9172
rect 50157 9163 50215 9169
rect 50157 9160 50169 9163
rect 50120 9132 50169 9160
rect 50120 9120 50126 9132
rect 50157 9129 50169 9132
rect 50203 9129 50215 9163
rect 50157 9123 50215 9129
rect 50890 9120 50896 9172
rect 50948 9160 50954 9172
rect 51261 9163 51319 9169
rect 51261 9160 51273 9163
rect 50948 9132 51273 9160
rect 50948 9120 50954 9132
rect 51261 9129 51273 9132
rect 51307 9129 51319 9163
rect 51261 9123 51319 9129
rect 35802 9052 35808 9104
rect 35860 9052 35866 9104
rect 49418 9092 49424 9104
rect 47780 9064 49424 9092
rect 32861 9027 32919 9033
rect 32861 8993 32873 9027
rect 32907 9024 32919 9027
rect 35820 9024 35848 9052
rect 37185 9027 37243 9033
rect 37185 9024 37197 9027
rect 32907 8996 33548 9024
rect 35820 8996 37197 9024
rect 32907 8993 32919 8996
rect 32861 8987 32919 8993
rect 29549 8959 29607 8965
rect 29549 8956 29561 8959
rect 29104 8928 29561 8956
rect 29549 8925 29561 8928
rect 29595 8925 29607 8959
rect 29549 8919 29607 8925
rect 30469 8959 30527 8965
rect 30469 8925 30481 8959
rect 30515 8956 30527 8959
rect 33042 8956 33048 8968
rect 30515 8928 33048 8956
rect 30515 8925 30527 8928
rect 30469 8919 30527 8925
rect 33042 8916 33048 8928
rect 33100 8916 33106 8968
rect 33134 8916 33140 8968
rect 33192 8956 33198 8968
rect 33520 8965 33548 8996
rect 37185 8993 37197 8996
rect 37231 9024 37243 9027
rect 39945 9027 40003 9033
rect 39945 9024 39957 9027
rect 37231 8996 39957 9024
rect 37231 8993 37243 8996
rect 37185 8987 37243 8993
rect 39945 8993 39957 8996
rect 39991 9024 40003 9027
rect 40310 9024 40316 9036
rect 39991 8996 40316 9024
rect 39991 8993 40003 8996
rect 39945 8987 40003 8993
rect 40310 8984 40316 8996
rect 40368 8984 40374 9036
rect 47780 9033 47808 9064
rect 49418 9052 49424 9064
rect 49476 9052 49482 9104
rect 49694 9052 49700 9104
rect 49752 9092 49758 9104
rect 50798 9092 50804 9104
rect 49752 9064 50804 9092
rect 49752 9052 49758 9064
rect 50798 9052 50804 9064
rect 50856 9092 50862 9104
rect 50856 9064 51074 9092
rect 50856 9052 50862 9064
rect 47765 9027 47823 9033
rect 47765 8993 47777 9027
rect 47811 8993 47823 9027
rect 48958 9024 48964 9036
rect 48871 8996 48964 9024
rect 47765 8987 47823 8993
rect 48958 8984 48964 8996
rect 49016 8984 49022 9036
rect 49053 9027 49111 9033
rect 49053 8993 49065 9027
rect 49099 9024 49111 9027
rect 49099 8996 50568 9024
rect 49099 8993 49111 8996
rect 49053 8987 49111 8993
rect 33321 8959 33379 8965
rect 33321 8956 33333 8959
rect 33192 8928 33333 8956
rect 33192 8916 33198 8928
rect 33321 8925 33333 8928
rect 33367 8925 33379 8959
rect 33321 8919 33379 8925
rect 33505 8959 33563 8965
rect 33505 8925 33517 8959
rect 33551 8925 33563 8959
rect 44174 8956 44180 8968
rect 44135 8928 44180 8956
rect 33505 8919 33563 8925
rect 44174 8916 44180 8928
rect 44232 8916 44238 8968
rect 47946 8956 47952 8968
rect 47907 8928 47952 8956
rect 47946 8916 47952 8928
rect 48004 8916 48010 8968
rect 48593 8959 48651 8965
rect 48593 8925 48605 8959
rect 48639 8925 48651 8959
rect 48774 8956 48780 8968
rect 48735 8928 48780 8956
rect 48593 8919 48651 8925
rect 23474 8888 23480 8900
rect 17144 8860 20944 8888
rect 22020 8860 23480 8888
rect 17144 8820 17172 8860
rect 16776 8792 17172 8820
rect 17773 8823 17831 8829
rect 16669 8783 16727 8789
rect 17773 8789 17785 8823
rect 17819 8820 17831 8823
rect 18230 8820 18236 8832
rect 17819 8792 18236 8820
rect 17819 8789 17831 8792
rect 17773 8783 17831 8789
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 20806 8820 20812 8832
rect 20767 8792 20812 8820
rect 20806 8780 20812 8792
rect 20864 8780 20870 8832
rect 20916 8820 20944 8860
rect 23474 8848 23480 8860
rect 23532 8888 23538 8900
rect 27982 8888 27988 8900
rect 23532 8860 27988 8888
rect 23532 8848 23538 8860
rect 27982 8848 27988 8860
rect 28040 8848 28046 8900
rect 28108 8891 28166 8897
rect 28108 8857 28120 8891
rect 28154 8888 28166 8891
rect 28154 8860 28856 8888
rect 28154 8857 28166 8860
rect 28108 8851 28166 8857
rect 22094 8820 22100 8832
rect 20916 8792 22100 8820
rect 22094 8780 22100 8792
rect 22152 8820 22158 8832
rect 28828 8829 28856 8860
rect 30558 8848 30564 8900
rect 30616 8888 30622 8900
rect 30714 8891 30772 8897
rect 30714 8888 30726 8891
rect 30616 8860 30726 8888
rect 30616 8848 30622 8860
rect 30714 8857 30726 8860
rect 30760 8857 30772 8891
rect 30714 8851 30772 8857
rect 32306 8848 32312 8900
rect 32364 8888 32370 8900
rect 32493 8891 32551 8897
rect 32493 8888 32505 8891
rect 32364 8860 32505 8888
rect 32364 8848 32370 8860
rect 32493 8857 32505 8860
rect 32539 8857 32551 8891
rect 32493 8851 32551 8857
rect 32674 8848 32680 8900
rect 32732 8888 32738 8900
rect 33965 8891 34023 8897
rect 33965 8888 33977 8891
rect 32732 8860 33977 8888
rect 32732 8848 32738 8860
rect 33965 8857 33977 8860
rect 34011 8857 34023 8891
rect 33965 8851 34023 8857
rect 36446 8848 36452 8900
rect 36504 8848 36510 8900
rect 36906 8888 36912 8900
rect 36867 8860 36912 8888
rect 36906 8848 36912 8860
rect 36964 8848 36970 8900
rect 40221 8891 40279 8897
rect 40221 8857 40233 8891
rect 40267 8888 40279 8891
rect 40494 8888 40500 8900
rect 40267 8860 40500 8888
rect 40267 8857 40279 8860
rect 40221 8851 40279 8857
rect 40494 8848 40500 8860
rect 40552 8848 40558 8900
rect 40954 8848 40960 8900
rect 41012 8848 41018 8900
rect 47762 8848 47768 8900
rect 47820 8888 47826 8900
rect 48608 8888 48636 8919
rect 48774 8916 48780 8928
rect 48832 8916 48838 8968
rect 48976 8956 49004 8984
rect 50540 8968 50568 8996
rect 49602 8956 49608 8968
rect 48976 8928 49608 8956
rect 49602 8916 49608 8928
rect 49660 8956 49666 8968
rect 50341 8959 50399 8965
rect 50341 8956 50353 8959
rect 49660 8928 50353 8956
rect 49660 8916 49666 8928
rect 50341 8925 50353 8928
rect 50387 8925 50399 8959
rect 50522 8956 50528 8968
rect 50483 8928 50528 8956
rect 50341 8919 50399 8925
rect 50522 8916 50528 8928
rect 50580 8916 50586 8968
rect 50617 8959 50675 8965
rect 50617 8925 50629 8959
rect 50663 8956 50675 8959
rect 50890 8956 50896 8968
rect 50663 8928 50896 8956
rect 50663 8925 50675 8928
rect 50617 8919 50675 8925
rect 50890 8916 50896 8928
rect 50948 8916 50954 8968
rect 51046 8956 51074 9064
rect 51046 8928 51488 8956
rect 49510 8888 49516 8900
rect 47820 8860 49516 8888
rect 47820 8848 47826 8860
rect 49510 8848 49516 8860
rect 49568 8848 49574 8900
rect 50982 8848 50988 8900
rect 51040 8888 51046 8900
rect 51460 8897 51488 8928
rect 51229 8891 51287 8897
rect 51229 8888 51241 8891
rect 51040 8860 51241 8888
rect 51040 8848 51046 8860
rect 51229 8857 51241 8860
rect 51275 8857 51287 8891
rect 51229 8851 51287 8857
rect 51445 8891 51503 8897
rect 51445 8857 51457 8891
rect 51491 8857 51503 8891
rect 51445 8851 51503 8857
rect 22465 8823 22523 8829
rect 22465 8820 22477 8823
rect 22152 8792 22477 8820
rect 22152 8780 22158 8792
rect 22465 8789 22477 8792
rect 22511 8789 22523 8823
rect 22465 8783 22523 8789
rect 28813 8823 28871 8829
rect 28813 8789 28825 8823
rect 28859 8789 28871 8823
rect 35434 8820 35440 8832
rect 35395 8792 35440 8820
rect 28813 8783 28871 8789
rect 35434 8780 35440 8792
rect 35492 8780 35498 8832
rect 41690 8820 41696 8832
rect 41651 8792 41696 8820
rect 41690 8780 41696 8792
rect 41748 8780 41754 8832
rect 44266 8820 44272 8832
rect 44227 8792 44272 8820
rect 44266 8780 44272 8792
rect 44324 8780 44330 8832
rect 48133 8823 48191 8829
rect 48133 8789 48145 8823
rect 48179 8820 48191 8823
rect 48498 8820 48504 8832
rect 48179 8792 48504 8820
rect 48179 8789 48191 8792
rect 48133 8783 48191 8789
rect 48498 8780 48504 8792
rect 48556 8780 48562 8832
rect 50706 8780 50712 8832
rect 50764 8820 50770 8832
rect 51077 8823 51135 8829
rect 51077 8820 51089 8823
rect 50764 8792 51089 8820
rect 50764 8780 50770 8792
rect 51077 8789 51089 8792
rect 51123 8789 51135 8823
rect 51077 8783 51135 8789
rect 1104 8730 68816 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 68816 8730
rect 1104 8656 68816 8678
rect 6365 8619 6423 8625
rect 6365 8585 6377 8619
rect 6411 8585 6423 8619
rect 6365 8579 6423 8585
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 6380 8480 6408 8579
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 6733 8619 6791 8625
rect 6733 8616 6745 8619
rect 6696 8588 6745 8616
rect 6696 8576 6702 8588
rect 6733 8585 6745 8588
rect 6779 8585 6791 8619
rect 6733 8579 6791 8585
rect 6822 8576 6828 8628
rect 6880 8616 6886 8628
rect 7561 8619 7619 8625
rect 7561 8616 7573 8619
rect 6880 8588 7573 8616
rect 6880 8576 6886 8588
rect 7561 8585 7573 8588
rect 7607 8585 7619 8619
rect 7561 8579 7619 8585
rect 8757 8619 8815 8625
rect 8757 8585 8769 8619
rect 8803 8616 8815 8619
rect 9030 8616 9036 8628
rect 8803 8588 9036 8616
rect 8803 8585 8815 8588
rect 8757 8579 8815 8585
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 11609 8619 11667 8625
rect 11609 8585 11621 8619
rect 11655 8616 11667 8619
rect 14090 8616 14096 8628
rect 11655 8588 14096 8616
rect 11655 8585 11667 8588
rect 11609 8579 11667 8585
rect 9766 8548 9772 8560
rect 9727 8520 9772 8548
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 5491 8452 6408 8480
rect 9125 8483 9183 8489
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 9125 8449 9137 8483
rect 9171 8480 9183 8483
rect 9784 8480 9812 8508
rect 9171 8452 9812 8480
rect 10781 8483 10839 8489
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 7374 8412 7380 8424
rect 7055 8384 7380 8412
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 7374 8372 7380 8384
rect 7432 8412 7438 8424
rect 7926 8412 7932 8424
rect 7432 8384 7932 8412
rect 7432 8372 7438 8384
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 9217 8415 9275 8421
rect 9217 8381 9229 8415
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 9232 8344 9260 8375
rect 9582 8372 9588 8424
rect 9640 8412 9646 8424
rect 10152 8412 10180 8466
rect 10781 8449 10793 8483
rect 10827 8480 10839 8483
rect 11624 8480 11652 8579
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 21818 8616 21824 8628
rect 14200 8588 20760 8616
rect 21779 8588 21824 8616
rect 11974 8508 11980 8560
rect 12032 8548 12038 8560
rect 12032 8520 13768 8548
rect 12032 8508 12038 8520
rect 12342 8480 12348 8492
rect 10827 8452 11652 8480
rect 12303 8452 12348 8480
rect 10827 8449 10839 8452
rect 10781 8443 10839 8449
rect 12342 8440 12348 8452
rect 12400 8440 12406 8492
rect 13740 8489 13768 8520
rect 14200 8489 14228 8588
rect 14553 8551 14611 8557
rect 14553 8517 14565 8551
rect 14599 8548 14611 8551
rect 16114 8548 16120 8560
rect 14599 8520 15424 8548
rect 16075 8520 16120 8548
rect 14599 8517 14611 8520
rect 14553 8511 14611 8517
rect 15396 8492 15424 8520
rect 16114 8508 16120 8520
rect 16172 8508 16178 8560
rect 17862 8548 17868 8560
rect 16684 8520 17868 8548
rect 13725 8483 13783 8489
rect 13725 8449 13737 8483
rect 13771 8480 13783 8483
rect 14185 8483 14243 8489
rect 14185 8480 14197 8483
rect 13771 8452 14197 8480
rect 13771 8449 13783 8452
rect 13725 8443 13783 8449
rect 14185 8449 14197 8452
rect 14231 8449 14243 8483
rect 14185 8443 14243 8449
rect 14339 8483 14397 8489
rect 14339 8449 14351 8483
rect 14385 8480 14397 8483
rect 14734 8480 14740 8492
rect 14385 8452 14740 8480
rect 14385 8449 14397 8452
rect 14339 8443 14397 8449
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 15378 8480 15384 8492
rect 15339 8452 15384 8480
rect 15378 8440 15384 8452
rect 15436 8440 15442 8492
rect 16574 8440 16580 8492
rect 16632 8480 16638 8492
rect 16684 8489 16712 8520
rect 17862 8508 17868 8520
rect 17920 8508 17926 8560
rect 20349 8551 20407 8557
rect 20349 8517 20361 8551
rect 20395 8548 20407 8551
rect 20622 8548 20628 8560
rect 20395 8520 20628 8548
rect 20395 8517 20407 8520
rect 20349 8511 20407 8517
rect 20622 8508 20628 8520
rect 20680 8508 20686 8560
rect 16942 8489 16948 8492
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 16632 8452 16681 8480
rect 16632 8440 16638 8452
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 16936 8443 16948 8489
rect 17000 8480 17006 8492
rect 17000 8452 17036 8480
rect 16942 8440 16948 8443
rect 17000 8440 17006 8452
rect 20162 8440 20168 8492
rect 20220 8480 20226 8492
rect 20732 8480 20760 8588
rect 21818 8576 21824 8588
rect 21876 8576 21882 8628
rect 25774 8616 25780 8628
rect 25735 8588 25780 8616
rect 25774 8576 25780 8588
rect 25832 8576 25838 8628
rect 26326 8616 26332 8628
rect 26287 8588 26332 8616
rect 26326 8576 26332 8588
rect 26384 8576 26390 8628
rect 27617 8619 27675 8625
rect 27617 8585 27629 8619
rect 27663 8616 27675 8619
rect 27982 8616 27988 8628
rect 27663 8588 27988 8616
rect 27663 8585 27675 8588
rect 27617 8579 27675 8585
rect 27982 8576 27988 8588
rect 28040 8576 28046 8628
rect 28077 8619 28135 8625
rect 28077 8585 28089 8619
rect 28123 8616 28135 8619
rect 28994 8616 29000 8628
rect 28123 8588 29000 8616
rect 28123 8585 28135 8588
rect 28077 8579 28135 8585
rect 28994 8576 29000 8588
rect 29052 8576 29058 8628
rect 29733 8619 29791 8625
rect 29733 8585 29745 8619
rect 29779 8616 29791 8619
rect 29822 8616 29828 8628
rect 29779 8588 29828 8616
rect 29779 8585 29791 8588
rect 29733 8579 29791 8585
rect 29822 8576 29828 8588
rect 29880 8576 29886 8628
rect 30377 8619 30435 8625
rect 30377 8585 30389 8619
rect 30423 8616 30435 8619
rect 31202 8616 31208 8628
rect 30423 8588 31208 8616
rect 30423 8585 30435 8588
rect 30377 8579 30435 8585
rect 31202 8576 31208 8588
rect 31260 8576 31266 8628
rect 31938 8576 31944 8628
rect 31996 8616 32002 8628
rect 32125 8619 32183 8625
rect 32125 8616 32137 8619
rect 31996 8588 32137 8616
rect 31996 8576 32002 8588
rect 32125 8585 32137 8588
rect 32171 8616 32183 8619
rect 33042 8616 33048 8628
rect 32171 8588 33048 8616
rect 32171 8585 32183 8588
rect 32125 8579 32183 8585
rect 33042 8576 33048 8588
rect 33100 8576 33106 8628
rect 36081 8619 36139 8625
rect 36081 8585 36093 8619
rect 36127 8616 36139 8619
rect 36906 8616 36912 8628
rect 36127 8588 36912 8616
rect 36127 8585 36139 8588
rect 36081 8579 36139 8585
rect 36906 8576 36912 8588
rect 36964 8576 36970 8628
rect 40218 8576 40224 8628
rect 40276 8616 40282 8628
rect 40405 8619 40463 8625
rect 40405 8616 40417 8619
rect 40276 8588 40417 8616
rect 40276 8576 40282 8588
rect 40405 8585 40417 8588
rect 40451 8585 40463 8619
rect 40405 8579 40463 8585
rect 40494 8576 40500 8628
rect 40552 8616 40558 8628
rect 40865 8619 40923 8625
rect 40865 8616 40877 8619
rect 40552 8588 40877 8616
rect 40552 8576 40558 8588
rect 40865 8585 40877 8588
rect 40911 8585 40923 8619
rect 40865 8579 40923 8585
rect 43533 8619 43591 8625
rect 43533 8585 43545 8619
rect 43579 8585 43591 8619
rect 43533 8579 43591 8585
rect 24857 8551 24915 8557
rect 24857 8548 24869 8551
rect 22112 8520 24869 8548
rect 22112 8492 22140 8520
rect 24857 8517 24869 8520
rect 24903 8548 24915 8551
rect 32674 8548 32680 8560
rect 24903 8520 25452 8548
rect 24903 8517 24915 8520
rect 24857 8511 24915 8517
rect 22094 8480 22100 8492
rect 20220 8452 20576 8480
rect 20732 8452 21956 8480
rect 22055 8452 22100 8480
rect 20220 8440 20226 8452
rect 12250 8412 12256 8424
rect 9640 8384 10180 8412
rect 12211 8384 12256 8412
rect 9640 8372 9646 8384
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 12710 8412 12716 8424
rect 12671 8384 12716 8412
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 15654 8412 15660 8424
rect 15519 8384 15660 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 19521 8415 19579 8421
rect 19521 8381 19533 8415
rect 19567 8412 19579 8415
rect 20438 8412 20444 8424
rect 19567 8384 20444 8412
rect 19567 8381 19579 8384
rect 19521 8375 19579 8381
rect 20438 8372 20444 8384
rect 20496 8372 20502 8424
rect 20548 8421 20576 8452
rect 20533 8415 20591 8421
rect 20533 8381 20545 8415
rect 20579 8381 20591 8415
rect 20533 8375 20591 8381
rect 20622 8372 20628 8424
rect 20680 8412 20686 8424
rect 21821 8415 21879 8421
rect 21821 8412 21833 8415
rect 20680 8384 21833 8412
rect 20680 8372 20686 8384
rect 21821 8381 21833 8384
rect 21867 8381 21879 8415
rect 21821 8375 21879 8381
rect 9674 8344 9680 8356
rect 9232 8316 9680 8344
rect 9674 8304 9680 8316
rect 9732 8344 9738 8356
rect 10778 8344 10784 8356
rect 9732 8316 10784 8344
rect 9732 8304 9738 8316
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 15013 8347 15071 8353
rect 15013 8344 15025 8347
rect 13780 8316 15025 8344
rect 13780 8304 13786 8316
rect 15013 8313 15025 8316
rect 15059 8313 15071 8347
rect 18046 8344 18052 8356
rect 18007 8316 18052 8344
rect 15013 8307 15071 8313
rect 18046 8304 18052 8316
rect 18104 8304 18110 8356
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 19981 8347 20039 8353
rect 19981 8344 19993 8347
rect 19300 8316 19993 8344
rect 19300 8304 19306 8316
rect 19981 8313 19993 8316
rect 20027 8313 20039 8347
rect 21928 8344 21956 8452
rect 22094 8440 22100 8452
rect 22152 8440 22158 8492
rect 22646 8480 22652 8492
rect 22607 8452 22652 8480
rect 22646 8440 22652 8452
rect 22704 8440 22710 8492
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8449 22891 8483
rect 23290 8480 23296 8492
rect 23251 8452 23296 8480
rect 22833 8443 22891 8449
rect 22848 8412 22876 8443
rect 23290 8440 23296 8452
rect 23348 8440 23354 8492
rect 23474 8480 23480 8492
rect 23435 8452 23480 8480
rect 23474 8440 23480 8452
rect 23532 8440 23538 8492
rect 25314 8480 25320 8492
rect 25275 8452 25320 8480
rect 25314 8440 25320 8452
rect 25372 8440 25378 8492
rect 25424 8480 25452 8520
rect 26252 8520 32680 8548
rect 26252 8489 26280 8520
rect 32674 8508 32680 8520
rect 32732 8508 32738 8560
rect 35434 8548 35440 8560
rect 34164 8520 35440 8548
rect 26237 8483 26295 8489
rect 26237 8480 26249 8483
rect 25424 8452 26249 8480
rect 26237 8449 26249 8452
rect 26283 8449 26295 8483
rect 26237 8443 26295 8449
rect 26326 8440 26332 8492
rect 26384 8480 26390 8492
rect 26421 8483 26479 8489
rect 26421 8480 26433 8483
rect 26384 8452 26433 8480
rect 26384 8440 26390 8452
rect 26421 8449 26433 8452
rect 26467 8449 26479 8483
rect 26421 8443 26479 8449
rect 27709 8483 27767 8489
rect 27709 8449 27721 8483
rect 27755 8480 27767 8483
rect 28258 8480 28264 8492
rect 27755 8452 28264 8480
rect 27755 8449 27767 8452
rect 27709 8443 27767 8449
rect 28258 8440 28264 8452
rect 28316 8440 28322 8492
rect 28799 8484 28857 8489
rect 28799 8483 28948 8484
rect 28460 8452 28764 8480
rect 23385 8415 23443 8421
rect 23385 8412 23397 8415
rect 22848 8384 23397 8412
rect 23385 8381 23397 8384
rect 23431 8381 23443 8415
rect 24946 8412 24952 8424
rect 23385 8375 23443 8381
rect 24228 8384 24952 8412
rect 24228 8344 24256 8384
rect 24946 8372 24952 8384
rect 25004 8412 25010 8424
rect 25774 8412 25780 8424
rect 25004 8384 25780 8412
rect 25004 8372 25010 8384
rect 25774 8372 25780 8384
rect 25832 8372 25838 8424
rect 27246 8372 27252 8424
rect 27304 8412 27310 8424
rect 27525 8415 27583 8421
rect 27525 8412 27537 8415
rect 27304 8384 27537 8412
rect 27304 8372 27310 8384
rect 27525 8381 27537 8384
rect 27571 8412 27583 8415
rect 28460 8412 28488 8452
rect 27571 8384 28488 8412
rect 28629 8415 28687 8421
rect 27571 8381 27583 8384
rect 27525 8375 27583 8381
rect 28629 8381 28641 8415
rect 28675 8381 28687 8415
rect 28736 8412 28764 8452
rect 28799 8449 28811 8483
rect 28845 8480 28948 8483
rect 29086 8480 29092 8492
rect 28845 8456 29092 8480
rect 28845 8449 28857 8456
rect 28920 8452 29092 8456
rect 28799 8443 28857 8449
rect 29086 8440 29092 8452
rect 29144 8440 29150 8492
rect 29638 8480 29644 8492
rect 29599 8452 29644 8480
rect 29638 8440 29644 8452
rect 29696 8440 29702 8492
rect 32306 8480 32312 8492
rect 32364 8489 32370 8492
rect 32364 8483 32397 8489
rect 31496 8452 32312 8480
rect 30926 8412 30932 8424
rect 28736 8384 30932 8412
rect 28629 8375 28687 8381
rect 21928 8316 24256 8344
rect 24305 8347 24363 8353
rect 19981 8307 20039 8313
rect 24305 8313 24317 8347
rect 24351 8344 24363 8347
rect 24394 8344 24400 8356
rect 24351 8316 24400 8344
rect 24351 8313 24363 8316
rect 24305 8307 24363 8313
rect 24394 8304 24400 8316
rect 24452 8344 24458 8356
rect 24452 8316 25544 8344
rect 24452 8304 24458 8316
rect 5261 8279 5319 8285
rect 5261 8245 5273 8279
rect 5307 8276 5319 8279
rect 5350 8276 5356 8288
rect 5307 8248 5356 8276
rect 5307 8245 5319 8248
rect 5261 8239 5319 8245
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 21910 8236 21916 8288
rect 21968 8276 21974 8288
rect 22005 8279 22063 8285
rect 22005 8276 22017 8279
rect 21968 8248 22017 8276
rect 21968 8236 21974 8248
rect 22005 8245 22017 8248
rect 22051 8245 22063 8279
rect 22005 8239 22063 8245
rect 22833 8279 22891 8285
rect 22833 8245 22845 8279
rect 22879 8276 22891 8279
rect 23014 8276 23020 8288
rect 22879 8248 23020 8276
rect 22879 8245 22891 8248
rect 22833 8239 22891 8245
rect 23014 8236 23020 8248
rect 23072 8236 23078 8288
rect 25406 8276 25412 8288
rect 25367 8248 25412 8276
rect 25406 8236 25412 8248
rect 25464 8236 25470 8288
rect 25516 8276 25544 8316
rect 26418 8304 26424 8356
rect 26476 8344 26482 8356
rect 28166 8344 28172 8356
rect 26476 8316 28172 8344
rect 26476 8304 26482 8316
rect 28166 8304 28172 8316
rect 28224 8344 28230 8356
rect 28644 8344 28672 8375
rect 30926 8372 30932 8384
rect 30984 8372 30990 8424
rect 31113 8415 31171 8421
rect 31113 8381 31125 8415
rect 31159 8412 31171 8415
rect 31294 8412 31300 8424
rect 31159 8384 31300 8412
rect 31159 8381 31171 8384
rect 31113 8375 31171 8381
rect 31294 8372 31300 8384
rect 31352 8412 31358 8424
rect 31496 8412 31524 8452
rect 32306 8440 32312 8452
rect 32385 8449 32397 8483
rect 32364 8443 32397 8449
rect 32364 8440 32370 8443
rect 32490 8440 32496 8492
rect 32548 8480 32554 8492
rect 34164 8489 34192 8520
rect 35434 8508 35440 8520
rect 35492 8508 35498 8560
rect 41690 8548 41696 8560
rect 41064 8520 41696 8548
rect 33137 8483 33195 8489
rect 32548 8452 32593 8480
rect 32548 8440 32554 8452
rect 33137 8449 33149 8483
rect 33183 8449 33195 8483
rect 33137 8443 33195 8449
rect 34149 8483 34207 8489
rect 34149 8449 34161 8483
rect 34195 8449 34207 8483
rect 34149 8443 34207 8449
rect 34425 8483 34483 8489
rect 34425 8449 34437 8483
rect 34471 8449 34483 8483
rect 34425 8443 34483 8449
rect 34609 8483 34667 8489
rect 34609 8449 34621 8483
rect 34655 8480 34667 8483
rect 35345 8483 35403 8489
rect 35345 8480 35357 8483
rect 34655 8452 35357 8480
rect 34655 8449 34667 8452
rect 34609 8443 34667 8449
rect 35345 8449 35357 8452
rect 35391 8449 35403 8483
rect 35345 8443 35403 8449
rect 39669 8483 39727 8489
rect 39669 8449 39681 8483
rect 39715 8480 39727 8483
rect 40034 8480 40040 8492
rect 39715 8452 40040 8480
rect 39715 8449 39727 8452
rect 39669 8443 39727 8449
rect 33152 8412 33180 8443
rect 31352 8384 31524 8412
rect 31588 8384 33180 8412
rect 31352 8372 31358 8384
rect 28224 8316 28672 8344
rect 29089 8347 29147 8353
rect 28224 8304 28230 8316
rect 29089 8313 29101 8347
rect 29135 8344 29147 8347
rect 30650 8344 30656 8356
rect 29135 8316 30656 8344
rect 29135 8313 29147 8316
rect 29089 8307 29147 8313
rect 30650 8304 30656 8316
rect 30708 8304 30714 8356
rect 31588 8353 31616 8384
rect 33594 8372 33600 8424
rect 33652 8412 33658 8424
rect 34440 8412 34468 8443
rect 40034 8440 40040 8452
rect 40092 8440 40098 8492
rect 41064 8489 41092 8520
rect 41690 8508 41696 8520
rect 41748 8508 41754 8560
rect 40129 8483 40187 8489
rect 40129 8449 40141 8483
rect 40175 8480 40187 8483
rect 41049 8483 41107 8489
rect 40175 8452 40356 8480
rect 40175 8449 40187 8452
rect 40129 8443 40187 8449
rect 33652 8384 34468 8412
rect 35069 8415 35127 8421
rect 33652 8372 33658 8384
rect 35069 8381 35081 8415
rect 35115 8381 35127 8415
rect 35069 8375 35127 8381
rect 31573 8347 31631 8353
rect 31573 8313 31585 8347
rect 31619 8313 31631 8347
rect 31573 8307 31631 8313
rect 29546 8276 29552 8288
rect 25516 8248 29552 8276
rect 29546 8236 29552 8248
rect 29604 8236 29610 8288
rect 32950 8276 32956 8288
rect 32911 8248 32956 8276
rect 32950 8236 32956 8248
rect 33008 8236 33014 8288
rect 34238 8276 34244 8288
rect 34199 8248 34244 8276
rect 34238 8236 34244 8248
rect 34296 8236 34302 8288
rect 34698 8236 34704 8288
rect 34756 8276 34762 8288
rect 35084 8276 35112 8375
rect 40218 8344 40224 8356
rect 40179 8316 40224 8344
rect 40218 8304 40224 8316
rect 40276 8304 40282 8356
rect 35710 8276 35716 8288
rect 34756 8248 35716 8276
rect 34756 8236 34762 8248
rect 35710 8236 35716 8248
rect 35768 8236 35774 8288
rect 39574 8276 39580 8288
rect 39535 8248 39580 8276
rect 39574 8236 39580 8248
rect 39632 8236 39638 8288
rect 40328 8276 40356 8452
rect 41049 8449 41061 8483
rect 41095 8449 41107 8483
rect 41049 8443 41107 8449
rect 41325 8483 41383 8489
rect 41325 8449 41337 8483
rect 41371 8449 41383 8483
rect 41325 8443 41383 8449
rect 42705 8483 42763 8489
rect 42705 8449 42717 8483
rect 42751 8480 42763 8483
rect 43254 8480 43260 8492
rect 42751 8452 43260 8480
rect 42751 8449 42763 8452
rect 42705 8443 42763 8449
rect 40405 8415 40463 8421
rect 40405 8381 40417 8415
rect 40451 8412 40463 8415
rect 40954 8412 40960 8424
rect 40451 8384 40960 8412
rect 40451 8381 40463 8384
rect 40405 8375 40463 8381
rect 40954 8372 40960 8384
rect 41012 8372 41018 8424
rect 41340 8412 41368 8443
rect 43254 8440 43260 8452
rect 43312 8480 43318 8492
rect 43548 8480 43576 8579
rect 43714 8576 43720 8628
rect 43772 8616 43778 8628
rect 50154 8616 50160 8628
rect 43772 8588 45324 8616
rect 50115 8588 50160 8616
rect 43772 8576 43778 8588
rect 44266 8508 44272 8560
rect 44324 8508 44330 8560
rect 45296 8489 45324 8588
rect 50154 8576 50160 8588
rect 50212 8576 50218 8628
rect 50325 8619 50383 8625
rect 50325 8616 50337 8619
rect 50264 8588 50337 8616
rect 48866 8508 48872 8560
rect 48924 8548 48930 8560
rect 49237 8551 49295 8557
rect 49237 8548 49249 8551
rect 48924 8520 49249 8548
rect 48924 8508 48930 8520
rect 49237 8517 49249 8520
rect 49283 8517 49295 8551
rect 49237 8511 49295 8517
rect 49326 8508 49332 8560
rect 49384 8548 49390 8560
rect 50264 8548 50292 8588
rect 50325 8585 50337 8588
rect 50371 8616 50383 8619
rect 50890 8616 50896 8628
rect 50371 8588 50896 8616
rect 50371 8585 50383 8588
rect 50325 8579 50383 8585
rect 50890 8576 50896 8588
rect 50948 8576 50954 8628
rect 49384 8520 50292 8548
rect 50525 8551 50583 8557
rect 49384 8508 49390 8520
rect 50525 8517 50537 8551
rect 50571 8548 50583 8551
rect 50798 8548 50804 8560
rect 50571 8520 50804 8548
rect 50571 8517 50583 8520
rect 50525 8511 50583 8517
rect 50798 8508 50804 8520
rect 50856 8508 50862 8560
rect 43312 8452 43576 8480
rect 45281 8483 45339 8489
rect 43312 8440 43318 8452
rect 45281 8449 45293 8483
rect 45327 8449 45339 8483
rect 45281 8443 45339 8449
rect 48314 8440 48320 8492
rect 48372 8480 48378 8492
rect 48501 8483 48559 8489
rect 48501 8480 48513 8483
rect 48372 8452 48513 8480
rect 48372 8440 48378 8452
rect 48501 8449 48513 8452
rect 48547 8480 48559 8483
rect 48958 8480 48964 8492
rect 48547 8452 48964 8480
rect 48547 8449 48559 8452
rect 48501 8443 48559 8449
rect 48958 8440 48964 8452
rect 49016 8440 49022 8492
rect 49418 8480 49424 8492
rect 49379 8452 49424 8480
rect 49418 8440 49424 8452
rect 49476 8440 49482 8492
rect 49513 8483 49571 8489
rect 49513 8449 49525 8483
rect 49559 8480 49571 8483
rect 49694 8480 49700 8492
rect 49559 8452 49700 8480
rect 49559 8449 49571 8452
rect 49513 8443 49571 8449
rect 49694 8440 49700 8452
rect 49752 8440 49758 8492
rect 41782 8412 41788 8424
rect 41340 8384 41788 8412
rect 41782 8372 41788 8384
rect 41840 8412 41846 8424
rect 42613 8415 42671 8421
rect 42613 8412 42625 8415
rect 41840 8384 42625 8412
rect 41840 8372 41846 8384
rect 42613 8381 42625 8384
rect 42659 8381 42671 8415
rect 45005 8415 45063 8421
rect 45005 8412 45017 8415
rect 42613 8375 42671 8381
rect 43088 8384 45017 8412
rect 41138 8344 41144 8356
rect 41099 8316 41144 8344
rect 41138 8304 41144 8316
rect 41196 8304 41202 8356
rect 41230 8304 41236 8356
rect 41288 8344 41294 8356
rect 43088 8353 43116 8384
rect 45005 8381 45017 8384
rect 45051 8381 45063 8415
rect 45005 8375 45063 8381
rect 48590 8372 48596 8424
rect 48648 8412 48654 8424
rect 48777 8415 48835 8421
rect 48777 8412 48789 8415
rect 48648 8384 48789 8412
rect 48648 8372 48654 8384
rect 48777 8381 48789 8384
rect 48823 8412 48835 8415
rect 48823 8384 49740 8412
rect 48823 8381 48835 8384
rect 48777 8375 48835 8381
rect 43073 8347 43131 8353
rect 41288 8316 41333 8344
rect 41288 8304 41294 8316
rect 43073 8313 43085 8347
rect 43119 8313 43131 8347
rect 43073 8307 43131 8313
rect 48685 8347 48743 8353
rect 48685 8313 48697 8347
rect 48731 8344 48743 8347
rect 49602 8344 49608 8356
rect 48731 8316 49608 8344
rect 48731 8313 48743 8316
rect 48685 8307 48743 8313
rect 49602 8304 49608 8316
rect 49660 8304 49666 8356
rect 49712 8353 49740 8384
rect 49697 8347 49755 8353
rect 49697 8313 49709 8347
rect 49743 8313 49755 8347
rect 49697 8307 49755 8313
rect 41248 8276 41276 8304
rect 48590 8276 48596 8288
rect 40328 8248 41276 8276
rect 48503 8248 48596 8276
rect 48590 8236 48596 8248
rect 48648 8276 48654 8288
rect 49326 8276 49332 8288
rect 48648 8248 49332 8276
rect 48648 8236 48654 8248
rect 49326 8236 49332 8248
rect 49384 8236 49390 8288
rect 49513 8279 49571 8285
rect 49513 8245 49525 8279
rect 49559 8276 49571 8279
rect 49970 8276 49976 8288
rect 49559 8248 49976 8276
rect 49559 8245 49571 8248
rect 49513 8239 49571 8245
rect 49970 8236 49976 8248
rect 50028 8236 50034 8288
rect 50341 8279 50399 8285
rect 50341 8245 50353 8279
rect 50387 8276 50399 8279
rect 50614 8276 50620 8288
rect 50387 8248 50620 8276
rect 50387 8245 50399 8248
rect 50341 8239 50399 8245
rect 50614 8236 50620 8248
rect 50672 8236 50678 8288
rect 1104 8186 68816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 65654 8186
rect 65706 8134 65718 8186
rect 65770 8134 65782 8186
rect 65834 8134 65846 8186
rect 65898 8134 65910 8186
rect 65962 8134 68816 8186
rect 1104 8112 68816 8134
rect 6457 8075 6515 8081
rect 6457 8041 6469 8075
rect 6503 8072 6515 8075
rect 6638 8072 6644 8084
rect 6503 8044 6644 8072
rect 6503 8041 6515 8044
rect 6457 8035 6515 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9582 8072 9588 8084
rect 8352 8044 9588 8072
rect 8352 8032 8358 8044
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 9861 8075 9919 8081
rect 9861 8041 9873 8075
rect 9907 8072 9919 8075
rect 9950 8072 9956 8084
rect 9907 8044 9956 8072
rect 9907 8041 9919 8044
rect 9861 8035 9919 8041
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10413 8075 10471 8081
rect 10413 8041 10425 8075
rect 10459 8072 10471 8075
rect 10459 8044 14780 8072
rect 10459 8041 10471 8044
rect 10413 8035 10471 8041
rect 4706 7896 4712 7948
rect 4764 7936 4770 7948
rect 5077 7939 5135 7945
rect 5077 7936 5089 7939
rect 4764 7908 5089 7936
rect 4764 7896 4770 7908
rect 5077 7905 5089 7908
rect 5123 7905 5135 7939
rect 5077 7899 5135 7905
rect 5350 7877 5356 7880
rect 5344 7868 5356 7877
rect 5311 7840 5356 7868
rect 5344 7831 5356 7840
rect 5350 7828 5356 7831
rect 5408 7828 5414 7880
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 9214 7868 9220 7880
rect 8067 7840 9220 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 10428 7868 10456 8035
rect 10962 8004 10968 8016
rect 10923 7976 10968 8004
rect 10962 7964 10968 7976
rect 11020 7964 11026 8016
rect 12345 8007 12403 8013
rect 12345 7973 12357 8007
rect 12391 8004 12403 8007
rect 13262 8004 13268 8016
rect 12391 7976 13268 8004
rect 12391 7973 12403 7976
rect 12345 7967 12403 7973
rect 13262 7964 13268 7976
rect 13320 7964 13326 8016
rect 14752 8004 14780 8044
rect 14826 8032 14832 8084
rect 14884 8072 14890 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 14884 8044 15117 8072
rect 14884 8032 14890 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 16393 8075 16451 8081
rect 16393 8041 16405 8075
rect 16439 8072 16451 8075
rect 16439 8044 16896 8072
rect 16439 8041 16451 8044
rect 16393 8035 16451 8041
rect 14752 7976 16344 8004
rect 12069 7939 12127 7945
rect 12069 7905 12081 7939
rect 12115 7936 12127 7939
rect 13722 7936 13728 7948
rect 12115 7908 13728 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 13722 7896 13728 7908
rect 13780 7896 13786 7948
rect 14642 7896 14648 7948
rect 14700 7936 14706 7948
rect 15749 7939 15807 7945
rect 15749 7936 15761 7939
rect 14700 7908 15761 7936
rect 14700 7896 14706 7908
rect 15749 7905 15761 7908
rect 15795 7905 15807 7939
rect 15749 7899 15807 7905
rect 9447 7840 10456 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 11422 7828 11428 7880
rect 11480 7868 11486 7880
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 11480 7840 11989 7868
rect 11480 7828 11486 7840
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 12618 7828 12624 7880
rect 12676 7868 12682 7880
rect 12805 7871 12863 7877
rect 12805 7868 12817 7871
rect 12676 7840 12817 7868
rect 12676 7828 12682 7840
rect 12805 7837 12817 7840
rect 12851 7837 12863 7871
rect 12805 7831 12863 7837
rect 12989 7871 13047 7877
rect 12989 7837 13001 7871
rect 13035 7868 13047 7871
rect 13541 7871 13599 7877
rect 13541 7868 13553 7871
rect 13035 7840 13553 7868
rect 13035 7837 13047 7840
rect 12989 7831 13047 7837
rect 13541 7837 13553 7840
rect 13587 7868 13599 7871
rect 14918 7868 14924 7880
rect 13587 7840 14924 7868
rect 13587 7837 13599 7840
rect 13541 7831 13599 7837
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 10870 7760 10876 7812
rect 10928 7800 10934 7812
rect 11149 7803 11207 7809
rect 11149 7800 11161 7803
rect 10928 7772 11161 7800
rect 10928 7760 10934 7772
rect 11149 7769 11161 7772
rect 11195 7769 11207 7803
rect 11149 7763 11207 7769
rect 11333 7803 11391 7809
rect 11333 7769 11345 7803
rect 11379 7800 11391 7803
rect 12897 7803 12955 7809
rect 12897 7800 12909 7803
rect 11379 7772 12909 7800
rect 11379 7769 11391 7772
rect 11333 7763 11391 7769
rect 12897 7769 12909 7772
rect 12943 7769 12955 7803
rect 14734 7800 14740 7812
rect 14695 7772 14740 7800
rect 12897 7763 12955 7769
rect 14734 7760 14740 7772
rect 14792 7760 14798 7812
rect 16316 7800 16344 7976
rect 16868 7877 16896 8044
rect 16942 8032 16948 8084
rect 17000 8072 17006 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 17000 8044 17049 8072
rect 17000 8032 17006 8044
rect 17037 8041 17049 8044
rect 17083 8041 17095 8075
rect 17037 8035 17095 8041
rect 19429 8075 19487 8081
rect 19429 8041 19441 8075
rect 19475 8072 19487 8075
rect 20162 8072 20168 8084
rect 19475 8044 20168 8072
rect 19475 8041 19487 8044
rect 19429 8035 19487 8041
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20806 8032 20812 8084
rect 20864 8072 20870 8084
rect 21269 8075 21327 8081
rect 21269 8072 21281 8075
rect 20864 8044 21281 8072
rect 20864 8032 20870 8044
rect 21269 8041 21281 8044
rect 21315 8072 21327 8075
rect 21818 8072 21824 8084
rect 21315 8044 21824 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 22646 8032 22652 8084
rect 22704 8072 22710 8084
rect 23201 8075 23259 8081
rect 23201 8072 23213 8075
rect 22704 8044 23213 8072
rect 22704 8032 22710 8044
rect 23201 8041 23213 8044
rect 23247 8041 23259 8075
rect 23201 8035 23259 8041
rect 24581 8075 24639 8081
rect 24581 8041 24593 8075
rect 24627 8072 24639 8075
rect 24670 8072 24676 8084
rect 24627 8044 24676 8072
rect 24627 8041 24639 8044
rect 24581 8035 24639 8041
rect 24670 8032 24676 8044
rect 24728 8032 24734 8084
rect 25314 8072 25320 8084
rect 25275 8044 25320 8072
rect 25314 8032 25320 8044
rect 25372 8032 25378 8084
rect 25774 8072 25780 8084
rect 25735 8044 25780 8072
rect 25774 8032 25780 8044
rect 25832 8032 25838 8084
rect 28258 8032 28264 8084
rect 28316 8072 28322 8084
rect 28445 8075 28503 8081
rect 28445 8072 28457 8075
rect 28316 8044 28457 8072
rect 28316 8032 28322 8044
rect 28445 8041 28457 8044
rect 28491 8072 28503 8075
rect 28626 8072 28632 8084
rect 28491 8044 28632 8072
rect 28491 8041 28503 8044
rect 28445 8035 28503 8041
rect 28626 8032 28632 8044
rect 28684 8032 28690 8084
rect 29638 8072 29644 8084
rect 29599 8044 29644 8072
rect 29638 8032 29644 8044
rect 29696 8032 29702 8084
rect 30558 8072 30564 8084
rect 30519 8044 30564 8072
rect 30558 8032 30564 8044
rect 30616 8032 30622 8084
rect 33781 8075 33839 8081
rect 33781 8072 33793 8075
rect 30760 8044 33793 8072
rect 20898 7964 20904 8016
rect 20956 8004 20962 8016
rect 21729 8007 21787 8013
rect 21729 8004 21741 8007
rect 20956 7976 21741 8004
rect 20956 7964 20962 7976
rect 21729 7973 21741 7976
rect 21775 7973 21787 8007
rect 25332 8004 25360 8032
rect 26234 8004 26240 8016
rect 25332 7976 26240 8004
rect 21729 7967 21787 7973
rect 26234 7964 26240 7976
rect 26292 7964 26298 8016
rect 26326 7964 26332 8016
rect 26384 8004 26390 8016
rect 26421 8007 26479 8013
rect 26421 8004 26433 8007
rect 26384 7976 26433 8004
rect 26384 7964 26390 7976
rect 26421 7973 26433 7976
rect 26467 7973 26479 8007
rect 26421 7967 26479 7973
rect 27801 8007 27859 8013
rect 27801 7973 27813 8007
rect 27847 8004 27859 8007
rect 30760 8004 30788 8044
rect 33781 8041 33793 8044
rect 33827 8041 33839 8075
rect 33781 8035 33839 8041
rect 33919 8075 33977 8081
rect 33919 8041 33931 8075
rect 33965 8072 33977 8075
rect 34238 8072 34244 8084
rect 33965 8044 34244 8072
rect 33965 8041 33977 8044
rect 33919 8035 33977 8041
rect 34238 8032 34244 8044
rect 34296 8072 34302 8084
rect 34790 8072 34796 8084
rect 34296 8044 34796 8072
rect 34296 8032 34302 8044
rect 34790 8032 34796 8044
rect 34848 8032 34854 8084
rect 35253 8075 35311 8081
rect 35253 8041 35265 8075
rect 35299 8072 35311 8075
rect 35342 8072 35348 8084
rect 35299 8044 35348 8072
rect 35299 8041 35311 8044
rect 35253 8035 35311 8041
rect 35342 8032 35348 8044
rect 35400 8032 35406 8084
rect 35710 8072 35716 8084
rect 35671 8044 35716 8072
rect 35710 8032 35716 8044
rect 35768 8032 35774 8084
rect 39301 8075 39359 8081
rect 39301 8041 39313 8075
rect 39347 8072 39359 8075
rect 40218 8072 40224 8084
rect 39347 8044 40224 8072
rect 39347 8041 39359 8044
rect 39301 8035 39359 8041
rect 40218 8032 40224 8044
rect 40276 8032 40282 8084
rect 40497 8075 40555 8081
rect 40497 8041 40509 8075
rect 40543 8041 40555 8075
rect 40497 8035 40555 8041
rect 27847 7976 30788 8004
rect 31205 8007 31263 8013
rect 27847 7973 27859 7976
rect 27801 7967 27859 7973
rect 31205 7973 31217 8007
rect 31251 8004 31263 8007
rect 31294 8004 31300 8016
rect 31251 7976 31300 8004
rect 31251 7973 31263 7976
rect 31205 7967 31263 7973
rect 31294 7964 31300 7976
rect 31352 7964 31358 8016
rect 40512 8004 40540 8035
rect 40954 8032 40960 8084
rect 41012 8072 41018 8084
rect 41417 8075 41475 8081
rect 41417 8072 41429 8075
rect 41012 8044 41429 8072
rect 41012 8032 41018 8044
rect 41417 8041 41429 8044
rect 41463 8041 41475 8075
rect 41690 8072 41696 8084
rect 41651 8044 41696 8072
rect 41417 8035 41475 8041
rect 41690 8032 41696 8044
rect 41748 8032 41754 8084
rect 49329 8075 49387 8081
rect 49329 8041 49341 8075
rect 49375 8072 49387 8075
rect 50154 8072 50160 8084
rect 49375 8044 50160 8072
rect 49375 8041 49387 8044
rect 49329 8035 49387 8041
rect 50154 8032 50160 8044
rect 50212 8032 50218 8084
rect 40862 8004 40868 8016
rect 39316 7976 40868 8004
rect 17862 7896 17868 7948
rect 17920 7936 17926 7948
rect 19150 7936 19156 7948
rect 17920 7908 19156 7936
rect 17920 7896 17926 7908
rect 19150 7896 19156 7908
rect 19208 7936 19214 7948
rect 19889 7939 19947 7945
rect 19889 7936 19901 7939
rect 19208 7908 19901 7936
rect 19208 7896 19214 7908
rect 19889 7905 19901 7908
rect 19935 7905 19947 7939
rect 22462 7936 22468 7948
rect 19889 7899 19947 7905
rect 20916 7908 22468 7936
rect 16853 7871 16911 7877
rect 16853 7837 16865 7871
rect 16899 7837 16911 7871
rect 18417 7871 18475 7877
rect 18417 7868 18429 7871
rect 16853 7831 16911 7837
rect 18064 7840 18429 7868
rect 18064 7800 18092 7840
rect 18417 7837 18429 7840
rect 18463 7837 18475 7871
rect 19242 7868 19248 7880
rect 19203 7840 19248 7868
rect 18417 7831 18475 7837
rect 18230 7800 18236 7812
rect 16316 7772 18092 7800
rect 18191 7772 18236 7800
rect 18230 7760 18236 7772
rect 18288 7760 18294 7812
rect 18432 7800 18460 7831
rect 19242 7828 19248 7840
rect 19300 7828 19306 7880
rect 19904 7868 19932 7899
rect 20916 7868 20944 7908
rect 22462 7896 22468 7908
rect 22520 7896 22526 7948
rect 27338 7936 27344 7948
rect 27299 7908 27344 7936
rect 27338 7896 27344 7908
rect 27396 7896 27402 7948
rect 32582 7936 32588 7948
rect 32543 7908 32588 7936
rect 32582 7896 32588 7908
rect 32640 7896 32646 7948
rect 34885 7939 34943 7945
rect 34885 7905 34897 7939
rect 34931 7936 34943 7939
rect 35434 7936 35440 7948
rect 34931 7908 35440 7936
rect 34931 7905 34943 7908
rect 34885 7899 34943 7905
rect 21910 7868 21916 7880
rect 19904 7840 20944 7868
rect 21871 7840 21916 7868
rect 21910 7828 21916 7840
rect 21968 7828 21974 7880
rect 22005 7871 22063 7877
rect 22005 7837 22017 7871
rect 22051 7868 22063 7871
rect 22186 7868 22192 7880
rect 22051 7840 22192 7868
rect 22051 7837 22063 7840
rect 22005 7831 22063 7837
rect 22186 7828 22192 7840
rect 22244 7828 22250 7880
rect 22281 7871 22339 7877
rect 22281 7837 22293 7871
rect 22327 7837 22339 7871
rect 23382 7868 23388 7880
rect 23343 7840 23388 7868
rect 22281 7831 22339 7837
rect 19426 7800 19432 7812
rect 18432 7772 19432 7800
rect 19426 7760 19432 7772
rect 19484 7760 19490 7812
rect 20162 7809 20168 7812
rect 20156 7800 20168 7809
rect 20123 7772 20168 7800
rect 20156 7763 20168 7772
rect 20162 7760 20168 7763
rect 20220 7760 20226 7812
rect 20438 7760 20444 7812
rect 20496 7800 20502 7812
rect 21928 7800 21956 7828
rect 22094 7800 22100 7812
rect 20496 7772 21956 7800
rect 22055 7772 22100 7800
rect 20496 7760 20502 7772
rect 22094 7760 22100 7772
rect 22152 7760 22158 7812
rect 7834 7732 7840 7744
rect 7795 7704 7840 7732
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 14277 7735 14335 7741
rect 14277 7701 14289 7735
rect 14323 7732 14335 7735
rect 15930 7732 15936 7744
rect 14323 7704 15936 7732
rect 14323 7701 14335 7704
rect 14277 7695 14335 7701
rect 15930 7692 15936 7704
rect 15988 7692 15994 7744
rect 16025 7735 16083 7741
rect 16025 7701 16037 7735
rect 16071 7732 16083 7735
rect 18046 7732 18052 7744
rect 16071 7704 18052 7732
rect 16071 7701 16083 7704
rect 16025 7695 16083 7701
rect 18046 7692 18052 7704
rect 18104 7692 18110 7744
rect 21818 7692 21824 7744
rect 21876 7732 21882 7744
rect 22296 7732 22324 7831
rect 23382 7828 23388 7840
rect 23440 7828 23446 7880
rect 23474 7828 23480 7880
rect 23532 7868 23538 7880
rect 24394 7868 24400 7880
rect 23532 7840 23577 7868
rect 24355 7840 24400 7868
rect 23532 7828 23538 7840
rect 24394 7828 24400 7840
rect 24452 7828 24458 7880
rect 27430 7868 27436 7880
rect 27391 7840 27436 7868
rect 27430 7828 27436 7840
rect 27488 7828 27494 7880
rect 30374 7868 30380 7880
rect 28184 7840 30236 7868
rect 30335 7840 30380 7868
rect 25774 7760 25780 7812
rect 25832 7800 25838 7812
rect 26789 7803 26847 7809
rect 26789 7800 26801 7803
rect 25832 7772 26801 7800
rect 25832 7760 25838 7772
rect 26789 7769 26801 7772
rect 26835 7800 26847 7803
rect 28184 7800 28212 7840
rect 28350 7800 28356 7812
rect 26835 7772 28212 7800
rect 28311 7772 28356 7800
rect 26835 7769 26847 7772
rect 26789 7763 26847 7769
rect 28350 7760 28356 7772
rect 28408 7760 28414 7812
rect 30208 7800 30236 7840
rect 30374 7828 30380 7840
rect 30432 7828 30438 7880
rect 32329 7871 32387 7877
rect 32329 7837 32341 7871
rect 32375 7868 32387 7871
rect 32950 7868 32956 7880
rect 32375 7840 32956 7868
rect 32375 7837 32387 7840
rect 32329 7831 32387 7837
rect 32950 7828 32956 7840
rect 33008 7828 33014 7880
rect 33594 7868 33600 7880
rect 33555 7840 33600 7868
rect 33594 7828 33600 7840
rect 33652 7828 33658 7880
rect 34057 7871 34115 7877
rect 34057 7837 34069 7871
rect 34103 7868 34115 7871
rect 34900 7868 34928 7899
rect 35434 7896 35440 7908
rect 35492 7896 35498 7948
rect 34103 7840 34928 7868
rect 35069 7871 35127 7877
rect 34103 7837 34115 7840
rect 34057 7831 34115 7837
rect 35069 7837 35081 7871
rect 35115 7837 35127 7871
rect 35069 7831 35127 7837
rect 30208 7772 31754 7800
rect 21876 7704 22324 7732
rect 26329 7735 26387 7741
rect 21876 7692 21882 7704
rect 26329 7701 26341 7735
rect 26375 7732 26387 7735
rect 26418 7732 26424 7744
rect 26375 7704 26424 7732
rect 26375 7701 26387 7704
rect 26329 7695 26387 7701
rect 26418 7692 26424 7704
rect 26476 7692 26482 7744
rect 31726 7732 31754 7772
rect 34790 7760 34796 7812
rect 34848 7800 34854 7812
rect 35084 7800 35112 7831
rect 35526 7828 35532 7880
rect 35584 7868 35590 7880
rect 35897 7871 35955 7877
rect 35897 7868 35909 7871
rect 35584 7840 35909 7868
rect 35584 7828 35590 7840
rect 35897 7837 35909 7840
rect 35943 7837 35955 7871
rect 35897 7831 35955 7837
rect 39025 7871 39083 7877
rect 39025 7837 39037 7871
rect 39071 7837 39083 7871
rect 39025 7831 39083 7837
rect 34848 7772 35112 7800
rect 39040 7800 39068 7831
rect 39206 7828 39212 7880
rect 39264 7868 39270 7880
rect 39316 7877 39344 7976
rect 40862 7964 40868 7976
rect 40920 7964 40926 8016
rect 46934 7964 46940 8016
rect 46992 8004 46998 8016
rect 54662 8004 54668 8016
rect 46992 7976 54668 8004
rect 46992 7964 46998 7976
rect 54662 7964 54668 7976
rect 54720 7964 54726 8016
rect 41138 7896 41144 7948
rect 41196 7936 41202 7948
rect 49421 7939 49479 7945
rect 41196 7908 43944 7936
rect 41196 7896 41202 7908
rect 39301 7871 39359 7877
rect 39301 7868 39313 7871
rect 39264 7840 39313 7868
rect 39264 7828 39270 7840
rect 39301 7837 39313 7840
rect 39347 7837 39359 7871
rect 41598 7868 41604 7880
rect 39301 7831 39359 7837
rect 40236 7840 40540 7868
rect 41559 7840 41604 7868
rect 40034 7800 40040 7812
rect 39040 7772 40040 7800
rect 34848 7760 34854 7772
rect 40034 7760 40040 7772
rect 40092 7800 40098 7812
rect 40236 7800 40264 7840
rect 40092 7772 40264 7800
rect 40313 7803 40371 7809
rect 40092 7760 40098 7772
rect 40313 7769 40325 7803
rect 40359 7800 40371 7803
rect 40402 7800 40408 7812
rect 40359 7772 40408 7800
rect 40359 7769 40371 7772
rect 40313 7763 40371 7769
rect 32398 7732 32404 7744
rect 31726 7704 32404 7732
rect 32398 7692 32404 7704
rect 32456 7732 32462 7744
rect 33045 7735 33103 7741
rect 33045 7732 33057 7735
rect 32456 7704 33057 7732
rect 32456 7692 32462 7704
rect 33045 7701 33057 7704
rect 33091 7701 33103 7735
rect 33045 7695 33103 7701
rect 33689 7735 33747 7741
rect 33689 7701 33701 7735
rect 33735 7732 33747 7735
rect 34422 7732 34428 7744
rect 33735 7704 34428 7732
rect 33735 7701 33747 7704
rect 33689 7695 33747 7701
rect 34422 7692 34428 7704
rect 34480 7692 34486 7744
rect 39117 7735 39175 7741
rect 39117 7701 39129 7735
rect 39163 7732 39175 7735
rect 40328 7732 40356 7763
rect 40402 7760 40408 7772
rect 40460 7760 40466 7812
rect 40512 7809 40540 7840
rect 41598 7828 41604 7840
rect 41656 7828 41662 7880
rect 41693 7871 41751 7877
rect 41693 7837 41705 7871
rect 41739 7837 41751 7871
rect 41693 7831 41751 7837
rect 42061 7871 42119 7877
rect 42061 7837 42073 7871
rect 42107 7868 42119 7871
rect 43254 7868 43260 7880
rect 42107 7840 43260 7868
rect 42107 7837 42119 7840
rect 42061 7831 42119 7837
rect 40512 7803 40571 7809
rect 40512 7772 40525 7803
rect 40513 7769 40525 7772
rect 40559 7800 40571 7803
rect 41708 7800 41736 7831
rect 43254 7828 43260 7840
rect 43312 7828 43318 7880
rect 43916 7877 43944 7908
rect 49421 7905 49433 7939
rect 49467 7936 49479 7939
rect 49694 7936 49700 7948
rect 49467 7908 49700 7936
rect 49467 7905 49479 7908
rect 49421 7899 49479 7905
rect 49694 7896 49700 7908
rect 49752 7896 49758 7948
rect 43901 7871 43959 7877
rect 43901 7837 43913 7871
rect 43947 7837 43959 7871
rect 44177 7871 44235 7877
rect 44177 7868 44189 7871
rect 43901 7831 43959 7837
rect 44008 7840 44189 7868
rect 40559 7772 41736 7800
rect 40559 7769 40571 7772
rect 40513 7763 40571 7769
rect 43070 7760 43076 7812
rect 43128 7800 43134 7812
rect 44008 7800 44036 7840
rect 44177 7837 44189 7840
rect 44223 7868 44235 7871
rect 45002 7868 45008 7880
rect 44223 7840 45008 7868
rect 44223 7837 44235 7840
rect 44177 7831 44235 7837
rect 45002 7828 45008 7840
rect 45060 7828 45066 7880
rect 45189 7871 45247 7877
rect 45189 7837 45201 7871
rect 45235 7868 45247 7871
rect 45554 7868 45560 7880
rect 45235 7840 45560 7868
rect 45235 7837 45247 7840
rect 45189 7831 45247 7837
rect 45554 7828 45560 7840
rect 45612 7828 45618 7880
rect 48314 7868 48320 7880
rect 48275 7840 48320 7868
rect 48314 7828 48320 7840
rect 48372 7828 48378 7880
rect 48501 7871 48559 7877
rect 48501 7837 48513 7871
rect 48547 7868 48559 7871
rect 48590 7868 48596 7880
rect 48547 7840 48596 7868
rect 48547 7837 48559 7840
rect 48501 7831 48559 7837
rect 48590 7828 48596 7840
rect 48648 7828 48654 7880
rect 49145 7871 49203 7877
rect 49145 7837 49157 7871
rect 49191 7868 49203 7871
rect 49326 7868 49332 7880
rect 49191 7840 49332 7868
rect 49191 7837 49203 7840
rect 49145 7831 49203 7837
rect 49326 7828 49332 7840
rect 49384 7828 49390 7880
rect 50341 7871 50399 7877
rect 50341 7837 50353 7871
rect 50387 7868 50399 7871
rect 50706 7868 50712 7880
rect 50387 7840 50712 7868
rect 50387 7837 50399 7840
rect 50341 7831 50399 7837
rect 50706 7828 50712 7840
rect 50764 7828 50770 7880
rect 43128 7772 44036 7800
rect 48409 7803 48467 7809
rect 43128 7760 43134 7772
rect 48409 7769 48421 7803
rect 48455 7800 48467 7803
rect 49970 7800 49976 7812
rect 48455 7772 49976 7800
rect 48455 7769 48467 7772
rect 48409 7763 48467 7769
rect 49970 7760 49976 7772
rect 50028 7760 50034 7812
rect 39163 7704 40356 7732
rect 40681 7735 40739 7741
rect 39163 7701 39175 7704
rect 39117 7695 39175 7701
rect 40681 7701 40693 7735
rect 40727 7732 40739 7735
rect 41230 7732 41236 7744
rect 40727 7704 41236 7732
rect 40727 7701 40739 7704
rect 40681 7695 40739 7701
rect 41230 7692 41236 7704
rect 41288 7692 41294 7744
rect 43717 7735 43775 7741
rect 43717 7701 43729 7735
rect 43763 7732 43775 7735
rect 43990 7732 43996 7744
rect 43763 7704 43996 7732
rect 43763 7701 43775 7704
rect 43717 7695 43775 7701
rect 43990 7692 43996 7704
rect 44048 7692 44054 7744
rect 44082 7692 44088 7744
rect 44140 7732 44146 7744
rect 45094 7732 45100 7744
rect 44140 7704 44185 7732
rect 45055 7704 45100 7732
rect 44140 7692 44146 7704
rect 45094 7692 45100 7704
rect 45152 7692 45158 7744
rect 48590 7692 48596 7744
rect 48648 7732 48654 7744
rect 48961 7735 49019 7741
rect 48961 7732 48973 7735
rect 48648 7704 48973 7732
rect 48648 7692 48654 7704
rect 48961 7701 48973 7704
rect 49007 7701 49019 7735
rect 48961 7695 49019 7701
rect 49694 7692 49700 7744
rect 49752 7732 49758 7744
rect 50157 7735 50215 7741
rect 50157 7732 50169 7735
rect 49752 7704 50169 7732
rect 49752 7692 49758 7704
rect 50157 7701 50169 7704
rect 50203 7701 50215 7735
rect 50157 7695 50215 7701
rect 1104 7642 68816 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 68816 7642
rect 1104 7568 68816 7590
rect 8757 7531 8815 7537
rect 8757 7497 8769 7531
rect 8803 7497 8815 7531
rect 9214 7528 9220 7540
rect 9175 7500 9220 7528
rect 8757 7491 8815 7497
rect 7644 7463 7702 7469
rect 7644 7429 7656 7463
rect 7690 7460 7702 7463
rect 7834 7460 7840 7472
rect 7690 7432 7840 7460
rect 7690 7429 7702 7432
rect 7644 7423 7702 7429
rect 7834 7420 7840 7432
rect 7892 7420 7898 7472
rect 8772 7460 8800 7491
rect 9214 7488 9220 7500
rect 9272 7488 9278 7540
rect 9306 7488 9312 7540
rect 9364 7528 9370 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 9364 7500 9597 7528
rect 9364 7488 9370 7500
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 9585 7491 9643 7497
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 10928 7500 11529 7528
rect 10928 7488 10934 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 20346 7488 20352 7540
rect 20404 7528 20410 7540
rect 20625 7531 20683 7537
rect 20625 7528 20637 7531
rect 20404 7500 20637 7528
rect 20404 7488 20410 7500
rect 20625 7497 20637 7500
rect 20671 7497 20683 7531
rect 21174 7528 21180 7540
rect 21087 7500 21180 7528
rect 20625 7491 20683 7497
rect 21174 7488 21180 7500
rect 21232 7528 21238 7540
rect 21818 7528 21824 7540
rect 21232 7500 21824 7528
rect 21232 7488 21238 7500
rect 21818 7488 21824 7500
rect 21876 7488 21882 7540
rect 28258 7528 28264 7540
rect 21928 7500 26234 7528
rect 28219 7500 28264 7528
rect 9324 7460 9352 7488
rect 8772 7432 9352 7460
rect 10965 7463 11023 7469
rect 10965 7429 10977 7463
rect 11011 7460 11023 7463
rect 11974 7460 11980 7472
rect 11011 7432 11980 7460
rect 11011 7429 11023 7432
rect 10965 7423 11023 7429
rect 11974 7420 11980 7432
rect 12032 7420 12038 7472
rect 14277 7463 14335 7469
rect 14277 7429 14289 7463
rect 14323 7460 14335 7463
rect 14734 7460 14740 7472
rect 14323 7432 14740 7460
rect 14323 7429 14335 7432
rect 14277 7423 14335 7429
rect 14734 7420 14740 7432
rect 14792 7420 14798 7472
rect 18230 7420 18236 7472
rect 18288 7460 18294 7472
rect 18601 7463 18659 7469
rect 18601 7460 18613 7463
rect 18288 7432 18613 7460
rect 18288 7420 18294 7432
rect 18601 7429 18613 7432
rect 18647 7460 18659 7463
rect 21928 7460 21956 7500
rect 18647 7432 21956 7460
rect 22097 7463 22155 7469
rect 18647 7429 18659 7432
rect 18601 7423 18659 7429
rect 22097 7429 22109 7463
rect 22143 7460 22155 7463
rect 22186 7460 22192 7472
rect 22143 7432 22192 7460
rect 22143 7429 22155 7432
rect 22097 7423 22155 7429
rect 22186 7420 22192 7432
rect 22244 7420 22250 7472
rect 22278 7420 22284 7472
rect 22336 7460 22342 7472
rect 23014 7460 23020 7472
rect 22336 7432 22381 7460
rect 22975 7432 23020 7460
rect 22336 7420 22342 7432
rect 23014 7420 23020 7432
rect 23072 7420 23078 7472
rect 25317 7463 25375 7469
rect 25317 7460 25329 7463
rect 24242 7432 25329 7460
rect 25317 7429 25329 7432
rect 25363 7429 25375 7463
rect 26206 7460 26234 7500
rect 28258 7488 28264 7500
rect 28316 7488 28322 7540
rect 28350 7488 28356 7540
rect 28408 7528 28414 7540
rect 28810 7528 28816 7540
rect 28408 7500 28816 7528
rect 28408 7488 28414 7500
rect 28810 7488 28816 7500
rect 28868 7488 28874 7540
rect 31202 7488 31208 7540
rect 31260 7528 31266 7540
rect 31389 7531 31447 7537
rect 31389 7528 31401 7531
rect 31260 7500 31401 7528
rect 31260 7488 31266 7500
rect 31389 7497 31401 7500
rect 31435 7497 31447 7531
rect 35526 7528 35532 7540
rect 35487 7500 35532 7528
rect 31389 7491 31447 7497
rect 35526 7488 35532 7500
rect 35584 7488 35590 7540
rect 41049 7531 41107 7537
rect 41049 7497 41061 7531
rect 41095 7528 41107 7531
rect 41138 7528 41144 7540
rect 41095 7500 41144 7528
rect 41095 7497 41107 7500
rect 41049 7491 41107 7497
rect 41138 7488 41144 7500
rect 41196 7488 41202 7540
rect 41598 7488 41604 7540
rect 41656 7488 41662 7540
rect 41782 7528 41788 7540
rect 41743 7500 41788 7528
rect 41782 7488 41788 7500
rect 41840 7488 41846 7540
rect 44082 7488 44088 7540
rect 44140 7528 44146 7540
rect 45465 7531 45523 7537
rect 45465 7528 45477 7531
rect 44140 7500 45477 7528
rect 44140 7488 44146 7500
rect 45465 7497 45477 7500
rect 45511 7528 45523 7531
rect 52730 7528 52736 7540
rect 45511 7500 52736 7528
rect 45511 7497 45523 7500
rect 45465 7491 45523 7497
rect 52730 7488 52736 7500
rect 52788 7488 52794 7540
rect 27341 7463 27399 7469
rect 27341 7460 27353 7463
rect 26206 7432 27353 7460
rect 25317 7423 25375 7429
rect 27341 7429 27353 7432
rect 27387 7460 27399 7463
rect 29178 7460 29184 7472
rect 27387 7432 29184 7460
rect 27387 7429 27399 7432
rect 27341 7423 27399 7429
rect 29178 7420 29184 7432
rect 29236 7420 29242 7472
rect 29546 7420 29552 7472
rect 29604 7460 29610 7472
rect 29604 7432 37320 7460
rect 29604 7420 29610 7432
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7392 6607 7395
rect 7190 7392 7196 7404
rect 6595 7364 7196 7392
rect 6595 7361 6607 7364
rect 6549 7355 6607 7361
rect 7190 7352 7196 7364
rect 7248 7352 7254 7404
rect 7926 7352 7932 7404
rect 7984 7392 7990 7404
rect 15470 7392 15476 7404
rect 7984 7364 9812 7392
rect 15431 7364 15476 7392
rect 7984 7352 7990 7364
rect 5350 7284 5356 7336
rect 5408 7324 5414 7336
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 5408 7296 7389 7324
rect 5408 7284 5414 7296
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 7377 7287 7435 7293
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 9784 7333 9812 7364
rect 15470 7352 15476 7364
rect 15528 7352 15534 7404
rect 19150 7352 19156 7404
rect 19208 7392 19214 7404
rect 19245 7395 19303 7401
rect 19245 7392 19257 7395
rect 19208 7364 19257 7392
rect 19208 7352 19214 7364
rect 19245 7361 19257 7364
rect 19291 7361 19303 7395
rect 19245 7355 19303 7361
rect 19334 7352 19340 7404
rect 19392 7392 19398 7404
rect 19501 7395 19559 7401
rect 19501 7392 19513 7395
rect 19392 7364 19513 7392
rect 19392 7352 19398 7364
rect 19501 7361 19513 7364
rect 19547 7361 19559 7395
rect 19501 7355 19559 7361
rect 19794 7352 19800 7404
rect 19852 7392 19858 7404
rect 20990 7392 20996 7404
rect 19852 7364 20996 7392
rect 19852 7352 19858 7364
rect 20990 7352 20996 7364
rect 21048 7392 21054 7404
rect 21085 7395 21143 7401
rect 21085 7392 21097 7395
rect 21048 7364 21097 7392
rect 21048 7352 21054 7364
rect 21085 7361 21097 7364
rect 21131 7361 21143 7395
rect 21085 7355 21143 7361
rect 24670 7352 24676 7404
rect 24728 7392 24734 7404
rect 25222 7392 25228 7404
rect 24728 7364 25228 7392
rect 24728 7352 24734 7364
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 26421 7395 26479 7401
rect 26421 7361 26433 7395
rect 26467 7392 26479 7395
rect 27706 7392 27712 7404
rect 26467 7364 27712 7392
rect 26467 7361 26479 7364
rect 26421 7355 26479 7361
rect 27706 7352 27712 7364
rect 27764 7352 27770 7404
rect 30650 7352 30656 7404
rect 30708 7392 30714 7404
rect 30745 7395 30803 7401
rect 30745 7392 30757 7395
rect 30708 7364 30757 7392
rect 30708 7352 30714 7364
rect 30745 7361 30757 7364
rect 30791 7392 30803 7395
rect 31297 7395 31355 7401
rect 31297 7392 31309 7395
rect 30791 7364 31309 7392
rect 30791 7361 30803 7364
rect 30745 7355 30803 7361
rect 31297 7361 31309 7364
rect 31343 7361 31355 7395
rect 32398 7392 32404 7404
rect 32359 7364 32404 7392
rect 31297 7355 31355 7361
rect 32398 7352 32404 7364
rect 32456 7352 32462 7404
rect 34422 7392 34428 7404
rect 34383 7364 34428 7392
rect 34422 7352 34428 7364
rect 34480 7352 34486 7404
rect 34698 7392 34704 7404
rect 34659 7364 34704 7392
rect 34698 7352 34704 7364
rect 34756 7352 34762 7404
rect 35342 7392 35348 7404
rect 35303 7364 35348 7392
rect 35342 7352 35348 7364
rect 35400 7352 35406 7404
rect 37292 7401 37320 7432
rect 39574 7420 39580 7472
rect 39632 7420 39638 7472
rect 40310 7420 40316 7472
rect 40368 7460 40374 7472
rect 41616 7460 41644 7488
rect 43990 7460 43996 7472
rect 40368 7432 40540 7460
rect 41616 7432 43024 7460
rect 43951 7432 43996 7460
rect 40368 7420 40374 7432
rect 37277 7395 37335 7401
rect 37277 7361 37289 7395
rect 37323 7392 37335 7395
rect 38010 7392 38016 7404
rect 37323 7364 38016 7392
rect 37323 7361 37335 7364
rect 37277 7355 37335 7361
rect 38010 7352 38016 7364
rect 38068 7352 38074 7404
rect 40512 7401 40540 7432
rect 40497 7395 40555 7401
rect 40497 7361 40509 7395
rect 40543 7361 40555 7395
rect 40497 7355 40555 7361
rect 40862 7352 40868 7404
rect 40920 7392 40926 7404
rect 40957 7395 41015 7401
rect 40957 7392 40969 7395
rect 40920 7364 40969 7392
rect 40920 7352 40926 7364
rect 40957 7361 40969 7364
rect 41003 7361 41015 7395
rect 40957 7355 41015 7361
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 9364 7296 9689 7324
rect 9364 7284 9370 7296
rect 9677 7293 9689 7296
rect 9723 7293 9735 7327
rect 9677 7287 9735 7293
rect 9769 7327 9827 7333
rect 9769 7293 9781 7327
rect 9815 7293 9827 7327
rect 13449 7327 13507 7333
rect 13449 7324 13461 7327
rect 9769 7287 9827 7293
rect 12820 7296 13461 7324
rect 10502 7216 10508 7268
rect 10560 7256 10566 7268
rect 11701 7259 11759 7265
rect 11701 7256 11713 7259
rect 10560 7228 11713 7256
rect 10560 7216 10566 7228
rect 11701 7225 11713 7228
rect 11747 7256 11759 7259
rect 12618 7256 12624 7268
rect 11747 7228 12624 7256
rect 11747 7225 11759 7228
rect 11701 7219 11759 7225
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 6362 7188 6368 7200
rect 6323 7160 6368 7188
rect 6362 7148 6368 7160
rect 6420 7148 6426 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12820 7188 12848 7296
rect 13449 7293 13461 7296
rect 13495 7324 13507 7327
rect 14369 7327 14427 7333
rect 14369 7324 14381 7327
rect 13495 7296 14381 7324
rect 13495 7293 13507 7296
rect 13449 7287 13507 7293
rect 14369 7293 14381 7296
rect 14415 7324 14427 7327
rect 14458 7324 14464 7336
rect 14415 7296 14464 7324
rect 14415 7293 14427 7296
rect 14369 7287 14427 7293
rect 14458 7284 14464 7296
rect 14516 7284 14522 7336
rect 14553 7327 14611 7333
rect 14553 7293 14565 7327
rect 14599 7324 14611 7327
rect 14642 7324 14648 7336
rect 14599 7296 14648 7324
rect 14599 7293 14611 7296
rect 14553 7287 14611 7293
rect 14642 7284 14648 7296
rect 14700 7324 14706 7336
rect 15197 7327 15255 7333
rect 15197 7324 15209 7327
rect 14700 7296 15209 7324
rect 14700 7284 14706 7296
rect 15197 7293 15209 7296
rect 15243 7293 15255 7327
rect 15378 7324 15384 7336
rect 15339 7296 15384 7324
rect 15197 7287 15255 7293
rect 15378 7284 15384 7296
rect 15436 7324 15442 7336
rect 16666 7324 16672 7336
rect 15436 7296 16672 7324
rect 15436 7284 15442 7296
rect 16666 7284 16672 7296
rect 16724 7284 16730 7336
rect 20254 7284 20260 7336
rect 20312 7324 20318 7336
rect 22094 7324 22100 7336
rect 20312 7296 22100 7324
rect 20312 7284 20318 7296
rect 22094 7284 22100 7296
rect 22152 7284 22158 7336
rect 22462 7284 22468 7336
rect 22520 7324 22526 7336
rect 22741 7327 22799 7333
rect 22741 7324 22753 7327
rect 22520 7296 22753 7324
rect 22520 7284 22526 7296
rect 22741 7293 22753 7296
rect 22787 7293 22799 7327
rect 24762 7324 24768 7336
rect 24675 7296 24768 7324
rect 22741 7287 22799 7293
rect 24762 7284 24768 7296
rect 24820 7324 24826 7336
rect 28626 7324 28632 7336
rect 24820 7296 28632 7324
rect 24820 7284 24826 7296
rect 28626 7284 28632 7296
rect 28684 7284 28690 7336
rect 32122 7324 32128 7336
rect 32083 7296 32128 7324
rect 32122 7284 32128 7296
rect 32180 7284 32186 7336
rect 35161 7327 35219 7333
rect 35161 7293 35173 7327
rect 35207 7324 35219 7327
rect 35434 7324 35440 7336
rect 35207 7296 35440 7324
rect 35207 7293 35219 7296
rect 35161 7287 35219 7293
rect 35434 7284 35440 7296
rect 35492 7284 35498 7336
rect 40218 7324 40224 7336
rect 40179 7296 40224 7324
rect 40218 7284 40224 7296
rect 40276 7284 40282 7336
rect 12897 7259 12955 7265
rect 12897 7225 12909 7259
rect 12943 7256 12955 7259
rect 14090 7256 14096 7268
rect 12943 7228 14096 7256
rect 12943 7225 12955 7228
rect 12897 7219 12955 7225
rect 14090 7216 14096 7228
rect 14148 7216 14154 7268
rect 15841 7259 15899 7265
rect 15841 7225 15853 7259
rect 15887 7256 15899 7259
rect 16758 7256 16764 7268
rect 15887 7228 16764 7256
rect 15887 7225 15899 7228
rect 15841 7219 15899 7225
rect 16758 7216 16764 7228
rect 16816 7216 16822 7268
rect 26234 7216 26240 7268
rect 26292 7256 26298 7268
rect 40972 7256 41000 7355
rect 41046 7352 41052 7404
rect 41104 7392 41110 7404
rect 41141 7395 41199 7401
rect 41141 7392 41153 7395
rect 41104 7364 41153 7392
rect 41104 7352 41110 7364
rect 41141 7361 41153 7364
rect 41187 7361 41199 7395
rect 41141 7355 41199 7361
rect 41230 7352 41236 7404
rect 41288 7392 41294 7404
rect 41601 7395 41659 7401
rect 41601 7392 41613 7395
rect 41288 7364 41613 7392
rect 41288 7352 41294 7364
rect 41601 7361 41613 7364
rect 41647 7361 41659 7395
rect 41782 7392 41788 7404
rect 41743 7364 41788 7392
rect 41601 7355 41659 7361
rect 41782 7352 41788 7364
rect 41840 7352 41846 7404
rect 42996 7392 43024 7432
rect 43990 7420 43996 7432
rect 44048 7420 44054 7472
rect 43070 7392 43076 7404
rect 42983 7364 43076 7392
rect 42996 7362 43076 7364
rect 43070 7352 43076 7362
rect 43128 7352 43134 7404
rect 43254 7392 43260 7404
rect 43215 7364 43260 7392
rect 43254 7352 43260 7364
rect 43312 7352 43318 7404
rect 45094 7352 45100 7404
rect 45152 7352 45158 7404
rect 48498 7392 48504 7404
rect 48459 7364 48504 7392
rect 48498 7352 48504 7364
rect 48556 7352 48562 7404
rect 49697 7395 49755 7401
rect 49697 7361 49709 7395
rect 49743 7392 49755 7395
rect 49786 7392 49792 7404
rect 49743 7364 49792 7392
rect 49743 7361 49755 7364
rect 49697 7355 49755 7361
rect 49786 7352 49792 7364
rect 49844 7352 49850 7404
rect 49970 7392 49976 7404
rect 49931 7364 49976 7392
rect 49970 7352 49976 7364
rect 50028 7352 50034 7404
rect 43714 7324 43720 7336
rect 43675 7296 43720 7324
rect 43714 7284 43720 7296
rect 43772 7284 43778 7336
rect 41230 7256 41236 7268
rect 26292 7228 26337 7256
rect 40972 7228 41236 7256
rect 26292 7216 26298 7228
rect 41230 7216 41236 7228
rect 41288 7216 41294 7268
rect 48961 7259 49019 7265
rect 48961 7256 48973 7259
rect 45020 7228 48973 7256
rect 13906 7188 13912 7200
rect 12032 7160 12848 7188
rect 13867 7160 13912 7188
rect 12032 7148 12038 7160
rect 13906 7148 13912 7160
rect 13964 7148 13970 7200
rect 33318 7148 33324 7200
rect 33376 7188 33382 7200
rect 33689 7191 33747 7197
rect 33689 7188 33701 7191
rect 33376 7160 33701 7188
rect 33376 7148 33382 7160
rect 33689 7157 33701 7160
rect 33735 7157 33747 7191
rect 37458 7188 37464 7200
rect 37419 7160 37464 7188
rect 33689 7151 33747 7157
rect 37458 7148 37464 7160
rect 37516 7148 37522 7200
rect 38749 7191 38807 7197
rect 38749 7157 38761 7191
rect 38795 7188 38807 7191
rect 40126 7188 40132 7200
rect 38795 7160 40132 7188
rect 38795 7157 38807 7160
rect 38749 7151 38807 7157
rect 40126 7148 40132 7160
rect 40184 7148 40190 7200
rect 43257 7191 43315 7197
rect 43257 7157 43269 7191
rect 43303 7188 43315 7191
rect 43990 7188 43996 7200
rect 43303 7160 43996 7188
rect 43303 7157 43315 7160
rect 43257 7151 43315 7157
rect 43990 7148 43996 7160
rect 44048 7148 44054 7200
rect 44450 7148 44456 7200
rect 44508 7188 44514 7200
rect 45020 7188 45048 7228
rect 48961 7225 48973 7228
rect 49007 7225 49019 7259
rect 48961 7219 49019 7225
rect 47854 7188 47860 7200
rect 44508 7160 45048 7188
rect 47815 7160 47860 7188
rect 44508 7148 44514 7160
rect 47854 7148 47860 7160
rect 47912 7148 47918 7200
rect 48314 7188 48320 7200
rect 48275 7160 48320 7188
rect 48314 7148 48320 7160
rect 48372 7148 48378 7200
rect 1104 7098 68816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 65654 7098
rect 65706 7046 65718 7098
rect 65770 7046 65782 7098
rect 65834 7046 65846 7098
rect 65898 7046 65910 7098
rect 65962 7046 68816 7098
rect 1104 7024 68816 7046
rect 7190 6984 7196 6996
rect 7151 6956 7196 6984
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 22097 6987 22155 6993
rect 22097 6953 22109 6987
rect 22143 6984 22155 6987
rect 22186 6984 22192 6996
rect 22143 6956 22192 6984
rect 22143 6953 22155 6956
rect 22097 6947 22155 6953
rect 22186 6944 22192 6956
rect 22244 6944 22250 6996
rect 22296 6956 23796 6984
rect 16666 6876 16672 6928
rect 16724 6916 16730 6928
rect 22296 6916 22324 6956
rect 16724 6888 22324 6916
rect 23569 6919 23627 6925
rect 16724 6876 16730 6888
rect 23569 6885 23581 6919
rect 23615 6914 23627 6919
rect 23768 6916 23796 6956
rect 23842 6944 23848 6996
rect 23900 6984 23906 6996
rect 24581 6987 24639 6993
rect 24581 6984 24593 6987
rect 23900 6956 24593 6984
rect 23900 6944 23906 6956
rect 24581 6953 24593 6956
rect 24627 6984 24639 6987
rect 26418 6984 26424 6996
rect 24627 6956 26424 6984
rect 24627 6953 24639 6956
rect 24581 6947 24639 6953
rect 26418 6944 26424 6956
rect 26476 6984 26482 6996
rect 27154 6984 27160 6996
rect 26476 6956 27160 6984
rect 26476 6944 26482 6956
rect 27154 6944 27160 6956
rect 27212 6944 27218 6996
rect 27246 6944 27252 6996
rect 27304 6984 27310 6996
rect 27430 6984 27436 6996
rect 27304 6956 27436 6984
rect 27304 6944 27310 6956
rect 27430 6944 27436 6956
rect 27488 6944 27494 6996
rect 34790 6984 34796 6996
rect 34751 6956 34796 6984
rect 34790 6944 34796 6956
rect 34848 6944 34854 6996
rect 37458 6944 37464 6996
rect 37516 6984 37522 6996
rect 37516 6956 40172 6984
rect 37516 6944 37522 6956
rect 29638 6916 29644 6928
rect 23615 6886 23649 6914
rect 23768 6888 29644 6916
rect 23615 6885 23627 6886
rect 23569 6879 23627 6885
rect 4706 6808 4712 6860
rect 4764 6848 4770 6860
rect 5350 6848 5356 6860
rect 4764 6820 5356 6848
rect 4764 6808 4770 6820
rect 5350 6808 5356 6820
rect 5408 6808 5414 6860
rect 7837 6851 7895 6857
rect 7837 6817 7849 6851
rect 7883 6848 7895 6851
rect 7926 6848 7932 6860
rect 7883 6820 7932 6848
rect 7883 6817 7895 6820
rect 7837 6811 7895 6817
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 10410 6808 10416 6860
rect 10468 6848 10474 6860
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 10468 6820 11529 6848
rect 10468 6808 10474 6820
rect 11517 6817 11529 6820
rect 11563 6848 11575 6851
rect 13078 6848 13084 6860
rect 11563 6820 13084 6848
rect 11563 6817 11575 6820
rect 11517 6811 11575 6817
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 16574 6848 16580 6860
rect 16071 6820 16580 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 17586 6808 17592 6860
rect 17644 6848 17650 6860
rect 20622 6848 20628 6860
rect 17644 6820 19288 6848
rect 20583 6820 20628 6848
rect 17644 6808 17650 6820
rect 5620 6783 5678 6789
rect 5620 6749 5632 6783
rect 5666 6780 5678 6783
rect 6362 6780 6368 6792
rect 5666 6752 6368 6780
rect 5666 6749 5678 6752
rect 5620 6743 5678 6749
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6780 7619 6783
rect 8386 6780 8392 6792
rect 7607 6752 8392 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 6733 6647 6791 6653
rect 6733 6613 6745 6647
rect 6779 6644 6791 6647
rect 7576 6644 7604 6743
rect 8386 6740 8392 6752
rect 8444 6740 8450 6792
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 10962 6780 10968 6792
rect 10735 6752 10968 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 10962 6740 10968 6752
rect 11020 6740 11026 6792
rect 11793 6783 11851 6789
rect 11793 6749 11805 6783
rect 11839 6780 11851 6783
rect 12342 6780 12348 6792
rect 11839 6752 12348 6780
rect 11839 6749 11851 6752
rect 11793 6743 11851 6749
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 13906 6780 13912 6792
rect 13403 6752 13912 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 16669 6783 16727 6789
rect 16448 6752 16620 6780
rect 16448 6740 16454 6752
rect 9306 6672 9312 6724
rect 9364 6712 9370 6724
rect 11701 6715 11759 6721
rect 11701 6712 11713 6715
rect 9364 6684 11713 6712
rect 9364 6672 9370 6684
rect 11701 6681 11713 6684
rect 11747 6712 11759 6715
rect 13998 6712 14004 6724
rect 11747 6684 14004 6712
rect 11747 6681 11759 6684
rect 11701 6675 11759 6681
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 14185 6715 14243 6721
rect 14185 6681 14197 6715
rect 14231 6712 14243 6715
rect 14458 6712 14464 6724
rect 14231 6684 14464 6712
rect 14231 6681 14243 6684
rect 14185 6675 14243 6681
rect 14458 6672 14464 6684
rect 14516 6712 14522 6724
rect 15194 6712 15200 6724
rect 14516 6684 15200 6712
rect 14516 6672 14522 6684
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 15780 6715 15838 6721
rect 15780 6681 15792 6715
rect 15826 6712 15838 6715
rect 16592 6712 16620 6752
rect 16669 6749 16681 6783
rect 16715 6780 16727 6783
rect 16758 6780 16764 6792
rect 16715 6752 16764 6780
rect 16715 6749 16727 6752
rect 16669 6743 16727 6749
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 18046 6740 18052 6792
rect 18104 6780 18110 6792
rect 19260 6789 19288 6820
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 23584 6848 23612 6879
rect 26528 6857 26556 6888
rect 26513 6851 26571 6857
rect 23124 6820 23612 6848
rect 23860 6820 24900 6848
rect 18509 6783 18567 6789
rect 18509 6780 18521 6783
rect 18104 6752 18521 6780
rect 18104 6740 18110 6752
rect 18509 6749 18521 6752
rect 18555 6749 18567 6783
rect 18509 6743 18567 6749
rect 19245 6783 19303 6789
rect 19245 6749 19257 6783
rect 19291 6749 19303 6783
rect 20254 6780 20260 6792
rect 20215 6752 20260 6780
rect 19245 6743 19303 6749
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 20441 6783 20499 6789
rect 20441 6749 20453 6783
rect 20487 6780 20499 6783
rect 21174 6780 21180 6792
rect 20487 6752 21180 6780
rect 20487 6749 20499 6752
rect 20441 6743 20499 6749
rect 21174 6740 21180 6752
rect 21232 6740 21238 6792
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6780 21603 6783
rect 22186 6780 22192 6792
rect 21591 6752 22192 6780
rect 21591 6749 21603 6752
rect 21545 6743 21603 6749
rect 22186 6740 22192 6752
rect 22244 6740 22250 6792
rect 23124 6789 23152 6820
rect 22925 6783 22983 6789
rect 22925 6749 22937 6783
rect 22971 6749 22983 6783
rect 22925 6743 22983 6749
rect 23109 6783 23167 6789
rect 23109 6749 23121 6783
rect 23155 6749 23167 6783
rect 23109 6743 23167 6749
rect 17129 6715 17187 6721
rect 17129 6712 17141 6715
rect 15826 6684 16528 6712
rect 16592 6684 17141 6712
rect 15826 6681 15838 6684
rect 15780 6675 15838 6681
rect 6779 6616 7604 6644
rect 6779 6613 6791 6616
rect 6733 6607 6791 6613
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 10042 6644 10048 6656
rect 7708 6616 7753 6644
rect 10003 6616 10048 6644
rect 7708 6604 7714 6616
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 10318 6604 10324 6656
rect 10376 6644 10382 6656
rect 10505 6647 10563 6653
rect 10505 6644 10517 6647
rect 10376 6616 10517 6644
rect 10376 6604 10382 6616
rect 10505 6613 10517 6616
rect 10551 6613 10563 6647
rect 10505 6607 10563 6613
rect 12066 6604 12072 6656
rect 12124 6644 12130 6656
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 12124 6616 12173 6644
rect 12124 6604 12130 6616
rect 12161 6613 12173 6616
rect 12207 6613 12219 6647
rect 12802 6644 12808 6656
rect 12763 6616 12808 6644
rect 12161 6607 12219 6613
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 13541 6647 13599 6653
rect 13541 6613 13553 6647
rect 13587 6644 13599 6647
rect 13630 6644 13636 6656
rect 13587 6616 13636 6644
rect 13587 6613 13599 6616
rect 13541 6607 13599 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 14645 6647 14703 6653
rect 14645 6613 14657 6647
rect 14691 6644 14703 6647
rect 15470 6644 15476 6656
rect 14691 6616 15476 6644
rect 14691 6613 14703 6616
rect 14645 6607 14703 6613
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 16500 6653 16528 6684
rect 17129 6681 17141 6684
rect 17175 6681 17187 6715
rect 19334 6712 19340 6724
rect 17129 6675 17187 6681
rect 18708 6684 19340 6712
rect 18708 6653 18736 6684
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 22940 6712 22968 6743
rect 23198 6740 23204 6792
rect 23256 6780 23262 6792
rect 23860 6789 23888 6820
rect 23845 6783 23903 6789
rect 23845 6780 23857 6783
rect 23256 6752 23857 6780
rect 23256 6740 23262 6752
rect 23845 6749 23857 6752
rect 23891 6749 23903 6783
rect 23845 6743 23903 6749
rect 24026 6740 24032 6792
rect 24084 6780 24090 6792
rect 24084 6752 24808 6780
rect 24084 6740 24090 6752
rect 23566 6712 23572 6724
rect 22940 6684 23152 6712
rect 23527 6684 23572 6712
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6613 16543 6647
rect 16485 6607 16543 6613
rect 18693 6647 18751 6653
rect 18693 6613 18705 6647
rect 18739 6613 18751 6647
rect 19426 6644 19432 6656
rect 19387 6616 19432 6644
rect 18693 6607 18751 6613
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 23014 6644 23020 6656
rect 22975 6616 23020 6644
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 23124 6644 23152 6684
rect 23566 6672 23572 6684
rect 23624 6672 23630 6724
rect 24780 6721 24808 6752
rect 24765 6715 24823 6721
rect 23676 6684 24440 6712
rect 23382 6644 23388 6656
rect 23124 6616 23388 6644
rect 23382 6604 23388 6616
rect 23440 6644 23446 6656
rect 23676 6644 23704 6684
rect 23440 6616 23704 6644
rect 23753 6647 23811 6653
rect 23440 6604 23446 6616
rect 23753 6613 23765 6647
rect 23799 6644 23811 6647
rect 23934 6644 23940 6656
rect 23799 6616 23940 6644
rect 23799 6613 23811 6616
rect 23753 6607 23811 6613
rect 23934 6604 23940 6616
rect 23992 6604 23998 6656
rect 24412 6653 24440 6684
rect 24765 6681 24777 6715
rect 24811 6681 24823 6715
rect 24872 6712 24900 6820
rect 26513 6817 26525 6851
rect 26559 6817 26571 6851
rect 26513 6811 26571 6817
rect 26697 6851 26755 6857
rect 26697 6817 26709 6851
rect 26743 6848 26755 6851
rect 27338 6848 27344 6860
rect 26743 6820 27344 6848
rect 26743 6817 26755 6820
rect 26697 6811 26755 6817
rect 27338 6808 27344 6820
rect 27396 6808 27402 6860
rect 28368 6857 28396 6888
rect 29638 6876 29644 6888
rect 29696 6876 29702 6928
rect 32122 6876 32128 6928
rect 32180 6916 32186 6928
rect 32766 6916 32772 6928
rect 32180 6888 32772 6916
rect 32180 6876 32186 6888
rect 32766 6876 32772 6888
rect 32824 6916 32830 6928
rect 33045 6919 33103 6925
rect 33045 6916 33057 6919
rect 32824 6888 33057 6916
rect 32824 6876 32830 6888
rect 33045 6885 33057 6888
rect 33091 6916 33103 6919
rect 39942 6916 39948 6928
rect 33091 6888 39948 6916
rect 33091 6885 33103 6888
rect 33045 6879 33103 6885
rect 39942 6876 39948 6888
rect 40000 6876 40006 6928
rect 40034 6876 40040 6928
rect 40092 6876 40098 6928
rect 40144 6916 40172 6956
rect 40218 6944 40224 6996
rect 40276 6984 40282 6996
rect 40405 6987 40463 6993
rect 40405 6984 40417 6987
rect 40276 6956 40417 6984
rect 40276 6944 40282 6956
rect 40405 6953 40417 6956
rect 40451 6953 40463 6987
rect 40405 6947 40463 6953
rect 40494 6944 40500 6996
rect 40552 6984 40558 6996
rect 45186 6984 45192 6996
rect 40552 6956 45192 6984
rect 40552 6944 40558 6956
rect 45186 6944 45192 6956
rect 45244 6944 45250 6996
rect 45554 6916 45560 6928
rect 40144 6888 45560 6916
rect 45554 6876 45560 6888
rect 45612 6916 45618 6928
rect 49970 6916 49976 6928
rect 45612 6888 45692 6916
rect 45612 6876 45618 6888
rect 28353 6851 28411 6857
rect 28353 6817 28365 6851
rect 28399 6848 28411 6851
rect 28399 6820 28433 6848
rect 28399 6817 28411 6820
rect 28353 6811 28411 6817
rect 28626 6808 28632 6860
rect 28684 6848 28690 6860
rect 35618 6848 35624 6860
rect 28684 6820 35624 6848
rect 28684 6808 28690 6820
rect 35618 6808 35624 6820
rect 35676 6808 35682 6860
rect 40052 6848 40080 6876
rect 40129 6851 40187 6857
rect 40129 6848 40141 6851
rect 40052 6820 40141 6848
rect 40129 6817 40141 6820
rect 40175 6848 40187 6851
rect 41138 6848 41144 6860
rect 40175 6820 41144 6848
rect 40175 6817 40187 6820
rect 40129 6811 40187 6817
rect 41138 6808 41144 6820
rect 41196 6808 41202 6860
rect 45002 6808 45008 6860
rect 45060 6848 45066 6860
rect 45097 6851 45155 6857
rect 45097 6848 45109 6851
rect 45060 6820 45109 6848
rect 45060 6808 45066 6820
rect 45097 6817 45109 6820
rect 45143 6817 45155 6851
rect 45097 6811 45155 6817
rect 25222 6780 25228 6792
rect 25183 6752 25228 6780
rect 25222 6740 25228 6752
rect 25280 6740 25286 6792
rect 26418 6780 26424 6792
rect 26379 6752 26424 6780
rect 26418 6740 26424 6752
rect 26476 6740 26482 6792
rect 29270 6780 29276 6792
rect 26528 6752 29276 6780
rect 26528 6712 26556 6752
rect 29270 6740 29276 6752
rect 29328 6740 29334 6792
rect 29638 6740 29644 6792
rect 29696 6780 29702 6792
rect 29733 6783 29791 6789
rect 29733 6780 29745 6783
rect 29696 6752 29745 6780
rect 29696 6740 29702 6752
rect 29733 6749 29745 6752
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 34790 6740 34796 6792
rect 34848 6780 34854 6792
rect 34885 6783 34943 6789
rect 34885 6780 34897 6783
rect 34848 6752 34897 6780
rect 34848 6740 34854 6752
rect 34885 6749 34897 6752
rect 34931 6780 34943 6783
rect 35342 6780 35348 6792
rect 34931 6752 35348 6780
rect 34931 6749 34943 6752
rect 34885 6743 34943 6749
rect 35342 6740 35348 6752
rect 35400 6740 35406 6792
rect 40037 6783 40095 6789
rect 40037 6749 40049 6783
rect 40083 6780 40095 6783
rect 40494 6780 40500 6792
rect 40083 6752 40500 6780
rect 40083 6749 40095 6752
rect 40037 6743 40095 6749
rect 40494 6740 40500 6752
rect 40552 6740 40558 6792
rect 41874 6740 41880 6792
rect 41932 6780 41938 6792
rect 43809 6783 43867 6789
rect 43809 6780 43821 6783
rect 41932 6752 43821 6780
rect 41932 6740 41938 6752
rect 43809 6749 43821 6752
rect 43855 6749 43867 6783
rect 43990 6780 43996 6792
rect 43951 6752 43996 6780
rect 43809 6743 43867 6749
rect 43990 6740 43996 6752
rect 44048 6740 44054 6792
rect 44266 6789 44272 6792
rect 44223 6783 44272 6789
rect 44223 6749 44235 6783
rect 44269 6749 44272 6783
rect 44223 6743 44272 6749
rect 44266 6740 44272 6743
rect 44324 6740 44330 6792
rect 24872 6684 26556 6712
rect 24765 6675 24823 6681
rect 27154 6672 27160 6724
rect 27212 6712 27218 6724
rect 27801 6715 27859 6721
rect 27801 6712 27813 6715
rect 27212 6684 27813 6712
rect 27212 6672 27218 6684
rect 27801 6681 27813 6684
rect 27847 6681 27859 6715
rect 27801 6675 27859 6681
rect 28718 6672 28724 6724
rect 28776 6712 28782 6724
rect 30650 6712 30656 6724
rect 28776 6684 30656 6712
rect 28776 6672 28782 6684
rect 30650 6672 30656 6684
rect 30708 6672 30714 6724
rect 40678 6712 40684 6724
rect 31726 6684 40684 6712
rect 24397 6647 24455 6653
rect 24397 6613 24409 6647
rect 24443 6613 24455 6647
rect 24397 6607 24455 6613
rect 24565 6647 24623 6653
rect 24565 6613 24577 6647
rect 24611 6644 24623 6647
rect 24946 6644 24952 6656
rect 24611 6616 24952 6644
rect 24611 6613 24623 6616
rect 24565 6607 24623 6613
rect 24946 6604 24952 6616
rect 25004 6604 25010 6656
rect 25222 6604 25228 6656
rect 25280 6644 25286 6656
rect 25317 6647 25375 6653
rect 25317 6644 25329 6647
rect 25280 6616 25329 6644
rect 25280 6604 25286 6616
rect 25317 6613 25329 6616
rect 25363 6613 25375 6647
rect 26050 6644 26056 6656
rect 26011 6616 26056 6644
rect 25317 6607 25375 6613
rect 26050 6604 26056 6616
rect 26108 6604 26114 6656
rect 27246 6644 27252 6656
rect 27207 6616 27252 6644
rect 27246 6604 27252 6616
rect 27304 6604 27310 6656
rect 29917 6647 29975 6653
rect 29917 6613 29929 6647
rect 29963 6644 29975 6647
rect 30282 6644 30288 6656
rect 29963 6616 30288 6644
rect 29963 6613 29975 6616
rect 29917 6607 29975 6613
rect 30282 6604 30288 6616
rect 30340 6604 30346 6656
rect 30469 6647 30527 6653
rect 30469 6613 30481 6647
rect 30515 6644 30527 6647
rect 31110 6644 31116 6656
rect 30515 6616 31116 6644
rect 30515 6613 30527 6616
rect 30469 6607 30527 6613
rect 31110 6604 31116 6616
rect 31168 6644 31174 6656
rect 31726 6644 31754 6684
rect 40678 6672 40684 6684
rect 40736 6672 40742 6724
rect 44085 6715 44143 6721
rect 44085 6681 44097 6715
rect 44131 6712 44143 6715
rect 45020 6712 45048 6808
rect 45186 6780 45192 6792
rect 45099 6752 45192 6780
rect 45186 6740 45192 6752
rect 45244 6740 45250 6792
rect 45664 6789 45692 6888
rect 49617 6888 49976 6916
rect 48406 6848 48412 6860
rect 47872 6820 48412 6848
rect 45649 6783 45707 6789
rect 45649 6749 45661 6783
rect 45695 6749 45707 6783
rect 45649 6743 45707 6749
rect 44131 6684 45048 6712
rect 45204 6712 45232 6740
rect 47486 6712 47492 6724
rect 45204 6684 47492 6712
rect 44131 6681 44143 6684
rect 44085 6675 44143 6681
rect 47486 6672 47492 6684
rect 47544 6672 47550 6724
rect 47872 6712 47900 6820
rect 48406 6808 48412 6820
rect 48464 6848 48470 6860
rect 48590 6848 48596 6860
rect 48464 6820 48596 6848
rect 48464 6808 48470 6820
rect 48590 6808 48596 6820
rect 48648 6808 48654 6860
rect 49617 6857 49645 6888
rect 49970 6876 49976 6888
rect 50028 6876 50034 6928
rect 49605 6851 49663 6857
rect 49605 6817 49617 6851
rect 49651 6817 49663 6851
rect 50801 6851 50859 6857
rect 50801 6848 50813 6851
rect 49605 6811 49663 6817
rect 49712 6820 50813 6848
rect 47949 6783 48007 6789
rect 47949 6749 47961 6783
rect 47995 6780 48007 6783
rect 48314 6780 48320 6792
rect 47995 6752 48320 6780
rect 47995 6749 48007 6752
rect 47949 6743 48007 6749
rect 48314 6740 48320 6752
rect 48372 6740 48378 6792
rect 49329 6783 49387 6789
rect 49329 6749 49341 6783
rect 49375 6749 49387 6783
rect 49329 6743 49387 6749
rect 48133 6715 48191 6721
rect 48133 6712 48145 6715
rect 47872 6684 48145 6712
rect 48133 6681 48145 6684
rect 48179 6681 48191 6715
rect 49344 6712 49372 6743
rect 49418 6740 49424 6792
rect 49476 6780 49482 6792
rect 49712 6780 49740 6820
rect 50801 6817 50813 6820
rect 50847 6817 50859 6851
rect 50801 6811 50859 6817
rect 50341 6783 50399 6789
rect 50341 6780 50353 6783
rect 49476 6752 49740 6780
rect 49804 6752 50353 6780
rect 49476 6740 49482 6752
rect 49694 6712 49700 6724
rect 48133 6675 48191 6681
rect 48424 6684 49280 6712
rect 49344 6684 49700 6712
rect 43346 6644 43352 6656
rect 31168 6616 31754 6644
rect 43307 6616 43352 6644
rect 31168 6604 31174 6616
rect 43346 6604 43352 6616
rect 43404 6604 43410 6656
rect 44174 6604 44180 6656
rect 44232 6644 44238 6656
rect 44361 6647 44419 6653
rect 44361 6644 44373 6647
rect 44232 6616 44373 6644
rect 44232 6604 44238 6616
rect 44361 6613 44373 6616
rect 44407 6613 44419 6647
rect 45738 6644 45744 6656
rect 45699 6616 45744 6644
rect 44361 6607 44419 6613
rect 45738 6604 45744 6616
rect 45796 6604 45802 6656
rect 47765 6647 47823 6653
rect 47765 6613 47777 6647
rect 47811 6644 47823 6647
rect 48424 6644 48452 6684
rect 47811 6616 48452 6644
rect 47811 6613 47823 6616
rect 47765 6607 47823 6613
rect 48498 6604 48504 6656
rect 48556 6644 48562 6656
rect 48593 6647 48651 6653
rect 48593 6644 48605 6647
rect 48556 6616 48605 6644
rect 48556 6604 48562 6616
rect 48593 6613 48605 6616
rect 48639 6613 48651 6647
rect 49252 6644 49280 6684
rect 49694 6672 49700 6684
rect 49752 6672 49758 6724
rect 49804 6644 49832 6752
rect 50341 6749 50353 6752
rect 50387 6749 50399 6783
rect 50341 6743 50399 6749
rect 49252 6616 49832 6644
rect 48593 6607 48651 6613
rect 49970 6604 49976 6656
rect 50028 6644 50034 6656
rect 50157 6647 50215 6653
rect 50157 6644 50169 6647
rect 50028 6616 50169 6644
rect 50028 6604 50034 6616
rect 50157 6613 50169 6616
rect 50203 6613 50215 6647
rect 50157 6607 50215 6613
rect 1104 6554 68816 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 68816 6554
rect 1104 6480 68816 6502
rect 7285 6443 7343 6449
rect 7285 6409 7297 6443
rect 7331 6440 7343 6443
rect 8294 6440 8300 6452
rect 7331 6412 8300 6440
rect 7331 6409 7343 6412
rect 7285 6403 7343 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 9306 6440 9312 6452
rect 9267 6412 9312 6440
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 9401 6443 9459 6449
rect 9401 6409 9413 6443
rect 9447 6440 9459 6443
rect 10502 6440 10508 6452
rect 9447 6412 10508 6440
rect 9447 6409 9459 6412
rect 9401 6403 9459 6409
rect 10502 6400 10508 6412
rect 10560 6400 10566 6452
rect 10962 6440 10968 6452
rect 10923 6412 10968 6440
rect 10962 6400 10968 6412
rect 11020 6400 11026 6452
rect 12342 6400 12348 6452
rect 12400 6440 12406 6452
rect 12897 6443 12955 6449
rect 12897 6440 12909 6443
rect 12400 6412 12909 6440
rect 12400 6400 12406 6412
rect 12897 6409 12909 6412
rect 12943 6409 12955 6443
rect 14734 6440 14740 6452
rect 14695 6412 14740 6440
rect 12897 6403 12955 6409
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 17402 6400 17408 6452
rect 17460 6440 17466 6452
rect 17586 6440 17592 6452
rect 17460 6412 17592 6440
rect 17460 6400 17466 6412
rect 17586 6400 17592 6412
rect 17644 6400 17650 6452
rect 18046 6440 18052 6452
rect 18007 6412 18052 6440
rect 18046 6400 18052 6412
rect 18104 6400 18110 6452
rect 19426 6400 19432 6452
rect 19484 6440 19490 6452
rect 25593 6443 25651 6449
rect 19484 6412 25452 6440
rect 19484 6400 19490 6412
rect 7377 6375 7435 6381
rect 7377 6341 7389 6375
rect 7423 6372 7435 6375
rect 7650 6372 7656 6384
rect 7423 6344 7656 6372
rect 7423 6341 7435 6344
rect 7377 6335 7435 6341
rect 7650 6332 7656 6344
rect 7708 6372 7714 6384
rect 8205 6375 8263 6381
rect 8205 6372 8217 6375
rect 7708 6344 8217 6372
rect 7708 6332 7714 6344
rect 8205 6341 8217 6344
rect 8251 6372 8263 6375
rect 10597 6375 10655 6381
rect 8251 6344 10088 6372
rect 8251 6341 8263 6344
rect 8205 6335 8263 6341
rect 10060 6316 10088 6344
rect 10597 6341 10609 6375
rect 10643 6372 10655 6375
rect 11422 6372 11428 6384
rect 10643 6344 11428 6372
rect 10643 6341 10655 6344
rect 10597 6335 10655 6341
rect 11422 6332 11428 6344
rect 11480 6332 11486 6384
rect 11514 6332 11520 6384
rect 11572 6372 11578 6384
rect 11572 6344 12434 6372
rect 11572 6332 11578 6344
rect 10042 6264 10048 6316
rect 10100 6304 10106 6316
rect 10100 6276 10548 6304
rect 10100 6264 10106 6276
rect 6454 6196 6460 6248
rect 6512 6236 6518 6248
rect 7469 6239 7527 6245
rect 7469 6236 7481 6239
rect 6512 6208 7481 6236
rect 6512 6196 6518 6208
rect 7469 6205 7481 6208
rect 7515 6236 7527 6239
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 7515 6208 9137 6236
rect 7515 6205 7527 6208
rect 7469 6199 7527 6205
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 10410 6236 10416 6248
rect 10371 6208 10416 6236
rect 9125 6199 9183 6205
rect 10410 6196 10416 6208
rect 10468 6196 10474 6248
rect 10520 6245 10548 6276
rect 11606 6264 11612 6316
rect 11664 6304 11670 6316
rect 11773 6307 11831 6313
rect 11773 6304 11785 6307
rect 11664 6276 11785 6304
rect 11664 6264 11670 6276
rect 11773 6273 11785 6276
rect 11819 6273 11831 6307
rect 12406 6304 12434 6344
rect 13998 6332 14004 6384
rect 14056 6372 14062 6384
rect 19794 6372 19800 6384
rect 14056 6344 19800 6372
rect 14056 6332 14062 6344
rect 13630 6313 13636 6316
rect 13357 6307 13415 6313
rect 13357 6304 13369 6307
rect 12406 6276 13369 6304
rect 11773 6267 11831 6273
rect 13357 6273 13369 6276
rect 13403 6273 13415 6307
rect 13624 6304 13636 6313
rect 13591 6276 13636 6304
rect 13357 6267 13415 6273
rect 13624 6267 13636 6276
rect 13630 6264 13636 6267
rect 13688 6264 13694 6316
rect 15194 6304 15200 6316
rect 15155 6276 15200 6304
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 15488 6313 15516 6344
rect 19794 6332 19800 6344
rect 19852 6332 19858 6384
rect 20990 6372 20996 6384
rect 20951 6344 20996 6372
rect 20990 6332 20996 6344
rect 21048 6372 21054 6384
rect 22189 6375 22247 6381
rect 22189 6372 22201 6375
rect 21048 6344 22201 6372
rect 21048 6332 21054 6344
rect 22189 6341 22201 6344
rect 22235 6341 22247 6375
rect 22189 6335 22247 6341
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6273 15531 6307
rect 15473 6267 15531 6273
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6304 17739 6307
rect 17954 6304 17960 6316
rect 17727 6276 17960 6304
rect 17727 6273 17739 6276
rect 17681 6267 17739 6273
rect 17954 6264 17960 6276
rect 18012 6304 18018 6316
rect 18506 6304 18512 6316
rect 18012 6276 18512 6304
rect 18012 6264 18018 6276
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 19061 6307 19119 6313
rect 19061 6273 19073 6307
rect 19107 6304 19119 6307
rect 19150 6304 19156 6316
rect 19107 6276 19156 6304
rect 19107 6273 19119 6276
rect 19061 6267 19119 6273
rect 19150 6264 19156 6276
rect 19208 6264 19214 6316
rect 22204 6304 22232 6335
rect 23014 6332 23020 6384
rect 23072 6372 23078 6384
rect 24121 6375 24179 6381
rect 24121 6372 24133 6375
rect 23072 6344 24133 6372
rect 23072 6332 23078 6344
rect 24121 6341 24133 6344
rect 24167 6341 24179 6375
rect 25424 6372 25452 6412
rect 25593 6409 25605 6443
rect 25639 6440 25651 6443
rect 27617 6443 27675 6449
rect 25639 6412 27476 6440
rect 25639 6409 25651 6412
rect 25593 6403 25651 6409
rect 27338 6372 27344 6384
rect 25424 6344 27344 6372
rect 24121 6335 24179 6341
rect 27338 6332 27344 6344
rect 27396 6332 27402 6384
rect 23293 6307 23351 6313
rect 23293 6304 23305 6307
rect 22204 6276 23305 6304
rect 23293 6273 23305 6276
rect 23339 6304 23351 6307
rect 23566 6304 23572 6316
rect 23339 6276 23572 6304
rect 23339 6273 23351 6276
rect 23293 6267 23351 6273
rect 23566 6264 23572 6276
rect 23624 6264 23630 6316
rect 25222 6264 25228 6316
rect 25280 6264 25286 6316
rect 27448 6304 27476 6412
rect 27617 6409 27629 6443
rect 27663 6440 27675 6443
rect 27982 6440 27988 6452
rect 27663 6412 27988 6440
rect 27663 6409 27675 6412
rect 27617 6403 27675 6409
rect 27982 6400 27988 6412
rect 28040 6400 28046 6452
rect 29638 6440 29644 6452
rect 29599 6412 29644 6440
rect 29638 6400 29644 6412
rect 29696 6400 29702 6452
rect 31573 6443 31631 6449
rect 31573 6409 31585 6443
rect 31619 6440 31631 6443
rect 32122 6440 32128 6452
rect 31619 6412 32128 6440
rect 31619 6409 31631 6412
rect 31573 6403 31631 6409
rect 32122 6400 32128 6412
rect 32180 6400 32186 6452
rect 34790 6440 34796 6452
rect 34751 6412 34796 6440
rect 34790 6400 34796 6412
rect 34848 6400 34854 6452
rect 41874 6440 41880 6452
rect 41835 6412 41880 6440
rect 41874 6400 41880 6412
rect 41932 6400 41938 6452
rect 43346 6400 43352 6452
rect 43404 6440 43410 6452
rect 44266 6440 44272 6452
rect 43404 6412 44272 6440
rect 43404 6400 43410 6412
rect 44266 6400 44272 6412
rect 44324 6440 44330 6452
rect 45649 6443 45707 6449
rect 45649 6440 45661 6443
rect 44324 6412 45661 6440
rect 44324 6400 44330 6412
rect 45649 6409 45661 6412
rect 45695 6440 45707 6443
rect 45695 6412 51074 6440
rect 45695 6409 45707 6412
rect 45649 6403 45707 6409
rect 27522 6332 27528 6384
rect 27580 6372 27586 6384
rect 28442 6372 28448 6384
rect 27580 6344 28448 6372
rect 27580 6332 27586 6344
rect 28442 6332 28448 6344
rect 28500 6372 28506 6384
rect 33318 6372 33324 6384
rect 28500 6344 31754 6372
rect 33279 6344 33324 6372
rect 28500 6332 28506 6344
rect 27706 6304 27712 6316
rect 27448 6276 27712 6304
rect 27706 6264 27712 6276
rect 27764 6264 27770 6316
rect 28718 6264 28724 6316
rect 28776 6304 28782 6316
rect 29181 6307 29239 6313
rect 29181 6304 29193 6307
rect 28776 6276 29193 6304
rect 28776 6264 28782 6276
rect 29181 6273 29193 6276
rect 29227 6273 29239 6307
rect 29181 6267 29239 6273
rect 29270 6264 29276 6316
rect 29328 6304 29334 6316
rect 30208 6313 30236 6344
rect 31726 6316 31754 6344
rect 33318 6332 33324 6344
rect 33376 6332 33382 6384
rect 33870 6332 33876 6384
rect 33928 6332 33934 6384
rect 44174 6372 44180 6384
rect 44135 6344 44180 6372
rect 44174 6332 44180 6344
rect 44232 6332 44238 6384
rect 45738 6372 45744 6384
rect 45402 6344 45744 6372
rect 45738 6332 45744 6344
rect 45796 6332 45802 6384
rect 50062 6332 50068 6384
rect 50120 6332 50126 6384
rect 30193 6307 30251 6313
rect 29328 6276 29421 6304
rect 29328 6264 29334 6276
rect 30193 6273 30205 6307
rect 30239 6273 30251 6307
rect 30193 6267 30251 6273
rect 30282 6264 30288 6316
rect 30340 6304 30346 6316
rect 30449 6307 30507 6313
rect 30449 6304 30461 6307
rect 30340 6276 30461 6304
rect 30340 6264 30346 6276
rect 30449 6273 30461 6276
rect 30495 6273 30507 6307
rect 31726 6276 31760 6316
rect 30449 6267 30507 6273
rect 31754 6264 31760 6276
rect 31812 6304 31818 6316
rect 32582 6304 32588 6316
rect 31812 6276 32588 6304
rect 31812 6264 31818 6276
rect 32582 6264 32588 6276
rect 32640 6304 32646 6316
rect 33045 6307 33103 6313
rect 33045 6304 33057 6307
rect 32640 6276 33057 6304
rect 32640 6264 32646 6276
rect 33045 6273 33057 6276
rect 33091 6273 33103 6307
rect 33045 6267 33103 6273
rect 37461 6307 37519 6313
rect 37461 6273 37473 6307
rect 37507 6304 37519 6307
rect 38654 6304 38660 6316
rect 37507 6276 38660 6304
rect 37507 6273 37519 6276
rect 37461 6267 37519 6273
rect 38654 6264 38660 6276
rect 38712 6264 38718 6316
rect 40954 6264 40960 6316
rect 41012 6313 41018 6316
rect 41012 6307 41033 6313
rect 41021 6273 41033 6307
rect 41230 6304 41236 6316
rect 41191 6276 41236 6304
rect 41012 6267 41033 6273
rect 41012 6264 41018 6267
rect 41230 6264 41236 6276
rect 41288 6264 41294 6316
rect 48314 6304 48320 6316
rect 48275 6276 48320 6304
rect 48314 6264 48320 6276
rect 48372 6264 48378 6316
rect 48958 6264 48964 6316
rect 49016 6304 49022 6316
rect 49053 6307 49111 6313
rect 49053 6304 49065 6307
rect 49016 6276 49065 6304
rect 49016 6264 49022 6276
rect 49053 6273 49065 6276
rect 49099 6273 49111 6307
rect 49878 6304 49884 6316
rect 49839 6276 49884 6304
rect 49053 6267 49111 6273
rect 49878 6264 49884 6276
rect 49936 6264 49942 6316
rect 50080 6304 50108 6332
rect 50157 6307 50215 6313
rect 50157 6304 50169 6307
rect 50080 6276 50169 6304
rect 50157 6273 50169 6276
rect 50203 6304 50215 6307
rect 50617 6307 50675 6313
rect 50617 6304 50629 6307
rect 50203 6276 50629 6304
rect 50203 6273 50215 6276
rect 50157 6267 50215 6273
rect 50617 6273 50629 6276
rect 50663 6273 50675 6307
rect 50617 6267 50675 6273
rect 10505 6239 10563 6245
rect 10505 6205 10517 6239
rect 10551 6236 10563 6239
rect 11054 6236 11060 6248
rect 10551 6208 11060 6236
rect 10551 6205 10563 6208
rect 10505 6199 10563 6205
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 11514 6236 11520 6248
rect 11475 6208 11520 6236
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 16758 6196 16764 6248
rect 16816 6236 16822 6248
rect 17402 6236 17408 6248
rect 16816 6208 17408 6236
rect 16816 6196 16822 6208
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 17589 6239 17647 6245
rect 17589 6205 17601 6239
rect 17635 6205 17647 6239
rect 17589 6199 17647 6205
rect 17604 6168 17632 6199
rect 22186 6196 22192 6248
rect 22244 6236 22250 6248
rect 22833 6239 22891 6245
rect 22833 6236 22845 6239
rect 22244 6208 22845 6236
rect 22244 6196 22250 6208
rect 22833 6205 22845 6208
rect 22879 6236 22891 6239
rect 23198 6236 23204 6248
rect 22879 6208 23204 6236
rect 22879 6205 22891 6208
rect 22833 6199 22891 6205
rect 23198 6196 23204 6208
rect 23256 6196 23262 6248
rect 23845 6239 23903 6245
rect 23845 6205 23857 6239
rect 23891 6205 23903 6239
rect 23845 6199 23903 6205
rect 15028 6140 17632 6168
rect 6914 6100 6920 6112
rect 6875 6072 6920 6100
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 9769 6103 9827 6109
rect 9769 6100 9781 6103
rect 9548 6072 9781 6100
rect 9548 6060 9554 6072
rect 9769 6069 9781 6072
rect 9815 6069 9827 6103
rect 9769 6063 9827 6069
rect 12158 6060 12164 6112
rect 12216 6100 12222 6112
rect 15028 6100 15056 6140
rect 12216 6072 15056 6100
rect 12216 6060 12222 6072
rect 16574 6060 16580 6112
rect 16632 6100 16638 6112
rect 16669 6103 16727 6109
rect 16669 6100 16681 6103
rect 16632 6072 16681 6100
rect 16632 6060 16638 6072
rect 16669 6069 16681 6072
rect 16715 6069 16727 6103
rect 16669 6063 16727 6069
rect 19245 6103 19303 6109
rect 19245 6069 19257 6103
rect 19291 6100 19303 6103
rect 19334 6100 19340 6112
rect 19291 6072 19340 6100
rect 19291 6069 19303 6072
rect 19245 6063 19303 6069
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 23860 6100 23888 6199
rect 27338 6196 27344 6248
rect 27396 6236 27402 6248
rect 27433 6239 27491 6245
rect 27433 6236 27445 6239
rect 27396 6208 27445 6236
rect 27396 6196 27402 6208
rect 27433 6205 27445 6208
rect 27479 6205 27491 6239
rect 27433 6199 27491 6205
rect 27525 6239 27583 6245
rect 27525 6205 27537 6239
rect 27571 6236 27583 6239
rect 27614 6236 27620 6248
rect 27571 6208 27620 6236
rect 27571 6205 27583 6208
rect 27525 6199 27583 6205
rect 26418 6168 26424 6180
rect 25148 6140 26424 6168
rect 25148 6100 25176 6140
rect 26418 6128 26424 6140
rect 26476 6128 26482 6180
rect 27448 6168 27476 6199
rect 27614 6196 27620 6208
rect 27672 6236 27678 6248
rect 28810 6236 28816 6248
rect 27672 6208 28816 6236
rect 27672 6196 27678 6208
rect 28810 6196 28816 6208
rect 28868 6196 28874 6248
rect 28997 6239 29055 6245
rect 28997 6205 29009 6239
rect 29043 6205 29055 6239
rect 28997 6199 29055 6205
rect 29012 6168 29040 6199
rect 27448 6140 29040 6168
rect 23860 6072 25176 6100
rect 26234 6060 26240 6112
rect 26292 6100 26298 6112
rect 26329 6103 26387 6109
rect 26329 6100 26341 6103
rect 26292 6072 26341 6100
rect 26292 6060 26298 6072
rect 26329 6069 26341 6072
rect 26375 6100 26387 6103
rect 27614 6100 27620 6112
rect 26375 6072 27620 6100
rect 26375 6069 26387 6072
rect 26329 6063 26387 6069
rect 27614 6060 27620 6072
rect 27672 6060 27678 6112
rect 27982 6100 27988 6112
rect 27943 6072 27988 6100
rect 27982 6060 27988 6072
rect 28040 6060 28046 6112
rect 29288 6100 29316 6264
rect 40034 6236 40040 6248
rect 39995 6208 40040 6236
rect 40034 6196 40040 6208
rect 40092 6196 40098 6248
rect 40218 6236 40224 6248
rect 40179 6208 40224 6236
rect 40218 6196 40224 6208
rect 40276 6196 40282 6248
rect 40310 6196 40316 6248
rect 40368 6236 40374 6248
rect 41074 6239 41132 6245
rect 41074 6236 41086 6239
rect 40368 6208 41086 6236
rect 40368 6196 40374 6208
rect 41074 6205 41086 6208
rect 41120 6205 41132 6239
rect 41074 6199 41132 6205
rect 43714 6196 43720 6248
rect 43772 6236 43778 6248
rect 43901 6239 43959 6245
rect 43901 6236 43913 6239
rect 43772 6208 43913 6236
rect 43772 6196 43778 6208
rect 43901 6205 43913 6208
rect 43947 6205 43959 6239
rect 43901 6199 43959 6205
rect 46845 6239 46903 6245
rect 46845 6205 46857 6239
rect 46891 6236 46903 6239
rect 47118 6236 47124 6248
rect 46891 6208 47124 6236
rect 46891 6205 46903 6208
rect 46845 6199 46903 6205
rect 47118 6196 47124 6208
rect 47176 6196 47182 6248
rect 48590 6196 48596 6248
rect 48648 6236 48654 6248
rect 51046 6236 51074 6412
rect 51442 6304 51448 6316
rect 51403 6276 51448 6304
rect 51442 6264 51448 6276
rect 51500 6264 51506 6316
rect 54018 6236 54024 6248
rect 48648 6208 48693 6236
rect 51046 6208 54024 6236
rect 48648 6196 48654 6208
rect 54018 6196 54024 6208
rect 54076 6196 54082 6248
rect 40681 6171 40739 6177
rect 40681 6137 40693 6171
rect 40727 6137 40739 6171
rect 50982 6168 50988 6180
rect 40681 6131 40739 6137
rect 50816 6140 50988 6168
rect 30374 6100 30380 6112
rect 29288 6072 30380 6100
rect 30374 6060 30380 6072
rect 30432 6060 30438 6112
rect 37366 6100 37372 6112
rect 37327 6072 37372 6100
rect 37366 6060 37372 6072
rect 37424 6060 37430 6112
rect 40696 6100 40724 6131
rect 41782 6100 41788 6112
rect 40696 6072 41788 6100
rect 41782 6060 41788 6072
rect 41840 6060 41846 6112
rect 46934 6060 46940 6112
rect 46992 6100 46998 6112
rect 47581 6103 47639 6109
rect 47581 6100 47593 6103
rect 46992 6072 47593 6100
rect 46992 6060 46998 6072
rect 47581 6069 47593 6072
rect 47627 6069 47639 6103
rect 47581 6063 47639 6069
rect 50062 6060 50068 6112
rect 50120 6100 50126 6112
rect 50816 6109 50844 6140
rect 50982 6128 50988 6140
rect 51040 6128 51046 6180
rect 50801 6103 50859 6109
rect 50801 6100 50813 6103
rect 50120 6072 50813 6100
rect 50120 6060 50126 6072
rect 50801 6069 50813 6072
rect 50847 6069 50859 6103
rect 50801 6063 50859 6069
rect 50890 6060 50896 6112
rect 50948 6100 50954 6112
rect 51261 6103 51319 6109
rect 51261 6100 51273 6103
rect 50948 6072 51273 6100
rect 50948 6060 50954 6072
rect 51261 6069 51273 6072
rect 51307 6069 51319 6103
rect 51261 6063 51319 6069
rect 1104 6010 68816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 65654 6010
rect 65706 5958 65718 6010
rect 65770 5958 65782 6010
rect 65834 5958 65846 6010
rect 65898 5958 65910 6010
rect 65962 5958 68816 6010
rect 1104 5936 68816 5958
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 7745 5899 7803 5905
rect 7745 5896 7757 5899
rect 7708 5868 7757 5896
rect 7708 5856 7714 5868
rect 7745 5865 7757 5868
rect 7791 5865 7803 5899
rect 11514 5896 11520 5908
rect 7745 5859 7803 5865
rect 10060 5868 11520 5896
rect 7193 5831 7251 5837
rect 7193 5797 7205 5831
rect 7239 5828 7251 5831
rect 8294 5828 8300 5840
rect 7239 5800 8300 5828
rect 7239 5797 7251 5800
rect 7193 5791 7251 5797
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 5350 5720 5356 5772
rect 5408 5760 5414 5772
rect 10060 5769 10088 5868
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 11885 5899 11943 5905
rect 11885 5896 11897 5899
rect 11664 5868 11897 5896
rect 11664 5856 11670 5868
rect 11885 5865 11897 5868
rect 11931 5865 11943 5899
rect 26234 5896 26240 5908
rect 11885 5859 11943 5865
rect 18800 5868 26240 5896
rect 11422 5828 11428 5840
rect 11383 5800 11428 5828
rect 11422 5788 11428 5800
rect 11480 5788 11486 5840
rect 5813 5763 5871 5769
rect 5813 5760 5825 5763
rect 5408 5732 5825 5760
rect 5408 5720 5414 5732
rect 5813 5729 5825 5732
rect 5859 5729 5871 5763
rect 10045 5763 10103 5769
rect 10045 5760 10057 5763
rect 5813 5723 5871 5729
rect 9140 5732 10057 5760
rect 5828 5692 5856 5723
rect 9140 5704 9168 5732
rect 10045 5729 10057 5732
rect 10091 5729 10103 5763
rect 10045 5723 10103 5729
rect 11054 5720 11060 5772
rect 11112 5760 11118 5772
rect 15013 5763 15071 5769
rect 15013 5760 15025 5763
rect 11112 5732 15025 5760
rect 11112 5720 11118 5732
rect 15013 5729 15025 5732
rect 15059 5760 15071 5763
rect 18598 5760 18604 5772
rect 15059 5732 18604 5760
rect 15059 5729 15071 5732
rect 15013 5723 15071 5729
rect 18598 5720 18604 5732
rect 18656 5720 18662 5772
rect 9122 5692 9128 5704
rect 5828 5664 9128 5692
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 9490 5692 9496 5704
rect 9451 5664 9496 5692
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 10318 5701 10324 5704
rect 10312 5692 10324 5701
rect 10279 5664 10324 5692
rect 10312 5655 10324 5664
rect 10318 5652 10324 5655
rect 10376 5652 10382 5704
rect 12066 5692 12072 5704
rect 12027 5664 12072 5692
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 12713 5695 12771 5701
rect 12713 5692 12725 5695
rect 12492 5664 12725 5692
rect 12492 5652 12498 5664
rect 12713 5661 12725 5664
rect 12759 5661 12771 5695
rect 12713 5655 12771 5661
rect 13262 5652 13268 5704
rect 13320 5692 13326 5704
rect 13357 5695 13415 5701
rect 13357 5692 13369 5695
rect 13320 5664 13369 5692
rect 13320 5652 13326 5664
rect 13357 5661 13369 5664
rect 13403 5661 13415 5695
rect 14090 5692 14096 5704
rect 14051 5664 14096 5692
rect 13357 5655 13415 5661
rect 14090 5652 14096 5664
rect 14148 5652 14154 5704
rect 15378 5692 15384 5704
rect 14844 5664 15384 5692
rect 6080 5627 6138 5633
rect 6080 5593 6092 5627
rect 6126 5624 6138 5627
rect 6362 5624 6368 5636
rect 6126 5596 6368 5624
rect 6126 5593 6138 5596
rect 6080 5587 6138 5593
rect 6362 5584 6368 5596
rect 6420 5584 6426 5636
rect 12802 5584 12808 5636
rect 12860 5624 12866 5636
rect 14844 5633 14872 5664
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5692 17463 5695
rect 17586 5692 17592 5704
rect 17451 5664 17592 5692
rect 17451 5661 17463 5664
rect 17405 5655 17463 5661
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 18049 5695 18107 5701
rect 18049 5661 18061 5695
rect 18095 5692 18107 5695
rect 18138 5692 18144 5704
rect 18095 5664 18144 5692
rect 18095 5661 18107 5664
rect 18049 5655 18107 5661
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 18690 5692 18696 5704
rect 18651 5664 18696 5692
rect 18690 5652 18696 5664
rect 18748 5652 18754 5704
rect 14829 5627 14887 5633
rect 14829 5624 14841 5627
rect 12860 5596 14841 5624
rect 12860 5584 12866 5596
rect 14829 5593 14841 5596
rect 14875 5593 14887 5627
rect 14829 5587 14887 5593
rect 15286 5584 15292 5636
rect 15344 5624 15350 5636
rect 15565 5627 15623 5633
rect 15565 5624 15577 5627
rect 15344 5596 15577 5624
rect 15344 5584 15350 5596
rect 15565 5593 15577 5596
rect 15611 5624 15623 5627
rect 15930 5624 15936 5636
rect 15611 5596 15936 5624
rect 15611 5593 15623 5596
rect 15565 5587 15623 5593
rect 15930 5584 15936 5596
rect 15988 5624 15994 5636
rect 16117 5627 16175 5633
rect 16117 5624 16129 5627
rect 15988 5596 16129 5624
rect 15988 5584 15994 5596
rect 16117 5593 16129 5596
rect 16163 5624 16175 5627
rect 18800 5624 18828 5868
rect 26234 5856 26240 5868
rect 26292 5856 26298 5908
rect 27706 5856 27712 5908
rect 27764 5896 27770 5908
rect 27801 5899 27859 5905
rect 27801 5896 27813 5899
rect 27764 5868 27813 5896
rect 27764 5856 27770 5868
rect 27801 5865 27813 5868
rect 27847 5865 27859 5899
rect 28718 5896 28724 5908
rect 28679 5868 28724 5896
rect 27801 5859 27859 5865
rect 28718 5856 28724 5868
rect 28776 5856 28782 5908
rect 31110 5856 31116 5908
rect 31168 5856 31174 5908
rect 32766 5896 32772 5908
rect 32727 5868 32772 5896
rect 32766 5856 32772 5868
rect 32824 5856 32830 5908
rect 33870 5896 33876 5908
rect 33831 5868 33876 5896
rect 33870 5856 33876 5868
rect 33928 5856 33934 5908
rect 37458 5896 37464 5908
rect 35452 5868 37464 5896
rect 20530 5828 20536 5840
rect 19812 5800 20536 5828
rect 19812 5772 19840 5800
rect 20530 5788 20536 5800
rect 20588 5788 20594 5840
rect 20622 5788 20628 5840
rect 20680 5828 20686 5840
rect 22097 5831 22155 5837
rect 22097 5828 22109 5831
rect 20680 5800 22109 5828
rect 20680 5788 20686 5800
rect 22097 5797 22109 5800
rect 22143 5797 22155 5831
rect 22097 5791 22155 5797
rect 24581 5831 24639 5837
rect 24581 5797 24593 5831
rect 24627 5828 24639 5831
rect 24946 5828 24952 5840
rect 24627 5800 24952 5828
rect 24627 5797 24639 5800
rect 24581 5791 24639 5797
rect 19794 5760 19800 5772
rect 19755 5732 19800 5760
rect 19794 5720 19800 5732
rect 19852 5720 19858 5772
rect 19978 5760 19984 5772
rect 19939 5732 19984 5760
rect 19978 5720 19984 5732
rect 20036 5720 20042 5772
rect 19705 5695 19763 5701
rect 19705 5661 19717 5695
rect 19751 5692 19763 5695
rect 20438 5692 20444 5704
rect 19751 5664 20444 5692
rect 19751 5661 19763 5664
rect 19705 5655 19763 5661
rect 20438 5652 20444 5664
rect 20496 5652 20502 5704
rect 22112 5692 22140 5791
rect 24946 5788 24952 5800
rect 25004 5788 25010 5840
rect 25961 5831 26019 5837
rect 25961 5797 25973 5831
rect 26007 5828 26019 5831
rect 30374 5828 30380 5840
rect 26007 5800 26234 5828
rect 26007 5797 26019 5800
rect 25961 5791 26019 5797
rect 23106 5760 23112 5772
rect 23067 5732 23112 5760
rect 23106 5720 23112 5732
rect 23164 5720 23170 5772
rect 22925 5695 22983 5701
rect 22925 5692 22937 5695
rect 22112 5664 22937 5692
rect 22925 5661 22937 5664
rect 22971 5661 22983 5695
rect 22925 5655 22983 5661
rect 23017 5695 23075 5701
rect 23017 5661 23029 5695
rect 23063 5692 23075 5695
rect 24118 5692 24124 5704
rect 23063 5664 24124 5692
rect 23063 5661 23075 5664
rect 23017 5655 23075 5661
rect 24118 5652 24124 5664
rect 24176 5652 24182 5704
rect 25777 5695 25835 5701
rect 25777 5661 25789 5695
rect 25823 5692 25835 5695
rect 26050 5692 26056 5704
rect 25823 5664 26056 5692
rect 25823 5661 25835 5664
rect 25777 5655 25835 5661
rect 26050 5652 26056 5664
rect 26108 5652 26114 5704
rect 20622 5624 20628 5636
rect 16163 5596 18828 5624
rect 18892 5596 20628 5624
rect 16163 5593 16175 5596
rect 16117 5587 16175 5593
rect 9309 5559 9367 5565
rect 9309 5525 9321 5559
rect 9355 5556 9367 5559
rect 9398 5556 9404 5568
rect 9355 5528 9404 5556
rect 9355 5525 9367 5528
rect 9309 5519 9367 5525
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 12894 5556 12900 5568
rect 12855 5528 12900 5556
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 13998 5556 14004 5568
rect 13587 5528 14004 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 13998 5516 14004 5528
rect 14056 5516 14062 5568
rect 14090 5516 14096 5568
rect 14148 5556 14154 5568
rect 14277 5559 14335 5565
rect 14277 5556 14289 5559
rect 14148 5528 14289 5556
rect 14148 5516 14154 5528
rect 14277 5525 14289 5528
rect 14323 5525 14335 5559
rect 14277 5519 14335 5525
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 16209 5559 16267 5565
rect 16209 5556 16221 5559
rect 14608 5528 16221 5556
rect 14608 5516 14614 5528
rect 16209 5525 16221 5528
rect 16255 5556 16267 5559
rect 18892 5556 18920 5596
rect 20622 5584 20628 5596
rect 20680 5584 20686 5636
rect 23753 5627 23811 5633
rect 23753 5593 23765 5627
rect 23799 5624 23811 5627
rect 23934 5624 23940 5636
rect 23799 5596 23940 5624
rect 23799 5593 23811 5596
rect 23753 5587 23811 5593
rect 23934 5584 23940 5596
rect 23992 5624 23998 5636
rect 25041 5627 25099 5633
rect 25041 5624 25053 5627
rect 23992 5596 25053 5624
rect 23992 5584 23998 5596
rect 25041 5593 25053 5596
rect 25087 5624 25099 5627
rect 26206 5624 26234 5800
rect 30024 5800 30380 5828
rect 30024 5769 30052 5800
rect 30374 5788 30380 5800
rect 30432 5828 30438 5840
rect 31128 5828 31156 5856
rect 30432 5800 31156 5828
rect 30432 5788 30438 5800
rect 30009 5763 30067 5769
rect 30009 5729 30021 5763
rect 30055 5729 30067 5763
rect 30009 5723 30067 5729
rect 30285 5763 30343 5769
rect 30285 5729 30297 5763
rect 30331 5729 30343 5763
rect 30285 5723 30343 5729
rect 31021 5763 31079 5769
rect 31021 5729 31033 5763
rect 31067 5760 31079 5763
rect 31754 5760 31760 5772
rect 31067 5732 31760 5760
rect 31067 5729 31079 5732
rect 31021 5723 31079 5729
rect 26418 5692 26424 5704
rect 26331 5664 26424 5692
rect 26418 5652 26424 5664
rect 26476 5692 26482 5704
rect 27522 5692 27528 5704
rect 26476 5664 27528 5692
rect 26476 5652 26482 5664
rect 27522 5652 27528 5664
rect 27580 5652 27586 5704
rect 29917 5695 29975 5701
rect 29917 5661 29929 5695
rect 29963 5661 29975 5695
rect 29917 5655 29975 5661
rect 26666 5627 26724 5633
rect 26666 5624 26678 5627
rect 25087 5596 26096 5624
rect 26206 5596 26678 5624
rect 25087 5593 25099 5596
rect 25041 5587 25099 5593
rect 16255 5528 18920 5556
rect 19337 5559 19395 5565
rect 16255 5525 16267 5528
rect 16209 5519 16267 5525
rect 19337 5525 19349 5559
rect 19383 5556 19395 5559
rect 19426 5556 19432 5568
rect 19383 5528 19432 5556
rect 19383 5525 19395 5528
rect 19337 5519 19395 5525
rect 19426 5516 19432 5528
rect 19484 5516 19490 5568
rect 22554 5556 22560 5568
rect 22515 5528 22560 5556
rect 22554 5516 22560 5528
rect 22612 5516 22618 5568
rect 26068 5556 26096 5596
rect 26666 5593 26678 5596
rect 26712 5593 26724 5627
rect 26666 5587 26724 5593
rect 29932 5556 29960 5655
rect 30300 5624 30328 5723
rect 31754 5720 31760 5732
rect 31812 5720 31818 5772
rect 33778 5692 33784 5704
rect 33691 5664 33784 5692
rect 33778 5652 33784 5664
rect 33836 5692 33842 5704
rect 35452 5692 35480 5868
rect 37458 5856 37464 5868
rect 37516 5856 37522 5908
rect 46109 5899 46167 5905
rect 46109 5865 46121 5899
rect 46155 5896 46167 5899
rect 46290 5896 46296 5908
rect 46155 5868 46296 5896
rect 46155 5865 46167 5868
rect 46109 5859 46167 5865
rect 46290 5856 46296 5868
rect 46348 5896 46354 5908
rect 48958 5896 48964 5908
rect 46348 5868 48964 5896
rect 46348 5856 46354 5868
rect 48958 5856 48964 5868
rect 49016 5856 49022 5908
rect 49053 5899 49111 5905
rect 49053 5865 49065 5899
rect 49099 5896 49111 5899
rect 51442 5896 51448 5908
rect 49099 5868 51448 5896
rect 49099 5865 49111 5868
rect 49053 5859 49111 5865
rect 51442 5856 51448 5868
rect 51500 5856 51506 5908
rect 35529 5763 35587 5769
rect 35529 5729 35541 5763
rect 35575 5760 35587 5763
rect 35802 5760 35808 5772
rect 35575 5732 35808 5760
rect 35575 5729 35587 5732
rect 35529 5723 35587 5729
rect 35802 5720 35808 5732
rect 35860 5720 35866 5772
rect 38378 5760 38384 5772
rect 38339 5732 38384 5760
rect 38378 5720 38384 5732
rect 38436 5720 38442 5772
rect 40126 5720 40132 5772
rect 40184 5760 40190 5772
rect 40865 5763 40923 5769
rect 40865 5760 40877 5763
rect 40184 5732 40877 5760
rect 40184 5720 40190 5732
rect 40865 5729 40877 5732
rect 40911 5729 40923 5763
rect 41138 5760 41144 5772
rect 41099 5732 41144 5760
rect 40865 5723 40923 5729
rect 41138 5720 41144 5732
rect 41196 5720 41202 5772
rect 48590 5720 48596 5772
rect 48648 5760 48654 5772
rect 50062 5760 50068 5772
rect 48648 5732 50068 5760
rect 48648 5720 48654 5732
rect 50062 5720 50068 5732
rect 50120 5720 50126 5772
rect 37366 5692 37372 5704
rect 33836 5664 35480 5692
rect 36938 5664 37372 5692
rect 33836 5652 33842 5664
rect 37366 5652 37372 5664
rect 37424 5652 37430 5704
rect 39298 5692 39304 5704
rect 39259 5664 39304 5692
rect 39298 5652 39304 5664
rect 39356 5652 39362 5704
rect 40402 5692 40408 5704
rect 40363 5664 40408 5692
rect 40402 5652 40408 5664
rect 40460 5652 40466 5704
rect 46474 5652 46480 5704
rect 46532 5692 46538 5704
rect 46569 5695 46627 5701
rect 46569 5692 46581 5695
rect 46532 5664 46581 5692
rect 46532 5652 46538 5664
rect 46569 5661 46581 5664
rect 46615 5661 46627 5695
rect 46569 5655 46627 5661
rect 48317 5695 48375 5701
rect 48317 5661 48329 5695
rect 48363 5692 48375 5695
rect 48406 5692 48412 5704
rect 48363 5664 48412 5692
rect 48363 5661 48375 5664
rect 48317 5655 48375 5661
rect 48406 5652 48412 5664
rect 48464 5652 48470 5704
rect 50890 5692 50896 5704
rect 48700 5664 49556 5692
rect 50851 5664 50896 5692
rect 31297 5627 31355 5633
rect 31297 5624 31309 5627
rect 30300 5596 31309 5624
rect 31297 5593 31309 5596
rect 31343 5593 31355 5627
rect 32674 5624 32680 5636
rect 32522 5596 32680 5624
rect 31297 5587 31355 5593
rect 32674 5584 32680 5596
rect 32732 5584 32738 5636
rect 35805 5627 35863 5633
rect 35805 5593 35817 5627
rect 35851 5624 35863 5627
rect 35894 5624 35900 5636
rect 35851 5596 35900 5624
rect 35851 5593 35863 5596
rect 35805 5587 35863 5593
rect 35894 5584 35900 5596
rect 35952 5584 35958 5636
rect 39850 5584 39856 5636
rect 39908 5624 39914 5636
rect 48700 5624 48728 5664
rect 39908 5596 48728 5624
rect 49237 5627 49295 5633
rect 39908 5584 39914 5596
rect 49237 5593 49249 5627
rect 49283 5593 49295 5627
rect 49237 5587 49295 5593
rect 49421 5627 49479 5633
rect 49421 5593 49433 5627
rect 49467 5593 49479 5627
rect 49528 5624 49556 5664
rect 50890 5652 50896 5664
rect 50948 5652 50954 5704
rect 50982 5652 50988 5704
rect 51040 5692 51046 5704
rect 51169 5695 51227 5701
rect 51169 5692 51181 5695
rect 51040 5664 51181 5692
rect 51040 5652 51046 5664
rect 51169 5661 51181 5664
rect 51215 5661 51227 5695
rect 51169 5655 51227 5661
rect 55214 5624 55220 5636
rect 49528 5596 55220 5624
rect 49421 5587 49479 5593
rect 30650 5556 30656 5568
rect 26068 5528 30656 5556
rect 30650 5516 30656 5528
rect 30708 5516 30714 5568
rect 37274 5556 37280 5568
rect 37235 5528 37280 5556
rect 37274 5516 37280 5528
rect 37332 5516 37338 5568
rect 37366 5516 37372 5568
rect 37424 5556 37430 5568
rect 37737 5559 37795 5565
rect 37737 5556 37749 5559
rect 37424 5528 37749 5556
rect 37424 5516 37430 5528
rect 37737 5525 37749 5528
rect 37783 5525 37795 5559
rect 38102 5556 38108 5568
rect 38063 5528 38108 5556
rect 37737 5519 37795 5525
rect 38102 5516 38108 5528
rect 38160 5516 38166 5568
rect 38197 5559 38255 5565
rect 38197 5525 38209 5559
rect 38243 5556 38255 5559
rect 38838 5556 38844 5568
rect 38243 5528 38844 5556
rect 38243 5525 38255 5528
rect 38197 5519 38255 5525
rect 38838 5516 38844 5528
rect 38896 5516 38902 5568
rect 39758 5516 39764 5568
rect 39816 5556 39822 5568
rect 40221 5559 40279 5565
rect 40221 5556 40233 5559
rect 39816 5528 40233 5556
rect 39816 5516 39822 5528
rect 40221 5525 40233 5528
rect 40267 5525 40279 5559
rect 40221 5519 40279 5525
rect 46566 5516 46572 5568
rect 46624 5556 46630 5568
rect 47581 5559 47639 5565
rect 47581 5556 47593 5559
rect 46624 5528 47593 5556
rect 46624 5516 46630 5528
rect 47581 5525 47593 5528
rect 47627 5525 47639 5559
rect 47581 5519 47639 5525
rect 48406 5516 48412 5568
rect 48464 5556 48470 5568
rect 49252 5556 49280 5587
rect 48464 5528 49280 5556
rect 49436 5556 49464 5587
rect 55214 5584 55220 5596
rect 55272 5624 55278 5636
rect 61378 5624 61384 5636
rect 55272 5596 61384 5624
rect 55272 5584 55278 5596
rect 61378 5584 61384 5596
rect 61436 5584 61442 5636
rect 49878 5556 49884 5568
rect 49436 5528 49884 5556
rect 48464 5516 48470 5528
rect 49878 5516 49884 5528
rect 49936 5516 49942 5568
rect 50154 5556 50160 5568
rect 50115 5528 50160 5556
rect 50154 5516 50160 5528
rect 50212 5516 50218 5568
rect 51350 5516 51356 5568
rect 51408 5556 51414 5568
rect 51629 5559 51687 5565
rect 51629 5556 51641 5559
rect 51408 5528 51641 5556
rect 51408 5516 51414 5528
rect 51629 5525 51641 5528
rect 51675 5525 51687 5559
rect 51629 5519 51687 5525
rect 1104 5466 68816 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 68816 5466
rect 1104 5392 68816 5414
rect 6362 5352 6368 5364
rect 6323 5324 6368 5352
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 10502 5352 10508 5364
rect 10463 5324 10508 5352
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 18601 5355 18659 5361
rect 18601 5321 18613 5355
rect 18647 5321 18659 5355
rect 20438 5352 20444 5364
rect 20399 5324 20444 5352
rect 18601 5315 18659 5321
rect 17954 5284 17960 5296
rect 15028 5256 17960 5284
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6914 5216 6920 5228
rect 6595 5188 6920 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 9122 5216 9128 5228
rect 9083 5188 9128 5216
rect 9122 5176 9128 5188
rect 9180 5176 9186 5228
rect 9398 5225 9404 5228
rect 9392 5216 9404 5225
rect 9359 5188 9404 5216
rect 9392 5179 9404 5188
rect 9398 5176 9404 5179
rect 9456 5176 9462 5228
rect 9858 5176 9864 5228
rect 9916 5216 9922 5228
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 9916 5188 12449 5216
rect 9916 5176 9922 5188
rect 12437 5185 12449 5188
rect 12483 5216 12495 5219
rect 13170 5216 13176 5228
rect 12483 5188 13176 5216
rect 12483 5185 12495 5188
rect 12437 5179 12495 5185
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 14918 5176 14924 5228
rect 14976 5216 14982 5228
rect 15028 5225 15056 5256
rect 17954 5244 17960 5256
rect 18012 5244 18018 5296
rect 18616 5284 18644 5315
rect 20438 5312 20444 5324
rect 20496 5312 20502 5364
rect 20530 5312 20536 5364
rect 20588 5352 20594 5364
rect 24673 5355 24731 5361
rect 24673 5352 24685 5355
rect 20588 5324 24685 5352
rect 20588 5312 20594 5324
rect 24673 5321 24685 5324
rect 24719 5321 24731 5355
rect 24673 5315 24731 5321
rect 28626 5312 28632 5364
rect 28684 5352 28690 5364
rect 28905 5355 28963 5361
rect 28905 5352 28917 5355
rect 28684 5324 28917 5352
rect 28684 5312 28690 5324
rect 28905 5321 28917 5324
rect 28951 5321 28963 5355
rect 31110 5352 31116 5364
rect 31071 5324 31116 5352
rect 28905 5315 28963 5321
rect 31110 5312 31116 5324
rect 31168 5312 31174 5364
rect 32674 5312 32680 5364
rect 32732 5352 32738 5364
rect 32769 5355 32827 5361
rect 32769 5352 32781 5355
rect 32732 5324 32781 5352
rect 32732 5312 32738 5324
rect 32769 5321 32781 5324
rect 32815 5321 32827 5355
rect 32769 5315 32827 5321
rect 35894 5312 35900 5364
rect 35952 5352 35958 5364
rect 35989 5355 36047 5361
rect 35989 5352 36001 5355
rect 35952 5324 36001 5352
rect 35952 5312 35958 5324
rect 35989 5321 36001 5324
rect 36035 5321 36047 5355
rect 35989 5315 36047 5321
rect 37274 5312 37280 5364
rect 37332 5352 37338 5364
rect 37645 5355 37703 5361
rect 37645 5352 37657 5355
rect 37332 5324 37657 5352
rect 37332 5312 37338 5324
rect 37645 5321 37657 5324
rect 37691 5321 37703 5355
rect 37645 5315 37703 5321
rect 19306 5287 19364 5293
rect 19306 5284 19318 5287
rect 18616 5256 19318 5284
rect 19306 5253 19318 5256
rect 19352 5253 19364 5287
rect 19306 5247 19364 5253
rect 19426 5244 19432 5296
rect 19484 5244 19490 5296
rect 24581 5287 24639 5293
rect 24581 5253 24593 5287
rect 24627 5284 24639 5287
rect 26326 5284 26332 5296
rect 24627 5256 26332 5284
rect 24627 5253 24639 5256
rect 24581 5247 24639 5253
rect 26326 5244 26332 5256
rect 26384 5244 26390 5296
rect 37660 5284 37688 5315
rect 40034 5312 40040 5364
rect 40092 5352 40098 5364
rect 40773 5355 40831 5361
rect 40773 5352 40785 5355
rect 40092 5324 40785 5352
rect 40092 5312 40098 5324
rect 40773 5321 40785 5324
rect 40819 5321 40831 5355
rect 40773 5315 40831 5321
rect 41141 5355 41199 5361
rect 41141 5321 41153 5355
rect 41187 5352 41199 5355
rect 41322 5352 41328 5364
rect 41187 5324 41328 5352
rect 41187 5321 41199 5324
rect 41141 5315 41199 5321
rect 41322 5312 41328 5324
rect 41380 5312 41386 5364
rect 48130 5312 48136 5364
rect 48188 5352 48194 5364
rect 48188 5324 51948 5352
rect 48188 5312 48194 5324
rect 41233 5287 41291 5293
rect 41233 5284 41245 5287
rect 37660 5256 41245 5284
rect 41233 5253 41245 5256
rect 41279 5284 41291 5287
rect 42426 5284 42432 5296
rect 41279 5256 42432 5284
rect 41279 5253 41291 5256
rect 41233 5247 41291 5253
rect 42426 5244 42432 5256
rect 42484 5244 42490 5296
rect 49510 5244 49516 5296
rect 49568 5284 49574 5296
rect 49568 5256 51856 5284
rect 49568 5244 49574 5256
rect 15013 5219 15071 5225
rect 15013 5216 15025 5219
rect 14976 5188 15025 5216
rect 14976 5176 14982 5188
rect 15013 5185 15025 5188
rect 15059 5185 15071 5219
rect 15746 5216 15752 5228
rect 15707 5188 15752 5216
rect 15013 5179 15071 5185
rect 15746 5176 15752 5188
rect 15804 5176 15810 5228
rect 18417 5219 18475 5225
rect 18417 5185 18429 5219
rect 18463 5216 18475 5219
rect 19444 5216 19472 5244
rect 18463 5188 19472 5216
rect 22465 5219 22523 5225
rect 18463 5185 18475 5188
rect 18417 5179 18475 5185
rect 22465 5185 22477 5219
rect 22511 5216 22523 5219
rect 22554 5216 22560 5228
rect 22511 5188 22560 5216
rect 22511 5185 22523 5188
rect 22465 5179 22523 5185
rect 22554 5176 22560 5188
rect 22612 5176 22618 5228
rect 23477 5219 23535 5225
rect 23477 5216 23489 5219
rect 22664 5188 23489 5216
rect 12066 5108 12072 5160
rect 12124 5148 12130 5160
rect 13354 5148 13360 5160
rect 12124 5120 13360 5148
rect 12124 5108 12130 5120
rect 13354 5108 13360 5120
rect 13412 5108 13418 5160
rect 14553 5151 14611 5157
rect 14553 5117 14565 5151
rect 14599 5148 14611 5151
rect 15930 5148 15936 5160
rect 14599 5120 15936 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 15930 5108 15936 5120
rect 15988 5108 15994 5160
rect 17862 5108 17868 5160
rect 17920 5148 17926 5160
rect 19061 5151 19119 5157
rect 19061 5148 19073 5151
rect 17920 5120 19073 5148
rect 17920 5108 17926 5120
rect 19061 5117 19073 5120
rect 19107 5117 19119 5151
rect 22664 5148 22692 5188
rect 23477 5185 23489 5188
rect 23523 5185 23535 5219
rect 25406 5216 25412 5228
rect 23477 5179 23535 5185
rect 24320 5188 25412 5216
rect 19061 5111 19119 5117
rect 22066 5120 22692 5148
rect 10410 5040 10416 5092
rect 10468 5080 10474 5092
rect 12434 5080 12440 5092
rect 10468 5052 12440 5080
rect 10468 5040 10474 5052
rect 12434 5040 12440 5052
rect 12492 5040 12498 5092
rect 13909 5083 13967 5089
rect 13909 5049 13921 5083
rect 13955 5080 13967 5083
rect 15010 5080 15016 5092
rect 13955 5052 15016 5080
rect 13955 5049 13967 5052
rect 13909 5043 13967 5049
rect 15010 5040 15016 5052
rect 15068 5040 15074 5092
rect 16022 5080 16028 5092
rect 15120 5052 16028 5080
rect 11977 5015 12035 5021
rect 11977 4981 11989 5015
rect 12023 5012 12035 5015
rect 12342 5012 12348 5024
rect 12023 4984 12348 5012
rect 12023 4981 12035 4984
rect 11977 4975 12035 4981
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 12618 5012 12624 5024
rect 12579 4984 12624 5012
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 13265 5015 13323 5021
rect 13265 4981 13277 5015
rect 13311 5012 13323 5015
rect 13814 5012 13820 5024
rect 13311 4984 13820 5012
rect 13311 4981 13323 4984
rect 13265 4975 13323 4981
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 15120 5021 15148 5052
rect 16022 5040 16028 5052
rect 16080 5040 16086 5092
rect 15105 5015 15163 5021
rect 15105 4981 15117 5015
rect 15151 4981 15163 5015
rect 15838 5012 15844 5024
rect 15799 4984 15844 5012
rect 15105 4975 15163 4981
rect 15838 4972 15844 4984
rect 15896 4972 15902 5024
rect 17313 5015 17371 5021
rect 17313 4981 17325 5015
rect 17359 5012 17371 5015
rect 17770 5012 17776 5024
rect 17359 4984 17776 5012
rect 17359 4981 17371 4984
rect 17313 4975 17371 4981
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 17957 5015 18015 5021
rect 17957 4981 17969 5015
rect 18003 5012 18015 5015
rect 18414 5012 18420 5024
rect 18003 4984 18420 5012
rect 18003 4981 18015 4984
rect 17957 4975 18015 4981
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 18598 4972 18604 5024
rect 18656 5012 18662 5024
rect 21913 5015 21971 5021
rect 21913 5012 21925 5015
rect 18656 4984 21925 5012
rect 18656 4972 18662 4984
rect 21913 4981 21925 4984
rect 21959 5012 21971 5015
rect 22066 5012 22094 5120
rect 23106 5108 23112 5160
rect 23164 5148 23170 5160
rect 23201 5151 23259 5157
rect 23201 5148 23213 5151
rect 23164 5120 23213 5148
rect 23164 5108 23170 5120
rect 23201 5117 23213 5120
rect 23247 5117 23259 5151
rect 23201 5111 23259 5117
rect 23385 5151 23443 5157
rect 23385 5117 23397 5151
rect 23431 5148 23443 5151
rect 24320 5148 24348 5188
rect 25406 5176 25412 5188
rect 25464 5216 25470 5228
rect 25774 5216 25780 5228
rect 25464 5188 25780 5216
rect 25464 5176 25470 5188
rect 25774 5176 25780 5188
rect 25832 5176 25838 5228
rect 27522 5216 27528 5228
rect 27483 5188 27528 5216
rect 27522 5176 27528 5188
rect 27580 5176 27586 5228
rect 27798 5225 27804 5228
rect 27792 5179 27804 5225
rect 27856 5216 27862 5228
rect 32861 5219 32919 5225
rect 27856 5188 27892 5216
rect 27798 5176 27804 5179
rect 27856 5176 27862 5188
rect 32861 5185 32873 5219
rect 32907 5216 32919 5219
rect 33778 5216 33784 5228
rect 32907 5188 33784 5216
rect 32907 5185 32919 5188
rect 32861 5179 32919 5185
rect 33778 5176 33784 5188
rect 33836 5176 33842 5228
rect 36173 5219 36231 5225
rect 36173 5185 36185 5219
rect 36219 5216 36231 5219
rect 37737 5219 37795 5225
rect 36219 5188 37320 5216
rect 36219 5185 36231 5188
rect 36173 5179 36231 5185
rect 23431 5120 24348 5148
rect 24397 5151 24455 5157
rect 23431 5117 23443 5120
rect 23385 5111 23443 5117
rect 24397 5117 24409 5151
rect 24443 5117 24455 5151
rect 24397 5111 24455 5117
rect 23216 5080 23244 5111
rect 24412 5080 24440 5111
rect 37292 5089 37320 5188
rect 37737 5185 37749 5219
rect 37783 5216 37795 5219
rect 38102 5216 38108 5228
rect 37783 5188 38108 5216
rect 37783 5185 37795 5188
rect 37737 5179 37795 5185
rect 38102 5176 38108 5188
rect 38160 5176 38166 5228
rect 38654 5216 38660 5228
rect 38615 5188 38660 5216
rect 38654 5176 38660 5188
rect 38712 5176 38718 5228
rect 38838 5176 38844 5228
rect 38896 5216 38902 5228
rect 39853 5219 39911 5225
rect 39853 5216 39865 5219
rect 38896 5188 39865 5216
rect 38896 5176 38902 5188
rect 39853 5185 39865 5188
rect 39899 5185 39911 5219
rect 39853 5179 39911 5185
rect 39942 5176 39948 5228
rect 40000 5216 40006 5228
rect 40000 5188 40045 5216
rect 40000 5176 40006 5188
rect 42794 5176 42800 5228
rect 42852 5216 42858 5228
rect 42889 5219 42947 5225
rect 42889 5216 42901 5219
rect 42852 5188 42901 5216
rect 42852 5176 42858 5188
rect 42889 5185 42901 5188
rect 42935 5216 42947 5219
rect 43441 5219 43499 5225
rect 43441 5216 43453 5219
rect 42935 5188 43453 5216
rect 42935 5185 42947 5188
rect 42889 5179 42947 5185
rect 43441 5185 43453 5188
rect 43487 5216 43499 5219
rect 49789 5219 49847 5225
rect 43487 5188 45324 5216
rect 43487 5185 43499 5188
rect 43441 5179 43499 5185
rect 37921 5151 37979 5157
rect 37921 5117 37933 5151
rect 37967 5148 37979 5151
rect 38378 5148 38384 5160
rect 37967 5120 38384 5148
rect 37967 5117 37979 5120
rect 37921 5111 37979 5117
rect 38378 5108 38384 5120
rect 38436 5148 38442 5160
rect 39761 5151 39819 5157
rect 38436 5120 39160 5148
rect 38436 5108 38442 5120
rect 23216 5052 24440 5080
rect 37277 5083 37335 5089
rect 37277 5049 37289 5083
rect 37323 5049 37335 5083
rect 37277 5043 37335 5049
rect 21959 4984 22094 5012
rect 22649 5015 22707 5021
rect 21959 4981 21971 4984
rect 21913 4975 21971 4981
rect 22649 4981 22661 5015
rect 22695 5012 22707 5015
rect 22738 5012 22744 5024
rect 22695 4984 22744 5012
rect 22695 4981 22707 4984
rect 22649 4975 22707 4981
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 23750 4972 23756 5024
rect 23808 5012 23814 5024
rect 23845 5015 23903 5021
rect 23845 5012 23857 5015
rect 23808 4984 23857 5012
rect 23808 4972 23814 4984
rect 23845 4981 23857 4984
rect 23891 4981 23903 5015
rect 23845 4975 23903 4981
rect 24578 4972 24584 5024
rect 24636 5012 24642 5024
rect 25041 5015 25099 5021
rect 25041 5012 25053 5015
rect 24636 4984 25053 5012
rect 24636 4972 24642 4984
rect 25041 4981 25053 4984
rect 25087 4981 25099 5015
rect 30650 5012 30656 5024
rect 30611 4984 30656 5012
rect 25041 4975 25099 4981
rect 30650 4972 30656 4984
rect 30708 4972 30714 5024
rect 37182 4972 37188 5024
rect 37240 5012 37246 5024
rect 38565 5015 38623 5021
rect 38565 5012 38577 5015
rect 37240 4984 38577 5012
rect 37240 4972 37246 4984
rect 38565 4981 38577 4984
rect 38611 4981 38623 5015
rect 39132 5012 39160 5120
rect 39761 5117 39773 5151
rect 39807 5117 39819 5151
rect 41322 5148 41328 5160
rect 39761 5111 39819 5117
rect 40144 5120 41328 5148
rect 39776 5080 39804 5111
rect 40144 5092 40172 5120
rect 41322 5108 41328 5120
rect 41380 5108 41386 5160
rect 43346 5108 43352 5160
rect 43404 5148 43410 5160
rect 45296 5157 45324 5188
rect 49789 5185 49801 5219
rect 49835 5216 49847 5219
rect 49878 5216 49884 5228
rect 49835 5188 49884 5216
rect 49835 5185 49847 5188
rect 49789 5179 49847 5185
rect 49878 5176 49884 5188
rect 49936 5176 49942 5228
rect 50062 5216 50068 5228
rect 50023 5188 50068 5216
rect 50062 5176 50068 5188
rect 50120 5176 50126 5228
rect 50614 5176 50620 5228
rect 50672 5216 50678 5228
rect 51828 5225 51856 5256
rect 51169 5219 51227 5225
rect 51169 5216 51181 5219
rect 50672 5188 51181 5216
rect 50672 5176 50678 5188
rect 51169 5185 51181 5188
rect 51215 5185 51227 5219
rect 51169 5179 51227 5185
rect 51813 5219 51871 5225
rect 51813 5185 51825 5219
rect 51859 5185 51871 5219
rect 51920 5216 51948 5324
rect 52733 5219 52791 5225
rect 52733 5216 52745 5219
rect 51920 5188 52745 5216
rect 51813 5179 51871 5185
rect 52733 5185 52745 5188
rect 52779 5216 52791 5219
rect 53377 5219 53435 5225
rect 53377 5216 53389 5219
rect 52779 5188 53389 5216
rect 52779 5185 52791 5188
rect 52733 5179 52791 5185
rect 53377 5185 53389 5188
rect 53423 5185 53435 5219
rect 53377 5179 53435 5185
rect 43901 5151 43959 5157
rect 43901 5148 43913 5151
rect 43404 5120 43913 5148
rect 43404 5108 43410 5120
rect 43901 5117 43913 5120
rect 43947 5117 43959 5151
rect 43901 5111 43959 5117
rect 45281 5151 45339 5157
rect 45281 5117 45293 5151
rect 45327 5148 45339 5151
rect 46290 5148 46296 5160
rect 45327 5120 46296 5148
rect 45327 5117 45339 5120
rect 45281 5111 45339 5117
rect 46290 5108 46296 5120
rect 46348 5108 46354 5160
rect 40126 5080 40132 5092
rect 39776 5052 40132 5080
rect 40126 5040 40132 5052
rect 40184 5040 40190 5092
rect 40310 5080 40316 5092
rect 40271 5052 40316 5080
rect 40310 5040 40316 5052
rect 40368 5040 40374 5092
rect 42613 5083 42671 5089
rect 42613 5049 42625 5083
rect 42659 5080 42671 5083
rect 46842 5080 46848 5092
rect 42659 5052 46848 5080
rect 42659 5049 42671 5052
rect 42613 5043 42671 5049
rect 46842 5040 46848 5052
rect 46900 5040 46906 5092
rect 47302 5040 47308 5092
rect 47360 5080 47366 5092
rect 48225 5083 48283 5089
rect 48225 5080 48237 5083
rect 47360 5052 48237 5080
rect 47360 5040 47366 5052
rect 48225 5049 48237 5052
rect 48271 5049 48283 5083
rect 48225 5043 48283 5049
rect 48682 5040 48688 5092
rect 48740 5080 48746 5092
rect 48740 5052 49188 5080
rect 48740 5040 48746 5052
rect 41782 5012 41788 5024
rect 39132 4984 41788 5012
rect 38565 4975 38623 4981
rect 41782 4972 41788 4984
rect 41840 5012 41846 5024
rect 42429 5015 42487 5021
rect 42429 5012 42441 5015
rect 41840 4984 42441 5012
rect 41840 4972 41846 4984
rect 42429 4981 42441 4984
rect 42475 4981 42487 5015
rect 42429 4975 42487 4981
rect 45646 4972 45652 5024
rect 45704 5012 45710 5024
rect 45741 5015 45799 5021
rect 45741 5012 45753 5015
rect 45704 4984 45753 5012
rect 45704 4972 45710 4984
rect 45741 4981 45753 4984
rect 45787 4981 45799 5015
rect 45741 4975 45799 4981
rect 45922 4972 45928 5024
rect 45980 5012 45986 5024
rect 46385 5015 46443 5021
rect 46385 5012 46397 5015
rect 45980 4984 46397 5012
rect 45980 4972 45986 4984
rect 46385 4981 46397 4984
rect 46431 4981 46443 5015
rect 46385 4975 46443 4981
rect 46750 4972 46756 5024
rect 46808 5012 46814 5024
rect 47581 5015 47639 5021
rect 47581 5012 47593 5015
rect 46808 4984 47593 5012
rect 46808 4972 46814 4984
rect 47581 4981 47593 4984
rect 47627 4981 47639 5015
rect 49050 5012 49056 5024
rect 49011 4984 49056 5012
rect 47581 4975 47639 4981
rect 49050 4972 49056 4984
rect 49108 4972 49114 5024
rect 49160 5012 49188 5052
rect 50525 5015 50583 5021
rect 50525 5012 50537 5015
rect 49160 4984 50537 5012
rect 50525 4981 50537 4984
rect 50571 4981 50583 5015
rect 50525 4975 50583 4981
rect 51353 5015 51411 5021
rect 51353 4981 51365 5015
rect 51399 5012 51411 5015
rect 51718 5012 51724 5024
rect 51399 4984 51724 5012
rect 51399 4981 51411 4984
rect 51353 4975 51411 4981
rect 51718 4972 51724 4984
rect 51776 4972 51782 5024
rect 52917 5015 52975 5021
rect 52917 4981 52929 5015
rect 52963 5012 52975 5015
rect 53282 5012 53288 5024
rect 52963 4984 53288 5012
rect 52963 4981 52975 4984
rect 52917 4975 52975 4981
rect 53282 4972 53288 4984
rect 53340 4972 53346 5024
rect 1104 4922 68816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 65654 4922
rect 65706 4870 65718 4922
rect 65770 4870 65782 4922
rect 65834 4870 65846 4922
rect 65898 4870 65910 4922
rect 65962 4870 68816 4922
rect 1104 4848 68816 4870
rect 9309 4811 9367 4817
rect 9309 4777 9321 4811
rect 9355 4808 9367 4811
rect 12710 4808 12716 4820
rect 9355 4780 12716 4808
rect 9355 4777 9367 4780
rect 9309 4771 9367 4777
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 14921 4811 14979 4817
rect 14921 4808 14933 4811
rect 14424 4780 14933 4808
rect 14424 4768 14430 4780
rect 14921 4777 14933 4780
rect 14967 4777 14979 4811
rect 14921 4771 14979 4777
rect 15654 4768 15660 4820
rect 15712 4808 15718 4820
rect 15841 4811 15899 4817
rect 15841 4808 15853 4811
rect 15712 4780 15853 4808
rect 15712 4768 15718 4780
rect 15841 4777 15853 4780
rect 15887 4777 15899 4811
rect 16025 4811 16083 4817
rect 16025 4808 16037 4811
rect 15841 4771 15899 4777
rect 15948 4780 16037 4808
rect 9858 4740 9864 4752
rect 9819 4712 9864 4740
rect 9858 4700 9864 4712
rect 9916 4700 9922 4752
rect 10410 4740 10416 4752
rect 10371 4712 10416 4740
rect 10410 4700 10416 4712
rect 10468 4700 10474 4752
rect 11609 4743 11667 4749
rect 11609 4709 11621 4743
rect 11655 4740 11667 4743
rect 14182 4740 14188 4752
rect 11655 4712 14188 4740
rect 11655 4709 11667 4712
rect 11609 4703 11667 4709
rect 14182 4700 14188 4712
rect 14240 4700 14246 4752
rect 14461 4743 14519 4749
rect 14461 4709 14473 4743
rect 14507 4740 14519 4743
rect 15746 4740 15752 4752
rect 14507 4712 15752 4740
rect 14507 4709 14519 4712
rect 14461 4703 14519 4709
rect 15746 4700 15752 4712
rect 15804 4700 15810 4752
rect 10965 4675 11023 4681
rect 10965 4641 10977 4675
rect 11011 4672 11023 4675
rect 13262 4672 13268 4684
rect 11011 4644 13268 4672
rect 11011 4641 11023 4644
rect 10965 4635 11023 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 13541 4675 13599 4681
rect 13541 4641 13553 4675
rect 13587 4672 13599 4675
rect 15654 4672 15660 4684
rect 13587 4644 15660 4672
rect 13587 4641 13599 4644
rect 13541 4635 13599 4641
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4604 8447 4607
rect 11422 4604 11428 4616
rect 8435 4576 11428 4604
rect 8435 4573 8447 4576
rect 8389 4567 8447 4573
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 12066 4604 12072 4616
rect 12027 4576 12072 4604
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 12710 4604 12716 4616
rect 12623 4576 12716 4604
rect 12710 4564 12716 4576
rect 12768 4604 12774 4616
rect 13446 4604 13452 4616
rect 12768 4576 13452 4604
rect 12768 4564 12774 4576
rect 13446 4564 13452 4576
rect 13504 4564 13510 4616
rect 14274 4604 14280 4616
rect 14235 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4573 14519 4607
rect 15948 4604 15976 4780
rect 16025 4777 16037 4780
rect 16071 4777 16083 4811
rect 16025 4771 16083 4777
rect 17037 4811 17095 4817
rect 17037 4777 17049 4811
rect 17083 4808 17095 4811
rect 17083 4780 20208 4808
rect 17083 4777 17095 4780
rect 17037 4771 17095 4777
rect 18049 4743 18107 4749
rect 18049 4709 18061 4743
rect 18095 4740 18107 4743
rect 18966 4740 18972 4752
rect 18095 4712 18972 4740
rect 18095 4709 18107 4712
rect 18049 4703 18107 4709
rect 18966 4700 18972 4712
rect 19024 4700 19030 4752
rect 20180 4740 20208 4780
rect 20254 4768 20260 4820
rect 20312 4808 20318 4820
rect 20625 4811 20683 4817
rect 20625 4808 20637 4811
rect 20312 4780 20637 4808
rect 20312 4768 20318 4780
rect 20625 4777 20637 4780
rect 20671 4777 20683 4811
rect 20625 4771 20683 4777
rect 23845 4811 23903 4817
rect 23845 4777 23857 4811
rect 23891 4808 23903 4811
rect 24118 4808 24124 4820
rect 23891 4780 24124 4808
rect 23891 4777 23903 4780
rect 23845 4771 23903 4777
rect 24118 4768 24124 4780
rect 24176 4768 24182 4820
rect 27709 4811 27767 4817
rect 27709 4777 27721 4811
rect 27755 4808 27767 4811
rect 27798 4808 27804 4820
rect 27755 4780 27804 4808
rect 27755 4777 27767 4780
rect 27709 4771 27767 4777
rect 27798 4768 27804 4780
rect 27856 4768 27862 4820
rect 40218 4768 40224 4820
rect 40276 4808 40282 4820
rect 40405 4811 40463 4817
rect 40405 4808 40417 4811
rect 40276 4780 40417 4808
rect 40276 4768 40282 4780
rect 40405 4777 40417 4780
rect 40451 4777 40463 4811
rect 40405 4771 40463 4777
rect 40954 4768 40960 4820
rect 41012 4808 41018 4820
rect 41601 4811 41659 4817
rect 41601 4808 41613 4811
rect 41012 4780 41613 4808
rect 41012 4768 41018 4780
rect 41601 4777 41613 4780
rect 41647 4777 41659 4811
rect 41601 4771 41659 4777
rect 48130 4768 48136 4820
rect 48188 4808 48194 4820
rect 50801 4811 50859 4817
rect 50801 4808 50813 4811
rect 48188 4780 50813 4808
rect 48188 4768 48194 4780
rect 50801 4777 50813 4780
rect 50847 4777 50859 4811
rect 54018 4808 54024 4820
rect 53979 4780 54024 4808
rect 50801 4771 50859 4777
rect 54018 4768 54024 4780
rect 54076 4768 54082 4820
rect 54570 4808 54576 4820
rect 54531 4780 54576 4808
rect 54570 4768 54576 4780
rect 54628 4768 54634 4820
rect 55306 4808 55312 4820
rect 55267 4780 55312 4808
rect 55306 4768 55312 4780
rect 55364 4768 55370 4820
rect 22002 4740 22008 4752
rect 20180 4712 22008 4740
rect 22002 4700 22008 4712
rect 22060 4700 22066 4752
rect 37553 4743 37611 4749
rect 37553 4709 37565 4743
rect 37599 4740 37611 4743
rect 38102 4740 38108 4752
rect 37599 4712 38108 4740
rect 37599 4709 37611 4712
rect 37553 4703 37611 4709
rect 38102 4700 38108 4712
rect 38160 4740 38166 4752
rect 41230 4740 41236 4752
rect 38160 4712 41236 4740
rect 38160 4700 38166 4712
rect 41230 4700 41236 4712
rect 41288 4700 41294 4752
rect 47210 4700 47216 4752
rect 47268 4740 47274 4752
rect 48869 4743 48927 4749
rect 48869 4740 48881 4743
rect 47268 4712 48881 4740
rect 47268 4700 47274 4712
rect 48869 4709 48881 4712
rect 48915 4709 48927 4743
rect 48869 4703 48927 4709
rect 49970 4700 49976 4752
rect 50028 4740 50034 4752
rect 52733 4743 52791 4749
rect 52733 4740 52745 4743
rect 50028 4712 52745 4740
rect 50028 4700 50034 4712
rect 52733 4709 52745 4712
rect 52779 4709 52791 4743
rect 52733 4703 52791 4709
rect 16022 4632 16028 4684
rect 16080 4672 16086 4684
rect 16117 4675 16175 4681
rect 16117 4672 16129 4675
rect 16080 4644 16129 4672
rect 16080 4632 16086 4644
rect 16117 4641 16129 4644
rect 16163 4672 16175 4675
rect 16666 4672 16672 4684
rect 16163 4644 16672 4672
rect 16163 4641 16175 4644
rect 16117 4635 16175 4641
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 17862 4632 17868 4684
rect 17920 4672 17926 4684
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 17920 4644 19257 4672
rect 17920 4632 17926 4644
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 22462 4672 22468 4684
rect 22423 4644 22468 4672
rect 19245 4635 19303 4641
rect 22462 4632 22468 4644
rect 22520 4632 22526 4684
rect 38381 4675 38439 4681
rect 38381 4641 38393 4675
rect 38427 4672 38439 4675
rect 38930 4672 38936 4684
rect 38427 4644 38936 4672
rect 38427 4641 38439 4644
rect 38381 4635 38439 4641
rect 38930 4632 38936 4644
rect 38988 4632 38994 4684
rect 41049 4675 41107 4681
rect 41049 4641 41061 4675
rect 41095 4672 41107 4675
rect 41138 4672 41144 4684
rect 41095 4644 41144 4672
rect 41095 4641 41107 4644
rect 41049 4635 41107 4641
rect 41138 4632 41144 4644
rect 41196 4632 41202 4684
rect 41322 4632 41328 4684
rect 41380 4672 41386 4684
rect 42153 4675 42211 4681
rect 42153 4672 42165 4675
rect 41380 4644 42165 4672
rect 41380 4632 41386 4644
rect 42153 4641 42165 4644
rect 42199 4641 42211 4675
rect 42153 4635 42211 4641
rect 44818 4632 44824 4684
rect 44876 4672 44882 4684
rect 45649 4675 45707 4681
rect 45649 4672 45661 4675
rect 44876 4644 45661 4672
rect 44876 4632 44882 4644
rect 45649 4641 45661 4644
rect 45695 4641 45707 4675
rect 45649 4635 45707 4641
rect 46198 4632 46204 4684
rect 46256 4672 46262 4684
rect 47581 4675 47639 4681
rect 47581 4672 47593 4675
rect 46256 4644 47593 4672
rect 46256 4632 46262 4644
rect 47581 4641 47593 4644
rect 47627 4641 47639 4675
rect 47581 4635 47639 4641
rect 47670 4632 47676 4684
rect 47728 4672 47734 4684
rect 50157 4675 50215 4681
rect 50157 4672 50169 4675
rect 47728 4644 50169 4672
rect 47728 4632 47734 4644
rect 50157 4641 50169 4644
rect 50203 4641 50215 4675
rect 50157 4635 50215 4641
rect 51166 4632 51172 4684
rect 51224 4672 51230 4684
rect 53377 4675 53435 4681
rect 53377 4672 53389 4675
rect 51224 4644 53389 4672
rect 51224 4632 51230 4644
rect 53377 4641 53389 4644
rect 53423 4641 53435 4675
rect 53377 4635 53435 4641
rect 16206 4604 16212 4616
rect 14461 4567 14519 4573
rect 15120 4576 15976 4604
rect 16167 4576 16212 4604
rect 11606 4496 11612 4548
rect 11664 4536 11670 4548
rect 14476 4536 14504 4567
rect 15120 4548 15148 4576
rect 16206 4564 16212 4576
rect 16264 4564 16270 4616
rect 16850 4604 16856 4616
rect 16592 4576 16856 4604
rect 14826 4536 14832 4548
rect 11664 4508 14832 4536
rect 11664 4496 11670 4508
rect 14826 4496 14832 4508
rect 14884 4496 14890 4548
rect 15102 4536 15108 4548
rect 15063 4508 15108 4536
rect 15102 4496 15108 4508
rect 15160 4496 15166 4548
rect 15289 4539 15347 4545
rect 15289 4505 15301 4539
rect 15335 4536 15347 4539
rect 16592 4536 16620 4576
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 18693 4607 18751 4613
rect 18693 4573 18705 4607
rect 18739 4604 18751 4607
rect 18739 4576 19288 4604
rect 18739 4573 18751 4576
rect 18693 4567 18751 4573
rect 19260 4548 19288 4576
rect 19334 4564 19340 4616
rect 19392 4604 19398 4616
rect 19501 4607 19559 4613
rect 19501 4604 19513 4607
rect 19392 4576 19513 4604
rect 19392 4564 19398 4576
rect 19501 4573 19513 4576
rect 19547 4573 19559 4607
rect 19501 4567 19559 4573
rect 21082 4564 21088 4616
rect 21140 4604 21146 4616
rect 22738 4613 22744 4616
rect 21269 4607 21327 4613
rect 21269 4604 21281 4607
rect 21140 4576 21281 4604
rect 21140 4564 21146 4576
rect 21269 4573 21281 4576
rect 21315 4604 21327 4607
rect 21729 4607 21787 4613
rect 21729 4604 21741 4607
rect 21315 4576 21741 4604
rect 21315 4573 21327 4576
rect 21269 4567 21327 4573
rect 21729 4573 21741 4576
rect 21775 4573 21787 4607
rect 22732 4604 22744 4613
rect 22699 4576 22744 4604
rect 21729 4567 21787 4573
rect 22732 4567 22744 4576
rect 22738 4564 22744 4567
rect 22796 4564 22802 4616
rect 24578 4604 24584 4616
rect 24539 4576 24584 4604
rect 24578 4564 24584 4576
rect 24636 4564 24642 4616
rect 27525 4607 27583 4613
rect 27525 4573 27537 4607
rect 27571 4604 27583 4607
rect 27982 4604 27988 4616
rect 27571 4576 27988 4604
rect 27571 4573 27583 4576
rect 27525 4567 27583 4573
rect 27982 4564 27988 4576
rect 28040 4564 28046 4616
rect 29914 4564 29920 4616
rect 29972 4604 29978 4616
rect 30009 4607 30067 4613
rect 30009 4604 30021 4607
rect 29972 4576 30021 4604
rect 29972 4564 29978 4576
rect 30009 4573 30021 4576
rect 30055 4573 30067 4607
rect 31110 4604 31116 4616
rect 31071 4576 31116 4604
rect 30009 4567 30067 4573
rect 31110 4564 31116 4576
rect 31168 4564 31174 4616
rect 31846 4564 31852 4616
rect 31904 4604 31910 4616
rect 31941 4607 31999 4613
rect 31941 4604 31953 4607
rect 31904 4576 31953 4604
rect 31904 4564 31910 4576
rect 31941 4573 31953 4576
rect 31987 4573 31999 4607
rect 35802 4604 35808 4616
rect 35763 4576 35808 4604
rect 31941 4567 31999 4573
rect 35802 4564 35808 4576
rect 35860 4564 35866 4616
rect 37182 4564 37188 4616
rect 37240 4564 37246 4616
rect 38746 4564 38752 4616
rect 38804 4604 38810 4616
rect 38841 4607 38899 4613
rect 38841 4604 38853 4607
rect 38804 4576 38853 4604
rect 38804 4564 38810 4576
rect 38841 4573 38853 4576
rect 38887 4573 38899 4607
rect 42794 4604 42800 4616
rect 38841 4567 38899 4573
rect 38948 4576 42800 4604
rect 15335 4508 16620 4536
rect 16669 4539 16727 4545
rect 15335 4505 15347 4508
rect 15289 4499 15347 4505
rect 16669 4505 16681 4539
rect 16715 4536 16727 4539
rect 16942 4536 16948 4548
rect 16715 4508 16948 4536
rect 16715 4505 16727 4508
rect 16669 4499 16727 4505
rect 16942 4496 16948 4508
rect 17000 4496 17006 4548
rect 19242 4496 19248 4548
rect 19300 4496 19306 4548
rect 36078 4536 36084 4548
rect 36039 4508 36084 4536
rect 36078 4496 36084 4508
rect 36136 4496 36142 4548
rect 12250 4468 12256 4480
rect 12211 4440 12256 4468
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 12897 4471 12955 4477
rect 12897 4437 12909 4471
rect 12943 4468 12955 4471
rect 15470 4468 15476 4480
rect 12943 4440 15476 4468
rect 12943 4437 12955 4440
rect 12897 4431 12955 4437
rect 15470 4428 15476 4440
rect 15528 4428 15534 4480
rect 20990 4428 20996 4480
rect 21048 4468 21054 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 21048 4440 21097 4468
rect 21048 4428 21054 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 24765 4471 24823 4477
rect 24765 4437 24777 4471
rect 24811 4468 24823 4471
rect 24946 4468 24952 4480
rect 24811 4440 24952 4468
rect 24811 4437 24823 4440
rect 24765 4431 24823 4437
rect 24946 4428 24952 4440
rect 25004 4428 25010 4480
rect 32950 4428 32956 4480
rect 33008 4468 33014 4480
rect 33597 4471 33655 4477
rect 33597 4468 33609 4471
rect 33008 4440 33609 4468
rect 33008 4428 33014 4440
rect 33597 4437 33609 4440
rect 33643 4468 33655 4471
rect 38948 4468 38976 4576
rect 42794 4564 42800 4576
rect 42852 4564 42858 4616
rect 42978 4604 42984 4616
rect 42939 4576 42984 4604
rect 42978 4564 42984 4576
rect 43036 4564 43042 4616
rect 43346 4564 43352 4616
rect 43404 4604 43410 4616
rect 43441 4607 43499 4613
rect 43441 4604 43453 4607
rect 43404 4576 43453 4604
rect 43404 4564 43410 4576
rect 43441 4573 43453 4576
rect 43487 4573 43499 4607
rect 44266 4604 44272 4616
rect 44227 4576 44272 4604
rect 43441 4567 43499 4573
rect 44266 4564 44272 4576
rect 44324 4564 44330 4616
rect 45094 4564 45100 4616
rect 45152 4604 45158 4616
rect 45189 4607 45247 4613
rect 45189 4604 45201 4607
rect 45152 4576 45201 4604
rect 45152 4564 45158 4576
rect 45189 4573 45201 4576
rect 45235 4573 45247 4607
rect 45189 4567 45247 4573
rect 45370 4564 45376 4616
rect 45428 4604 45434 4616
rect 46293 4607 46351 4613
rect 46293 4604 46305 4607
rect 45428 4576 46305 4604
rect 45428 4564 45434 4576
rect 46293 4573 46305 4576
rect 46339 4573 46351 4607
rect 46934 4604 46940 4616
rect 46895 4576 46940 4604
rect 46293 4567 46351 4573
rect 46934 4564 46940 4576
rect 46992 4564 46998 4616
rect 48038 4564 48044 4616
rect 48096 4604 48102 4616
rect 48225 4607 48283 4613
rect 48225 4604 48237 4607
rect 48096 4576 48237 4604
rect 48096 4564 48102 4576
rect 48225 4573 48237 4576
rect 48271 4573 48283 4607
rect 48225 4567 48283 4573
rect 48314 4564 48320 4616
rect 48372 4604 48378 4616
rect 49513 4607 49571 4613
rect 49513 4604 49525 4607
rect 48372 4576 49525 4604
rect 48372 4564 48378 4576
rect 49513 4573 49525 4576
rect 49559 4573 49571 4607
rect 49513 4567 49571 4573
rect 50890 4564 50896 4616
rect 50948 4604 50954 4616
rect 51445 4607 51503 4613
rect 51445 4604 51457 4607
rect 50948 4576 51457 4604
rect 50948 4564 50954 4576
rect 51445 4573 51457 4576
rect 51491 4573 51503 4607
rect 51445 4567 51503 4573
rect 52273 4607 52331 4613
rect 52273 4573 52285 4607
rect 52319 4573 52331 4607
rect 52273 4567 52331 4573
rect 40862 4536 40868 4548
rect 40823 4508 40868 4536
rect 40862 4496 40868 4508
rect 40920 4496 40926 4548
rect 41969 4539 42027 4545
rect 41969 4505 41981 4539
rect 42015 4536 42027 4539
rect 42518 4536 42524 4548
rect 42015 4508 42524 4536
rect 42015 4505 42027 4508
rect 41969 4499 42027 4505
rect 42518 4496 42524 4508
rect 42576 4496 42582 4548
rect 42610 4496 42616 4548
rect 42668 4536 42674 4548
rect 42668 4508 49648 4536
rect 42668 4496 42674 4508
rect 39850 4468 39856 4480
rect 33643 4440 38976 4468
rect 39811 4440 39856 4468
rect 33643 4437 33655 4440
rect 33597 4431 33655 4437
rect 39850 4428 39856 4440
rect 39908 4468 39914 4480
rect 40773 4471 40831 4477
rect 40773 4468 40785 4471
rect 39908 4440 40785 4468
rect 39908 4428 39914 4440
rect 40773 4437 40785 4440
rect 40819 4437 40831 4471
rect 40773 4431 40831 4437
rect 42061 4471 42119 4477
rect 42061 4437 42073 4471
rect 42107 4468 42119 4471
rect 42334 4468 42340 4480
rect 42107 4440 42340 4468
rect 42107 4437 42119 4440
rect 42061 4431 42119 4437
rect 42334 4428 42340 4440
rect 42392 4428 42398 4480
rect 42794 4468 42800 4480
rect 42755 4440 42800 4468
rect 42794 4428 42800 4440
rect 42852 4428 42858 4480
rect 43530 4468 43536 4480
rect 43491 4440 43536 4468
rect 43530 4428 43536 4440
rect 43588 4428 43594 4480
rect 44174 4468 44180 4480
rect 44135 4440 44180 4468
rect 44174 4428 44180 4440
rect 44232 4428 44238 4480
rect 45002 4468 45008 4480
rect 44963 4440 45008 4468
rect 45002 4428 45008 4440
rect 45060 4428 45066 4480
rect 47026 4428 47032 4480
rect 47084 4468 47090 4480
rect 47121 4471 47179 4477
rect 47121 4468 47133 4471
rect 47084 4440 47133 4468
rect 47084 4428 47090 4440
rect 47121 4437 47133 4440
rect 47167 4437 47179 4471
rect 48406 4468 48412 4480
rect 48367 4440 48412 4468
rect 47121 4431 47179 4437
rect 48406 4428 48412 4440
rect 48464 4428 48470 4480
rect 49620 4468 49648 4508
rect 50706 4496 50712 4548
rect 50764 4536 50770 4548
rect 52288 4536 52316 4567
rect 50764 4508 52316 4536
rect 50764 4496 50770 4508
rect 51626 4468 51632 4480
rect 49620 4440 51632 4468
rect 51626 4428 51632 4440
rect 51684 4428 51690 4480
rect 52086 4468 52092 4480
rect 52047 4440 52092 4468
rect 52086 4428 52092 4440
rect 52144 4428 52150 4480
rect 55950 4468 55956 4480
rect 55911 4440 55956 4468
rect 55950 4428 55956 4440
rect 56008 4428 56014 4480
rect 1104 4378 68816 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 68816 4378
rect 1104 4304 68816 4326
rect 9217 4267 9275 4273
rect 9217 4233 9229 4267
rect 9263 4264 9275 4267
rect 12066 4264 12072 4276
rect 9263 4236 12072 4264
rect 9263 4233 9275 4236
rect 9217 4227 9275 4233
rect 12066 4224 12072 4236
rect 12124 4224 12130 4276
rect 12713 4267 12771 4273
rect 12406 4236 12664 4264
rect 8662 4128 8668 4140
rect 8623 4100 8668 4128
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4128 9827 4131
rect 12406 4128 12434 4236
rect 12636 4196 12664 4236
rect 12713 4233 12725 4267
rect 12759 4264 12771 4267
rect 14274 4264 14280 4276
rect 12759 4236 14280 4264
rect 12759 4233 12771 4236
rect 12713 4227 12771 4233
rect 14274 4224 14280 4236
rect 14332 4224 14338 4276
rect 15838 4264 15844 4276
rect 15799 4236 15844 4264
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 16850 4224 16856 4276
rect 16908 4264 16914 4276
rect 17773 4267 17831 4273
rect 17773 4264 17785 4267
rect 16908 4236 17785 4264
rect 16908 4224 16914 4236
rect 17773 4233 17785 4236
rect 17819 4233 17831 4267
rect 17773 4227 17831 4233
rect 19521 4267 19579 4273
rect 19521 4233 19533 4267
rect 19567 4264 19579 4267
rect 20254 4264 20260 4276
rect 19567 4236 20260 4264
rect 19567 4233 19579 4236
rect 19521 4227 19579 4233
rect 20254 4224 20260 4236
rect 20312 4224 20318 4276
rect 26053 4267 26111 4273
rect 26053 4233 26065 4267
rect 26099 4264 26111 4267
rect 26326 4264 26332 4276
rect 26099 4236 26332 4264
rect 26099 4233 26111 4236
rect 26053 4227 26111 4233
rect 26326 4224 26332 4236
rect 26384 4224 26390 4276
rect 33042 4264 33048 4276
rect 33003 4236 33048 4264
rect 33042 4224 33048 4236
rect 33100 4224 33106 4276
rect 36078 4224 36084 4276
rect 36136 4264 36142 4276
rect 36541 4267 36599 4273
rect 36541 4264 36553 4267
rect 36136 4236 36553 4264
rect 36136 4224 36142 4236
rect 36541 4233 36553 4236
rect 36587 4233 36599 4267
rect 36541 4227 36599 4233
rect 41601 4267 41659 4273
rect 41601 4233 41613 4267
rect 41647 4264 41659 4267
rect 42610 4264 42616 4276
rect 41647 4236 42616 4264
rect 41647 4233 41659 4236
rect 41601 4227 41659 4233
rect 42610 4224 42616 4236
rect 42668 4224 42674 4276
rect 46382 4264 46388 4276
rect 46343 4236 46388 4264
rect 46382 4224 46388 4236
rect 46440 4224 46446 4276
rect 48406 4224 48412 4276
rect 48464 4264 48470 4276
rect 49510 4264 49516 4276
rect 48464 4236 49516 4264
rect 48464 4224 48470 4236
rect 49510 4224 49516 4236
rect 49568 4224 49574 4276
rect 49697 4267 49755 4273
rect 49697 4233 49709 4267
rect 49743 4264 49755 4267
rect 50890 4264 50896 4276
rect 49743 4236 50896 4264
rect 49743 4233 49755 4236
rect 49697 4227 49755 4233
rect 50890 4224 50896 4236
rect 50948 4224 50954 4276
rect 54018 4224 54024 4276
rect 54076 4264 54082 4276
rect 67174 4264 67180 4276
rect 54076 4236 67180 4264
rect 54076 4224 54082 4236
rect 67174 4224 67180 4236
rect 67232 4224 67238 4276
rect 13722 4196 13728 4208
rect 12636 4168 13728 4196
rect 13722 4156 13728 4168
rect 13780 4196 13786 4208
rect 13909 4199 13967 4205
rect 13909 4196 13921 4199
rect 13780 4168 13921 4196
rect 13780 4156 13786 4168
rect 13909 4165 13921 4168
rect 13955 4165 13967 4199
rect 14642 4196 14648 4208
rect 14603 4168 14648 4196
rect 13909 4159 13967 4165
rect 14642 4156 14648 4168
rect 14700 4156 14706 4208
rect 15378 4156 15384 4208
rect 15436 4196 15442 4208
rect 15657 4199 15715 4205
rect 15657 4196 15669 4199
rect 15436 4168 15669 4196
rect 15436 4156 15442 4168
rect 15657 4165 15669 4168
rect 15703 4196 15715 4199
rect 15703 4168 16160 4196
rect 15703 4165 15715 4168
rect 15657 4159 15715 4165
rect 9815 4100 12434 4128
rect 12529 4131 12587 4137
rect 9815 4097 9827 4100
rect 9769 4091 9827 4097
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 12802 4128 12808 4140
rect 12575 4100 12808 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 12802 4088 12808 4100
rect 12860 4128 12866 4140
rect 13538 4128 13544 4140
rect 12860 4100 13544 4128
rect 12860 4088 12866 4100
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4128 14151 4131
rect 15286 4128 15292 4140
rect 14139 4100 15292 4128
rect 14139 4097 14151 4100
rect 14093 4091 14151 4097
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 15470 4128 15476 4140
rect 15431 4100 15476 4128
rect 15470 4088 15476 4100
rect 15528 4088 15534 4140
rect 15746 4128 15752 4140
rect 15707 4100 15752 4128
rect 15746 4088 15752 4100
rect 15804 4088 15810 4140
rect 16132 4128 16160 4168
rect 16206 4156 16212 4208
rect 16264 4196 16270 4208
rect 17313 4199 17371 4205
rect 16264 4168 17080 4196
rect 16264 4156 16270 4168
rect 16482 4128 16488 4140
rect 16132 4100 16488 4128
rect 16482 4088 16488 4100
rect 16540 4088 16546 4140
rect 16666 4128 16672 4140
rect 16627 4100 16672 4128
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 17052 4137 17080 4168
rect 17313 4165 17325 4199
rect 17359 4196 17371 4199
rect 25038 4196 25044 4208
rect 17359 4168 25044 4196
rect 17359 4165 17371 4168
rect 17313 4159 17371 4165
rect 25038 4156 25044 4168
rect 25096 4156 25102 4208
rect 30208 4168 30420 4196
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17083 4100 17908 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 12069 4063 12127 4069
rect 12069 4029 12081 4063
rect 12115 4060 12127 4063
rect 13357 4063 13415 4069
rect 12115 4032 13216 4060
rect 12115 4029 12127 4032
rect 12069 4023 12127 4029
rect 10965 3995 11023 4001
rect 10965 3961 10977 3995
rect 11011 3992 11023 3995
rect 12802 3992 12808 4004
rect 11011 3964 12808 3992
rect 11011 3961 11023 3964
rect 10965 3955 11023 3961
rect 12802 3952 12808 3964
rect 12860 3952 12866 4004
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 13188 3924 13216 4032
rect 13357 4029 13369 4063
rect 13403 4060 13415 4063
rect 16850 4060 16856 4072
rect 13403 4032 16856 4060
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 17129 4063 17187 4069
rect 17129 4029 17141 4063
rect 17175 4029 17187 4063
rect 17880 4060 17908 4100
rect 17954 4088 17960 4140
rect 18012 4128 18018 4140
rect 18141 4131 18199 4137
rect 18012 4100 18057 4128
rect 18012 4088 18018 4100
rect 18141 4097 18153 4131
rect 18187 4128 18199 4131
rect 18230 4128 18236 4140
rect 18187 4100 18236 4128
rect 18187 4097 18199 4100
rect 18141 4091 18199 4097
rect 18156 4060 18184 4091
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 18598 4128 18604 4140
rect 18559 4100 18604 4128
rect 18598 4088 18604 4100
rect 18656 4128 18662 4140
rect 19613 4131 19671 4137
rect 19613 4128 19625 4131
rect 18656 4100 19625 4128
rect 18656 4088 18662 4100
rect 19613 4097 19625 4100
rect 19659 4097 19671 4131
rect 19613 4091 19671 4097
rect 19978 4088 19984 4140
rect 20036 4128 20042 4140
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 20036 4100 20821 4128
rect 20036 4088 20042 4100
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 20990 4128 20996 4140
rect 20951 4100 20996 4128
rect 20809 4091 20867 4097
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 23750 4128 23756 4140
rect 23711 4100 23756 4128
rect 23750 4088 23756 4100
rect 23808 4088 23814 4140
rect 24946 4137 24952 4140
rect 24940 4128 24952 4137
rect 24907 4100 24952 4128
rect 24940 4091 24952 4100
rect 24946 4088 24952 4091
rect 25004 4088 25010 4140
rect 29457 4131 29515 4137
rect 29457 4097 29469 4131
rect 29503 4128 29515 4131
rect 30208 4128 30236 4168
rect 29503 4100 30236 4128
rect 30285 4131 30343 4137
rect 29503 4097 29515 4100
rect 29457 4091 29515 4097
rect 30285 4097 30297 4131
rect 30331 4097 30343 4131
rect 30392 4128 30420 4168
rect 38838 4156 38844 4208
rect 38896 4196 38902 4208
rect 41509 4199 41567 4205
rect 41509 4196 41521 4199
rect 38896 4168 41521 4196
rect 38896 4156 38902 4168
rect 41509 4165 41521 4168
rect 41555 4196 41567 4199
rect 42242 4196 42248 4208
rect 41555 4168 42248 4196
rect 41555 4165 41567 4168
rect 41509 4159 41567 4165
rect 42242 4156 42248 4168
rect 42300 4156 42306 4208
rect 44174 4156 44180 4208
rect 44232 4156 44238 4208
rect 44913 4199 44971 4205
rect 44913 4165 44925 4199
rect 44959 4196 44971 4199
rect 45002 4196 45008 4208
rect 44959 4168 45008 4196
rect 44959 4165 44971 4168
rect 44913 4159 44971 4165
rect 45002 4156 45008 4168
rect 45060 4156 45066 4208
rect 30837 4131 30895 4137
rect 30837 4128 30849 4131
rect 30392 4100 30849 4128
rect 30285 4091 30343 4097
rect 30837 4097 30849 4100
rect 30883 4128 30895 4131
rect 31297 4131 31355 4137
rect 31297 4128 31309 4131
rect 30883 4100 31309 4128
rect 30883 4097 30895 4100
rect 30837 4091 30895 4097
rect 31297 4097 31309 4100
rect 31343 4128 31355 4131
rect 31754 4128 31760 4140
rect 31343 4100 31760 4128
rect 31343 4097 31355 4100
rect 31297 4091 31355 4097
rect 17880 4032 18184 4060
rect 19797 4063 19855 4069
rect 17129 4023 17187 4029
rect 19797 4029 19809 4063
rect 19843 4060 19855 4063
rect 19886 4060 19892 4072
rect 19843 4032 19892 4060
rect 19843 4029 19855 4032
rect 19797 4023 19855 4029
rect 13446 3952 13452 4004
rect 13504 3992 13510 4004
rect 14366 3992 14372 4004
rect 13504 3964 14372 3992
rect 13504 3952 13510 3964
rect 14366 3952 14372 3964
rect 14424 3952 14430 4004
rect 14918 3952 14924 4004
rect 14976 3992 14982 4004
rect 16942 3992 16948 4004
rect 14976 3964 16948 3992
rect 14976 3952 14982 3964
rect 16942 3952 16948 3964
rect 17000 3992 17006 4004
rect 17144 3992 17172 4023
rect 19886 4020 19892 4032
rect 19944 4020 19950 4072
rect 24673 4063 24731 4069
rect 24673 4029 24685 4063
rect 24719 4029 24731 4063
rect 30300 4060 30328 4091
rect 31754 4088 31760 4100
rect 31812 4128 31818 4140
rect 32217 4131 32275 4137
rect 32217 4128 32229 4131
rect 31812 4100 32229 4128
rect 31812 4088 31818 4100
rect 32217 4097 32229 4100
rect 32263 4097 32275 4131
rect 32217 4091 32275 4097
rect 33137 4131 33195 4137
rect 33137 4097 33149 4131
rect 33183 4128 33195 4131
rect 33873 4131 33931 4137
rect 33873 4128 33885 4131
rect 33183 4100 33885 4128
rect 33183 4097 33195 4100
rect 33137 4091 33195 4097
rect 33873 4097 33885 4100
rect 33919 4097 33931 4131
rect 33873 4091 33931 4097
rect 36725 4131 36783 4137
rect 36725 4097 36737 4131
rect 36771 4128 36783 4131
rect 37366 4128 37372 4140
rect 36771 4100 37372 4128
rect 36771 4097 36783 4100
rect 36725 4091 36783 4097
rect 32122 4060 32128 4072
rect 30300 4032 32128 4060
rect 24673 4023 24731 4029
rect 19150 3992 19156 4004
rect 17000 3964 17172 3992
rect 19111 3964 19156 3992
rect 17000 3952 17006 3964
rect 19150 3952 19156 3964
rect 19208 3952 19214 4004
rect 14550 3924 14556 3936
rect 13188 3896 14556 3924
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14734 3924 14740 3936
rect 14695 3896 14740 3924
rect 14734 3884 14740 3896
rect 14792 3884 14798 3936
rect 14826 3884 14832 3936
rect 14884 3924 14890 3936
rect 15562 3924 15568 3936
rect 14884 3896 15568 3924
rect 14884 3884 14890 3896
rect 15562 3884 15568 3896
rect 15620 3924 15626 3936
rect 15746 3924 15752 3936
rect 15620 3896 15752 3924
rect 15620 3884 15626 3896
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 16025 3927 16083 3933
rect 16025 3893 16037 3927
rect 16071 3924 16083 3927
rect 16758 3924 16764 3936
rect 16071 3896 16764 3924
rect 16071 3893 16083 3896
rect 16025 3887 16083 3893
rect 16758 3884 16764 3896
rect 16816 3884 16822 3936
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 20901 3927 20959 3933
rect 20901 3924 20913 3927
rect 20588 3896 20913 3924
rect 20588 3884 20594 3896
rect 20901 3893 20913 3896
rect 20947 3893 20959 3927
rect 20901 3887 20959 3893
rect 21726 3884 21732 3936
rect 21784 3924 21790 3936
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 21784 3896 21833 3924
rect 21784 3884 21790 3896
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 21821 3887 21879 3893
rect 23014 3884 23020 3936
rect 23072 3924 23078 3936
rect 23109 3927 23167 3933
rect 23109 3924 23121 3927
rect 23072 3896 23121 3924
rect 23072 3884 23078 3896
rect 23109 3893 23121 3896
rect 23155 3893 23167 3927
rect 23934 3924 23940 3936
rect 23895 3896 23940 3924
rect 23109 3887 23167 3893
rect 23934 3884 23940 3896
rect 23992 3884 23998 3936
rect 24394 3884 24400 3936
rect 24452 3924 24458 3936
rect 24688 3924 24716 4023
rect 32122 4020 32128 4032
rect 32180 4020 32186 4072
rect 32950 4020 32956 4072
rect 33008 4060 33014 4072
rect 33229 4063 33287 4069
rect 33229 4060 33241 4063
rect 33008 4032 33241 4060
rect 33008 4020 33014 4032
rect 33229 4029 33241 4032
rect 33275 4029 33287 4063
rect 33888 4060 33916 4091
rect 37366 4088 37372 4100
rect 37424 4088 37430 4140
rect 37458 4088 37464 4140
rect 37516 4128 37522 4140
rect 39850 4128 39856 4140
rect 37516 4100 37561 4128
rect 37844 4100 39856 4128
rect 37516 4088 37522 4100
rect 37844 4060 37872 4100
rect 39850 4088 39856 4100
rect 39908 4088 39914 4140
rect 40405 4131 40463 4137
rect 40405 4097 40417 4131
rect 40451 4128 40463 4131
rect 40586 4128 40592 4140
rect 40451 4100 40592 4128
rect 40451 4097 40463 4100
rect 40405 4091 40463 4097
rect 40586 4088 40592 4100
rect 40644 4088 40650 4140
rect 42426 4128 42432 4140
rect 42387 4100 42432 4128
rect 42426 4088 42432 4100
rect 42484 4088 42490 4140
rect 45830 4088 45836 4140
rect 45888 4128 45894 4140
rect 46566 4128 46572 4140
rect 45888 4100 46428 4128
rect 46527 4100 46572 4128
rect 45888 4088 45894 4100
rect 33888 4032 37872 4060
rect 33229 4023 33287 4029
rect 37918 4020 37924 4072
rect 37976 4060 37982 4072
rect 38565 4063 38623 4069
rect 38565 4060 38577 4063
rect 37976 4032 38577 4060
rect 37976 4020 37982 4032
rect 38565 4029 38577 4032
rect 38611 4029 38623 4063
rect 41782 4060 41788 4072
rect 41743 4032 41788 4060
rect 38565 4023 38623 4029
rect 41782 4020 41788 4032
rect 41840 4020 41846 4072
rect 45186 4060 45192 4072
rect 45147 4032 45192 4060
rect 45186 4020 45192 4032
rect 45244 4020 45250 4072
rect 46201 4063 46259 4069
rect 46201 4029 46213 4063
rect 46247 4060 46259 4063
rect 46290 4060 46296 4072
rect 46247 4032 46296 4060
rect 46247 4029 46259 4032
rect 46201 4023 46259 4029
rect 46290 4020 46296 4032
rect 46348 4020 46354 4072
rect 46400 4060 46428 4100
rect 46566 4088 46572 4100
rect 46624 4088 46630 4140
rect 47765 4131 47823 4137
rect 47765 4097 47777 4131
rect 47811 4128 47823 4131
rect 48222 4128 48228 4140
rect 47811 4100 48228 4128
rect 47811 4097 47823 4100
rect 47765 4091 47823 4097
rect 47780 4060 47808 4091
rect 48222 4088 48228 4100
rect 48280 4088 48286 4140
rect 48409 4131 48467 4137
rect 48409 4097 48421 4131
rect 48455 4128 48467 4131
rect 48590 4128 48596 4140
rect 48455 4100 48596 4128
rect 48455 4097 48467 4100
rect 48409 4091 48467 4097
rect 48590 4088 48596 4100
rect 48648 4088 48654 4140
rect 49050 4088 49056 4140
rect 49108 4128 49114 4140
rect 49326 4128 49332 4140
rect 49108 4100 49332 4128
rect 49108 4088 49114 4100
rect 49326 4088 49332 4100
rect 49384 4128 49390 4140
rect 50157 4131 50215 4137
rect 50157 4128 50169 4131
rect 49384 4100 50169 4128
rect 49384 4088 49390 4100
rect 50157 4097 50169 4100
rect 50203 4097 50215 4131
rect 51905 4131 51963 4137
rect 51905 4128 51917 4131
rect 50157 4091 50215 4097
rect 50264 4100 51917 4128
rect 46400 4032 47808 4060
rect 49694 4020 49700 4072
rect 49752 4060 49758 4072
rect 50264 4060 50292 4100
rect 51905 4097 51917 4100
rect 51951 4097 51963 4131
rect 54662 4128 54668 4140
rect 54623 4100 54668 4128
rect 51905 4091 51963 4097
rect 54662 4088 54668 4100
rect 54720 4088 54726 4140
rect 55214 4088 55220 4140
rect 55272 4128 55278 4140
rect 55766 4128 55772 4140
rect 55272 4100 55317 4128
rect 55727 4100 55772 4128
rect 55272 4088 55278 4100
rect 55766 4088 55772 4100
rect 55824 4088 55830 4140
rect 56318 4128 56324 4140
rect 56279 4100 56324 4128
rect 56318 4088 56324 4100
rect 56376 4088 56382 4140
rect 67358 4128 67364 4140
rect 67319 4100 67364 4128
rect 67358 4088 67364 4100
rect 67416 4088 67422 4140
rect 50614 4060 50620 4072
rect 49752 4032 50292 4060
rect 50575 4032 50620 4060
rect 49752 4020 49758 4032
rect 50614 4020 50620 4032
rect 50672 4020 50678 4072
rect 54021 4063 54079 4069
rect 54021 4060 54033 4063
rect 50724 4032 54033 4060
rect 26418 3992 26424 4004
rect 25608 3964 26424 3992
rect 25608 3924 25636 3964
rect 26418 3952 26424 3964
rect 26476 3952 26482 4004
rect 39022 3952 39028 4004
rect 39080 3992 39086 4004
rect 39850 3992 39856 4004
rect 39080 3964 39856 3992
rect 39080 3952 39086 3964
rect 39850 3952 39856 3964
rect 39908 3952 39914 4004
rect 40402 3952 40408 4004
rect 40460 3992 40466 4004
rect 41141 3995 41199 4001
rect 41141 3992 41153 3995
rect 40460 3964 41153 3992
rect 40460 3952 40466 3964
rect 41141 3961 41153 3964
rect 41187 3961 41199 3995
rect 41141 3955 41199 3961
rect 42426 3952 42432 4004
rect 42484 3992 42490 4004
rect 42484 3964 43576 3992
rect 42484 3952 42490 3964
rect 24452 3896 25636 3924
rect 24452 3884 24458 3896
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 27801 3927 27859 3933
rect 27801 3924 27813 3927
rect 27764 3896 27813 3924
rect 27764 3884 27770 3896
rect 27801 3893 27813 3896
rect 27847 3893 27859 3927
rect 28994 3924 29000 3936
rect 28955 3896 29000 3924
rect 27801 3887 27859 3893
rect 28994 3884 29000 3896
rect 29052 3884 29058 3936
rect 29546 3924 29552 3936
rect 29507 3896 29552 3924
rect 29546 3884 29552 3896
rect 29604 3884 29610 3936
rect 29638 3884 29644 3936
rect 29696 3924 29702 3936
rect 30101 3927 30159 3933
rect 30101 3924 30113 3927
rect 29696 3896 30113 3924
rect 29696 3884 29702 3896
rect 30101 3893 30113 3896
rect 30147 3893 30159 3927
rect 30101 3887 30159 3893
rect 31389 3927 31447 3933
rect 31389 3893 31401 3927
rect 31435 3924 31447 3927
rect 31478 3924 31484 3936
rect 31435 3896 31484 3924
rect 31435 3893 31447 3896
rect 31389 3887 31447 3893
rect 31478 3884 31484 3896
rect 31536 3884 31542 3936
rect 32214 3884 32220 3936
rect 32272 3924 32278 3936
rect 32677 3927 32735 3933
rect 32677 3924 32689 3927
rect 32272 3896 32689 3924
rect 32272 3884 32278 3896
rect 32677 3893 32689 3896
rect 32723 3893 32735 3927
rect 37366 3924 37372 3936
rect 37327 3896 37372 3924
rect 32677 3887 32735 3893
rect 37366 3884 37372 3896
rect 37424 3884 37430 3936
rect 37642 3884 37648 3936
rect 37700 3924 37706 3936
rect 37921 3927 37979 3933
rect 37921 3924 37933 3927
rect 37700 3896 37933 3924
rect 37700 3884 37706 3896
rect 37921 3893 37933 3896
rect 37967 3893 37979 3927
rect 37921 3887 37979 3893
rect 38470 3884 38476 3936
rect 38528 3924 38534 3936
rect 39209 3927 39267 3933
rect 39209 3924 39221 3927
rect 38528 3896 39221 3924
rect 38528 3884 38534 3896
rect 39209 3893 39221 3896
rect 39255 3893 39267 3927
rect 39209 3887 39267 3893
rect 40497 3927 40555 3933
rect 40497 3893 40509 3927
rect 40543 3924 40555 3927
rect 40586 3924 40592 3936
rect 40543 3896 40592 3924
rect 40543 3893 40555 3896
rect 40497 3887 40555 3893
rect 40586 3884 40592 3896
rect 40644 3884 40650 3936
rect 41782 3884 41788 3936
rect 41840 3924 41846 3936
rect 42613 3927 42671 3933
rect 42613 3924 42625 3927
rect 41840 3896 42625 3924
rect 41840 3884 41846 3896
rect 42613 3893 42625 3896
rect 42659 3893 42671 3927
rect 43438 3924 43444 3936
rect 43399 3896 43444 3924
rect 42613 3887 42671 3893
rect 43438 3884 43444 3896
rect 43496 3884 43502 3936
rect 43548 3924 43576 3964
rect 46106 3952 46112 4004
rect 46164 3992 46170 4004
rect 46934 3992 46940 4004
rect 46164 3964 46940 3992
rect 46164 3952 46170 3964
rect 46934 3952 46940 3964
rect 46992 3952 46998 4004
rect 49145 3995 49203 4001
rect 49145 3961 49157 3995
rect 49191 3992 49203 3995
rect 50062 3992 50068 4004
rect 49191 3964 50068 3992
rect 49191 3961 49203 3964
rect 49145 3955 49203 3961
rect 50062 3952 50068 3964
rect 50120 3952 50126 4004
rect 50154 3952 50160 4004
rect 50212 3992 50218 4004
rect 50724 3992 50752 4032
rect 54021 4029 54033 4032
rect 54067 4029 54079 4063
rect 54021 4023 54079 4029
rect 50212 3964 50752 3992
rect 50212 3952 50218 3964
rect 50798 3952 50804 4004
rect 50856 3992 50862 4004
rect 53377 3995 53435 4001
rect 53377 3992 53389 3995
rect 50856 3964 53389 3992
rect 50856 3952 50862 3964
rect 53377 3961 53389 3964
rect 53423 3961 53435 3995
rect 53377 3955 53435 3961
rect 45554 3924 45560 3936
rect 43548 3896 45560 3924
rect 45554 3884 45560 3896
rect 45612 3884 45618 3936
rect 46201 3927 46259 3933
rect 46201 3893 46213 3927
rect 46247 3924 46259 3927
rect 46658 3924 46664 3936
rect 46247 3896 46664 3924
rect 46247 3893 46259 3896
rect 46201 3887 46259 3893
rect 46658 3884 46664 3896
rect 46716 3924 46722 3936
rect 46842 3924 46848 3936
rect 46716 3896 46848 3924
rect 46716 3884 46722 3896
rect 46842 3884 46848 3896
rect 46900 3884 46906 3936
rect 47118 3884 47124 3936
rect 47176 3924 47182 3936
rect 47581 3927 47639 3933
rect 47581 3924 47593 3927
rect 47176 3896 47593 3924
rect 47176 3884 47182 3896
rect 47581 3893 47593 3896
rect 47627 3893 47639 3927
rect 48222 3924 48228 3936
rect 48183 3896 48228 3924
rect 47581 3887 47639 3893
rect 48222 3884 48228 3896
rect 48280 3884 48286 3936
rect 49326 3884 49332 3936
rect 49384 3924 49390 3936
rect 49513 3927 49571 3933
rect 49513 3924 49525 3927
rect 49384 3896 49525 3924
rect 49384 3884 49390 3896
rect 49513 3893 49525 3896
rect 49559 3893 49571 3927
rect 50246 3924 50252 3936
rect 50207 3896 50252 3924
rect 49513 3887 49571 3893
rect 50246 3884 50252 3896
rect 50304 3884 50310 3936
rect 50338 3884 50344 3936
rect 50396 3924 50402 3936
rect 51077 3927 51135 3933
rect 51077 3924 51089 3927
rect 50396 3896 51089 3924
rect 50396 3884 50402 3896
rect 51077 3893 51089 3896
rect 51123 3893 51135 3927
rect 51077 3887 51135 3893
rect 51258 3884 51264 3936
rect 51316 3924 51322 3936
rect 51721 3927 51779 3933
rect 51721 3924 51733 3927
rect 51316 3896 51733 3924
rect 51316 3884 51322 3896
rect 51721 3893 51733 3896
rect 51767 3893 51779 3927
rect 51721 3887 51779 3893
rect 51902 3884 51908 3936
rect 51960 3924 51966 3936
rect 52733 3927 52791 3933
rect 52733 3924 52745 3927
rect 51960 3896 52745 3924
rect 51960 3884 51966 3896
rect 52733 3893 52745 3896
rect 52779 3893 52791 3927
rect 67542 3924 67548 3936
rect 67503 3896 67548 3924
rect 52733 3887 52791 3893
rect 67542 3884 67548 3896
rect 67600 3884 67606 3936
rect 1104 3834 68816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 65654 3834
rect 65706 3782 65718 3834
rect 65770 3782 65782 3834
rect 65834 3782 65846 3834
rect 65898 3782 65910 3834
rect 65962 3782 68816 3834
rect 1104 3760 68816 3782
rect 11606 3720 11612 3732
rect 11567 3692 11612 3720
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 12158 3680 12164 3732
rect 12216 3720 12222 3732
rect 12253 3723 12311 3729
rect 12253 3720 12265 3723
rect 12216 3692 12265 3720
rect 12216 3680 12222 3692
rect 12253 3689 12265 3692
rect 12299 3689 12311 3723
rect 12253 3683 12311 3689
rect 12802 3680 12808 3732
rect 12860 3720 12866 3732
rect 13446 3720 13452 3732
rect 12860 3692 13452 3720
rect 12860 3680 12866 3692
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 14182 3720 14188 3732
rect 14143 3692 14188 3720
rect 14182 3680 14188 3692
rect 14240 3680 14246 3732
rect 14274 3680 14280 3732
rect 14332 3680 14338 3732
rect 14645 3723 14703 3729
rect 14645 3689 14657 3723
rect 14691 3720 14703 3723
rect 14918 3720 14924 3732
rect 14691 3692 14924 3720
rect 14691 3689 14703 3692
rect 14645 3683 14703 3689
rect 14918 3680 14924 3692
rect 14976 3680 14982 3732
rect 15286 3720 15292 3732
rect 15028 3692 15292 3720
rect 10321 3655 10379 3661
rect 10321 3621 10333 3655
rect 10367 3652 10379 3655
rect 12713 3655 12771 3661
rect 12713 3652 12725 3655
rect 10367 3624 12725 3652
rect 10367 3621 10379 3624
rect 10321 3615 10379 3621
rect 12713 3621 12725 3624
rect 12759 3621 12771 3655
rect 14292 3652 14320 3680
rect 15028 3652 15056 3692
rect 15286 3680 15292 3692
rect 15344 3720 15350 3732
rect 15746 3729 15752 3732
rect 15565 3723 15623 3729
rect 15565 3720 15577 3723
rect 15344 3692 15577 3720
rect 15344 3680 15350 3692
rect 15565 3689 15577 3692
rect 15611 3689 15623 3723
rect 15565 3683 15623 3689
rect 15703 3723 15752 3729
rect 15703 3689 15715 3723
rect 15749 3689 15752 3723
rect 15703 3683 15752 3689
rect 15746 3680 15752 3683
rect 15804 3680 15810 3732
rect 16482 3680 16488 3732
rect 16540 3720 16546 3732
rect 16945 3723 17003 3729
rect 16540 3692 16585 3720
rect 16540 3680 16546 3692
rect 16945 3689 16957 3723
rect 16991 3720 17003 3723
rect 17494 3720 17500 3732
rect 16991 3692 17500 3720
rect 16991 3689 17003 3692
rect 16945 3683 17003 3689
rect 17494 3680 17500 3692
rect 17552 3680 17558 3732
rect 20254 3720 20260 3732
rect 20215 3692 20260 3720
rect 20254 3680 20260 3692
rect 20312 3680 20318 3732
rect 25774 3720 25780 3732
rect 25735 3692 25780 3720
rect 25774 3680 25780 3692
rect 25832 3680 25838 3732
rect 30285 3723 30343 3729
rect 30285 3689 30297 3723
rect 30331 3720 30343 3723
rect 31570 3720 31576 3732
rect 30331 3692 31576 3720
rect 30331 3689 30343 3692
rect 30285 3683 30343 3689
rect 31570 3680 31576 3692
rect 31628 3680 31634 3732
rect 32493 3723 32551 3729
rect 32493 3689 32505 3723
rect 32539 3720 32551 3723
rect 32582 3720 32588 3732
rect 32539 3692 32588 3720
rect 32539 3689 32551 3692
rect 32493 3683 32551 3689
rect 32582 3680 32588 3692
rect 32640 3720 32646 3732
rect 33042 3720 33048 3732
rect 32640 3692 33048 3720
rect 32640 3680 32646 3692
rect 33042 3680 33048 3692
rect 33100 3680 33106 3732
rect 35529 3723 35587 3729
rect 35529 3689 35541 3723
rect 35575 3720 35587 3723
rect 39574 3720 39580 3732
rect 35575 3692 39580 3720
rect 35575 3689 35587 3692
rect 35529 3683 35587 3689
rect 39574 3680 39580 3692
rect 39632 3680 39638 3732
rect 42797 3723 42855 3729
rect 42797 3689 42809 3723
rect 42843 3720 42855 3723
rect 42978 3720 42984 3732
rect 42843 3692 42984 3720
rect 42843 3689 42855 3692
rect 42797 3683 42855 3689
rect 42978 3680 42984 3692
rect 43036 3680 43042 3732
rect 43806 3680 43812 3732
rect 43864 3720 43870 3732
rect 45005 3723 45063 3729
rect 43864 3692 44312 3720
rect 43864 3680 43870 3692
rect 14292 3624 15056 3652
rect 19705 3655 19763 3661
rect 12713 3615 12771 3621
rect 19705 3621 19717 3655
rect 19751 3652 19763 3655
rect 20622 3652 20628 3664
rect 19751 3624 20628 3652
rect 19751 3621 19763 3624
rect 19705 3615 19763 3621
rect 20622 3612 20628 3624
rect 20680 3612 20686 3664
rect 38197 3655 38255 3661
rect 38197 3621 38209 3655
rect 38243 3621 38255 3655
rect 38197 3615 38255 3621
rect 7837 3587 7895 3593
rect 7837 3553 7849 3587
rect 7883 3584 7895 3587
rect 10965 3587 11023 3593
rect 7883 3556 10364 3584
rect 7883 3553 7895 3556
rect 7837 3547 7895 3553
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 10137 3519 10195 3525
rect 10137 3516 10149 3519
rect 8168 3488 10149 3516
rect 8168 3476 8174 3488
rect 10137 3485 10149 3488
rect 10183 3485 10195 3519
rect 10336 3516 10364 3556
rect 10965 3553 10977 3587
rect 11011 3584 11023 3587
rect 11606 3584 11612 3596
rect 11011 3556 11612 3584
rect 11011 3553 11023 3556
rect 10965 3547 11023 3553
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 13998 3544 14004 3596
rect 14056 3584 14062 3596
rect 14274 3584 14280 3596
rect 14056 3556 14280 3584
rect 14056 3544 14062 3556
rect 14274 3544 14280 3556
rect 14332 3584 14338 3596
rect 14369 3587 14427 3593
rect 14369 3584 14381 3587
rect 14332 3556 14381 3584
rect 14332 3544 14338 3556
rect 14369 3553 14381 3556
rect 14415 3553 14427 3587
rect 15470 3584 15476 3596
rect 15431 3556 15476 3584
rect 14369 3547 14427 3553
rect 15470 3544 15476 3556
rect 15528 3584 15534 3596
rect 15528 3556 16160 3584
rect 15528 3544 15534 3556
rect 11425 3519 11483 3525
rect 11425 3516 11437 3519
rect 10336 3488 11437 3516
rect 10137 3479 10195 3485
rect 11425 3485 11437 3488
rect 11471 3516 11483 3519
rect 11882 3516 11888 3528
rect 11471 3488 11888 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 8386 3448 8392 3460
rect 8347 3420 8392 3448
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 9033 3451 9091 3457
rect 9033 3417 9045 3451
rect 9079 3448 9091 3451
rect 10152 3448 10180 3479
rect 11882 3476 11888 3488
rect 11940 3476 11946 3528
rect 12066 3516 12072 3528
rect 12027 3488 12072 3516
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 12894 3476 12900 3528
rect 12952 3516 12958 3528
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 12952 3488 13093 3516
rect 12952 3476 12958 3488
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13354 3476 13360 3528
rect 13412 3516 13418 3528
rect 13630 3516 13636 3528
rect 13412 3488 13636 3516
rect 13412 3476 13418 3488
rect 13630 3476 13636 3488
rect 13688 3476 13694 3528
rect 14090 3516 14096 3528
rect 14051 3488 14096 3516
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 15378 3476 15384 3528
rect 15436 3516 15442 3528
rect 16025 3519 16083 3525
rect 16025 3516 16037 3519
rect 15436 3488 16037 3516
rect 15436 3476 15442 3488
rect 16025 3485 16037 3488
rect 16071 3485 16083 3519
rect 16132 3516 16160 3556
rect 16482 3544 16488 3596
rect 16540 3584 16546 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 16540 3556 16589 3584
rect 16540 3544 16546 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 19334 3584 19340 3596
rect 18095 3556 19340 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 19334 3544 19340 3556
rect 19392 3544 19398 3596
rect 20530 3584 20536 3596
rect 20491 3556 20536 3584
rect 20530 3544 20536 3556
rect 20588 3544 20594 3596
rect 24394 3584 24400 3596
rect 24355 3556 24400 3584
rect 24394 3544 24400 3556
rect 24452 3544 24458 3596
rect 26418 3544 26424 3596
rect 26476 3584 26482 3596
rect 29086 3584 29092 3596
rect 26476 3556 29092 3584
rect 26476 3544 26482 3556
rect 29086 3544 29092 3556
rect 29144 3584 29150 3596
rect 30745 3587 30803 3593
rect 30745 3584 30757 3587
rect 29144 3556 30757 3584
rect 29144 3544 29150 3556
rect 30745 3553 30757 3556
rect 30791 3553 30803 3587
rect 30745 3547 30803 3553
rect 32306 3544 32312 3596
rect 32364 3584 32370 3596
rect 33965 3587 34023 3593
rect 33965 3584 33977 3587
rect 32364 3556 33977 3584
rect 32364 3544 32370 3556
rect 33965 3553 33977 3556
rect 34011 3553 34023 3587
rect 33965 3547 34023 3553
rect 35802 3544 35808 3596
rect 35860 3584 35866 3596
rect 35989 3587 36047 3593
rect 35989 3584 36001 3587
rect 35860 3556 36001 3584
rect 35860 3544 35866 3556
rect 35989 3553 36001 3556
rect 36035 3553 36047 3587
rect 35989 3547 36047 3553
rect 36265 3587 36323 3593
rect 36265 3553 36277 3587
rect 36311 3584 36323 3587
rect 38212 3584 38240 3615
rect 42610 3612 42616 3664
rect 42668 3652 42674 3664
rect 44177 3655 44235 3661
rect 44177 3652 44189 3655
rect 42668 3624 44189 3652
rect 42668 3612 42674 3624
rect 44177 3621 44189 3624
rect 44223 3621 44235 3655
rect 44284 3652 44312 3692
rect 45005 3689 45017 3723
rect 45051 3720 45063 3723
rect 45094 3720 45100 3732
rect 45051 3692 45100 3720
rect 45051 3689 45063 3692
rect 45005 3683 45063 3689
rect 45094 3680 45100 3692
rect 45152 3680 45158 3732
rect 46201 3723 46259 3729
rect 46201 3720 46213 3723
rect 45204 3692 46213 3720
rect 45204 3652 45232 3692
rect 46201 3689 46213 3692
rect 46247 3689 46259 3723
rect 46201 3683 46259 3689
rect 47305 3723 47363 3729
rect 47305 3689 47317 3723
rect 47351 3720 47363 3723
rect 47762 3720 47768 3732
rect 47351 3692 47768 3720
rect 47351 3689 47363 3692
rect 47305 3683 47363 3689
rect 47762 3680 47768 3692
rect 47820 3680 47826 3732
rect 48590 3720 48596 3732
rect 48551 3692 48596 3720
rect 48590 3680 48596 3692
rect 48648 3680 48654 3732
rect 50338 3720 50344 3732
rect 48700 3692 50344 3720
rect 46014 3652 46020 3664
rect 44284 3624 45232 3652
rect 45296 3624 46020 3652
rect 44177 3615 44235 3621
rect 36311 3556 38240 3584
rect 40129 3587 40187 3593
rect 36311 3553 36323 3556
rect 36265 3547 36323 3553
rect 40129 3553 40141 3587
rect 40175 3584 40187 3587
rect 40175 3556 41414 3584
rect 40175 3553 40187 3556
rect 40129 3547 40187 3553
rect 16761 3519 16819 3525
rect 16761 3516 16773 3519
rect 16132 3488 16773 3516
rect 16025 3479 16083 3485
rect 16761 3485 16773 3488
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 20070 3516 20076 3528
rect 18739 3488 20076 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 20070 3476 20076 3488
rect 20128 3476 20134 3528
rect 20625 3519 20683 3525
rect 20625 3485 20637 3519
rect 20671 3516 20683 3519
rect 21082 3516 21088 3528
rect 20671 3488 21088 3516
rect 20671 3485 20683 3488
rect 20625 3479 20683 3485
rect 21082 3476 21088 3488
rect 21140 3476 21146 3528
rect 21913 3519 21971 3525
rect 21913 3485 21925 3519
rect 21959 3516 21971 3519
rect 22002 3516 22008 3528
rect 21959 3488 22008 3516
rect 21959 3485 21971 3488
rect 21913 3479 21971 3485
rect 22002 3476 22008 3488
rect 22060 3476 22066 3528
rect 22373 3519 22431 3525
rect 22373 3485 22385 3519
rect 22419 3516 22431 3519
rect 22462 3516 22468 3528
rect 22419 3488 22468 3516
rect 22419 3485 22431 3488
rect 22373 3479 22431 3485
rect 22462 3476 22468 3488
rect 22520 3476 22526 3528
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3516 23259 3519
rect 23566 3516 23572 3528
rect 23247 3488 23572 3516
rect 23247 3485 23259 3488
rect 23201 3479 23259 3485
rect 23566 3476 23572 3488
rect 23624 3476 23630 3528
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 10686 3448 10692 3460
rect 9079 3420 10088 3448
rect 10152 3420 10692 3448
rect 9079 3417 9091 3420
rect 9033 3411 9091 3417
rect 9677 3383 9735 3389
rect 9677 3349 9689 3383
rect 9723 3380 9735 3383
rect 9950 3380 9956 3392
rect 9723 3352 9956 3380
rect 9723 3349 9735 3352
rect 9677 3343 9735 3349
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 10060 3380 10088 3420
rect 10686 3408 10692 3420
rect 10744 3408 10750 3460
rect 11330 3408 11336 3460
rect 11388 3448 11394 3460
rect 12989 3451 13047 3457
rect 12989 3448 13001 3451
rect 11388 3420 13001 3448
rect 11388 3408 11394 3420
rect 12989 3417 13001 3420
rect 13035 3417 13047 3451
rect 12989 3411 13047 3417
rect 13265 3451 13323 3457
rect 13265 3417 13277 3451
rect 13311 3448 13323 3451
rect 13311 3420 16436 3448
rect 13311 3417 13323 3420
rect 13265 3411 13323 3417
rect 12250 3380 12256 3392
rect 10060 3352 12256 3380
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 12897 3383 12955 3389
rect 12897 3380 12909 3383
rect 12676 3352 12909 3380
rect 12676 3340 12682 3352
rect 12897 3349 12909 3352
rect 12943 3349 12955 3383
rect 12897 3343 12955 3349
rect 15197 3383 15255 3389
rect 15197 3349 15209 3383
rect 15243 3380 15255 3383
rect 16114 3380 16120 3392
rect 15243 3352 16120 3380
rect 15243 3349 15255 3352
rect 15197 3343 15255 3349
rect 16114 3340 16120 3352
rect 16172 3340 16178 3392
rect 16408 3380 16436 3420
rect 16482 3408 16488 3460
rect 16540 3448 16546 3460
rect 20165 3451 20223 3457
rect 20165 3448 20177 3451
rect 16540 3420 16585 3448
rect 16776 3420 20177 3448
rect 16540 3408 16546 3420
rect 16776 3380 16804 3420
rect 20165 3417 20177 3420
rect 20211 3417 20223 3451
rect 23860 3448 23888 3479
rect 23934 3476 23940 3528
rect 23992 3516 23998 3528
rect 24653 3519 24711 3525
rect 24653 3516 24665 3519
rect 23992 3488 24665 3516
rect 23992 3476 23998 3488
rect 24653 3485 24665 3488
rect 24699 3485 24711 3519
rect 24653 3479 24711 3485
rect 26050 3476 26056 3528
rect 26108 3516 26114 3528
rect 26237 3519 26295 3525
rect 26237 3516 26249 3519
rect 26108 3488 26249 3516
rect 26108 3476 26114 3488
rect 26237 3485 26249 3488
rect 26283 3485 26295 3519
rect 26237 3479 26295 3485
rect 27065 3519 27123 3525
rect 27065 3485 27077 3519
rect 27111 3516 27123 3519
rect 27430 3516 27436 3528
rect 27111 3488 27436 3516
rect 27111 3485 27123 3488
rect 27065 3479 27123 3485
rect 27430 3476 27436 3488
rect 27488 3476 27494 3528
rect 27709 3519 27767 3525
rect 27709 3485 27721 3519
rect 27755 3516 27767 3519
rect 28258 3516 28264 3528
rect 27755 3488 28264 3516
rect 27755 3485 27767 3488
rect 27709 3479 27767 3485
rect 28258 3476 28264 3488
rect 28316 3476 28322 3528
rect 28353 3519 28411 3525
rect 28353 3485 28365 3519
rect 28399 3516 28411 3519
rect 28810 3516 28816 3528
rect 28399 3488 28816 3516
rect 28399 3485 28411 3488
rect 28353 3479 28411 3485
rect 28810 3476 28816 3488
rect 28868 3476 28874 3528
rect 28997 3519 29055 3525
rect 28997 3485 29009 3519
rect 29043 3516 29055 3519
rect 29454 3516 29460 3528
rect 29043 3488 29460 3516
rect 29043 3485 29055 3488
rect 28997 3479 29055 3485
rect 29454 3476 29460 3488
rect 29512 3476 29518 3528
rect 33226 3476 33232 3528
rect 33284 3516 33290 3528
rect 33321 3519 33379 3525
rect 33321 3516 33333 3519
rect 33284 3488 33333 3516
rect 33284 3476 33290 3488
rect 33321 3485 33333 3488
rect 33367 3485 33379 3519
rect 33321 3479 33379 3485
rect 37366 3476 37372 3528
rect 37424 3476 37430 3528
rect 38381 3519 38439 3525
rect 38381 3485 38393 3519
rect 38427 3516 38439 3519
rect 38562 3516 38568 3528
rect 38427 3488 38568 3516
rect 38427 3485 38439 3488
rect 38381 3479 38439 3485
rect 38562 3476 38568 3488
rect 38620 3476 38626 3528
rect 38933 3519 38991 3525
rect 38933 3485 38945 3519
rect 38979 3516 38991 3519
rect 39022 3516 39028 3528
rect 38979 3488 39028 3516
rect 38979 3485 38991 3488
rect 38933 3479 38991 3485
rect 39022 3476 39028 3488
rect 39080 3476 39086 3528
rect 39850 3516 39856 3528
rect 39811 3488 39856 3516
rect 39850 3476 39856 3488
rect 39908 3476 39914 3528
rect 41386 3516 41414 3556
rect 41966 3544 41972 3596
rect 42024 3584 42030 3596
rect 42245 3587 42303 3593
rect 42245 3584 42257 3587
rect 42024 3556 42257 3584
rect 42024 3544 42030 3556
rect 42245 3553 42257 3556
rect 42291 3584 42303 3587
rect 42426 3584 42432 3596
rect 42291 3556 42432 3584
rect 42291 3553 42303 3556
rect 42245 3547 42303 3553
rect 42426 3544 42432 3556
rect 42484 3544 42490 3596
rect 42518 3544 42524 3596
rect 42576 3584 42582 3596
rect 43438 3584 43444 3596
rect 42576 3556 43444 3584
rect 42576 3544 42582 3556
rect 43438 3544 43444 3556
rect 43496 3584 43502 3596
rect 43496 3556 44128 3584
rect 43496 3544 43502 3556
rect 42794 3516 42800 3528
rect 41386 3488 42800 3516
rect 42794 3476 42800 3488
rect 42852 3476 42858 3528
rect 43548 3525 43576 3556
rect 43533 3519 43591 3525
rect 43533 3485 43545 3519
rect 43579 3485 43591 3519
rect 43533 3479 43591 3485
rect 43993 3519 44051 3525
rect 43993 3485 44005 3519
rect 44039 3485 44051 3519
rect 43993 3479 44051 3485
rect 24394 3448 24400 3460
rect 23860 3420 24400 3448
rect 20165 3411 20223 3417
rect 24394 3408 24400 3420
rect 24452 3408 24458 3460
rect 31018 3448 31024 3460
rect 30979 3420 31024 3448
rect 31018 3408 31024 3420
rect 31076 3408 31082 3460
rect 31478 3408 31484 3460
rect 31536 3408 31542 3460
rect 37752 3420 40172 3448
rect 16408 3352 16804 3380
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 37752 3389 37780 3420
rect 20809 3383 20867 3389
rect 20809 3380 20821 3383
rect 18288 3352 20821 3380
rect 18288 3340 18294 3352
rect 20809 3349 20821 3352
rect 20855 3349 20867 3383
rect 20809 3343 20867 3349
rect 37737 3383 37795 3389
rect 37737 3349 37749 3383
rect 37783 3349 37795 3383
rect 39022 3380 39028 3392
rect 38983 3352 39028 3380
rect 37737 3343 37795 3349
rect 39022 3340 39028 3352
rect 39080 3340 39086 3392
rect 40144 3380 40172 3420
rect 40586 3408 40592 3460
rect 40644 3408 40650 3460
rect 44008 3448 44036 3479
rect 41524 3420 44036 3448
rect 44100 3448 44128 3556
rect 44542 3544 44548 3596
rect 44600 3584 44606 3596
rect 45296 3584 45324 3624
rect 46014 3612 46020 3624
rect 46072 3612 46078 3664
rect 44600 3556 45324 3584
rect 44600 3544 44606 3556
rect 45554 3544 45560 3596
rect 45612 3584 45618 3596
rect 45649 3587 45707 3593
rect 45649 3584 45661 3587
rect 45612 3556 45661 3584
rect 45612 3544 45618 3556
rect 45649 3553 45661 3556
rect 45695 3584 45707 3587
rect 46382 3584 46388 3596
rect 45695 3556 46388 3584
rect 45695 3553 45707 3556
rect 45649 3547 45707 3553
rect 46382 3544 46388 3556
rect 46440 3544 46446 3596
rect 47118 3584 47124 3596
rect 47079 3556 47124 3584
rect 47118 3544 47124 3556
rect 47176 3544 47182 3596
rect 47946 3544 47952 3596
rect 48004 3584 48010 3596
rect 48700 3584 48728 3692
rect 50338 3680 50344 3692
rect 50396 3680 50402 3732
rect 51810 3720 51816 3732
rect 51046 3692 51816 3720
rect 48774 3612 48780 3664
rect 48832 3652 48838 3664
rect 50709 3655 50767 3661
rect 50709 3652 50721 3655
rect 48832 3624 50721 3652
rect 48832 3612 48838 3624
rect 50709 3621 50721 3624
rect 50755 3652 50767 3655
rect 51046 3652 51074 3692
rect 51810 3680 51816 3692
rect 51868 3680 51874 3732
rect 67358 3720 67364 3732
rect 67319 3692 67364 3720
rect 67358 3680 67364 3692
rect 67416 3680 67422 3732
rect 50755 3624 51074 3652
rect 50755 3621 50767 3624
rect 50709 3615 50767 3621
rect 57238 3612 57244 3664
rect 57296 3652 57302 3664
rect 57885 3655 57943 3661
rect 57885 3652 57897 3655
rect 57296 3624 57897 3652
rect 57296 3612 57302 3624
rect 57885 3621 57897 3624
rect 57931 3621 57943 3655
rect 57885 3615 57943 3621
rect 48004 3556 48728 3584
rect 48004 3544 48010 3556
rect 48866 3544 48872 3596
rect 48924 3584 48930 3596
rect 48924 3556 49004 3584
rect 48924 3544 48930 3556
rect 47026 3516 47032 3528
rect 46987 3488 47032 3516
rect 47026 3476 47032 3488
rect 47084 3476 47090 3528
rect 47394 3476 47400 3528
rect 47452 3516 47458 3528
rect 48976 3525 49004 3556
rect 49050 3544 49056 3596
rect 49108 3584 49114 3596
rect 49145 3587 49203 3593
rect 49145 3584 49157 3587
rect 49108 3556 49157 3584
rect 49108 3544 49114 3556
rect 49145 3553 49157 3556
rect 49191 3553 49203 3587
rect 49145 3547 49203 3553
rect 49234 3544 49240 3596
rect 49292 3584 49298 3596
rect 49292 3556 51074 3584
rect 49292 3544 49298 3556
rect 47857 3519 47915 3525
rect 47857 3516 47869 3519
rect 47452 3488 47869 3516
rect 47452 3476 47458 3488
rect 47857 3485 47869 3488
rect 47903 3485 47915 3519
rect 47857 3479 47915 3485
rect 48961 3519 49019 3525
rect 48961 3485 48973 3519
rect 49007 3485 49019 3519
rect 48961 3479 49019 3485
rect 49786 3476 49792 3528
rect 49844 3516 49850 3528
rect 50798 3516 50804 3528
rect 49844 3488 50804 3516
rect 49844 3476 49850 3488
rect 50798 3476 50804 3488
rect 50856 3476 50862 3528
rect 51046 3516 51074 3556
rect 51718 3544 51724 3596
rect 51776 3584 51782 3596
rect 51776 3556 51821 3584
rect 51776 3544 51782 3556
rect 54478 3544 54484 3596
rect 54536 3584 54542 3596
rect 55309 3587 55367 3593
rect 55309 3584 55321 3587
rect 54536 3556 55321 3584
rect 54536 3544 54542 3556
rect 55309 3553 55321 3556
rect 55355 3553 55367 3587
rect 55309 3547 55367 3553
rect 55858 3544 55864 3596
rect 55916 3584 55922 3596
rect 56597 3587 56655 3593
rect 56597 3584 56609 3587
rect 55916 3556 56609 3584
rect 55916 3544 55922 3556
rect 56597 3553 56609 3556
rect 56643 3553 56655 3587
rect 56597 3547 56655 3553
rect 57606 3544 57612 3596
rect 57664 3584 57670 3596
rect 58529 3587 58587 3593
rect 58529 3584 58541 3587
rect 57664 3556 58541 3584
rect 57664 3544 57670 3556
rect 58529 3553 58541 3556
rect 58575 3553 58587 3587
rect 58529 3547 58587 3553
rect 51445 3519 51503 3525
rect 51046 3488 51396 3516
rect 45465 3451 45523 3457
rect 45465 3448 45477 3451
rect 44100 3420 45477 3448
rect 41138 3380 41144 3392
rect 40144 3352 41144 3380
rect 41138 3340 41144 3352
rect 41196 3380 41202 3392
rect 41524 3380 41552 3420
rect 45465 3417 45477 3420
rect 45511 3417 45523 3451
rect 45465 3411 45523 3417
rect 46382 3408 46388 3460
rect 46440 3448 46446 3460
rect 48038 3448 48044 3460
rect 46440 3420 48044 3448
rect 46440 3408 46446 3420
rect 48038 3408 48044 3420
rect 48096 3448 48102 3460
rect 49053 3451 49111 3457
rect 48096 3420 49004 3448
rect 48096 3408 48102 3420
rect 41196 3352 41552 3380
rect 41196 3340 41202 3352
rect 41598 3340 41604 3392
rect 41656 3380 41662 3392
rect 42334 3380 42340 3392
rect 41656 3352 42340 3380
rect 41656 3340 41662 3352
rect 42334 3340 42340 3352
rect 42392 3340 42398 3392
rect 42429 3383 42487 3389
rect 42429 3349 42441 3383
rect 42475 3380 42487 3383
rect 42518 3380 42524 3392
rect 42475 3352 42524 3380
rect 42475 3349 42487 3352
rect 42429 3343 42487 3349
rect 42518 3340 42524 3352
rect 42576 3340 42582 3392
rect 42702 3340 42708 3392
rect 42760 3380 42766 3392
rect 43349 3383 43407 3389
rect 43349 3380 43361 3383
rect 42760 3352 43361 3380
rect 42760 3340 42766 3352
rect 43349 3349 43361 3352
rect 43395 3349 43407 3383
rect 43349 3343 43407 3349
rect 43438 3340 43444 3392
rect 43496 3380 43502 3392
rect 45278 3380 45284 3392
rect 43496 3352 45284 3380
rect 43496 3340 43502 3352
rect 45278 3340 45284 3352
rect 45336 3340 45342 3392
rect 45373 3383 45431 3389
rect 45373 3349 45385 3383
rect 45419 3380 45431 3383
rect 48774 3380 48780 3392
rect 45419 3352 48780 3380
rect 45419 3349 45431 3352
rect 45373 3343 45431 3349
rect 48774 3340 48780 3352
rect 48832 3340 48838 3392
rect 48976 3380 49004 3420
rect 49053 3417 49065 3451
rect 49099 3448 49111 3451
rect 51258 3448 51264 3460
rect 49099 3420 51264 3448
rect 49099 3417 49111 3420
rect 49053 3411 49111 3417
rect 51258 3408 51264 3420
rect 51316 3408 51322 3460
rect 51368 3448 51396 3488
rect 51445 3485 51457 3519
rect 51491 3516 51503 3519
rect 52086 3516 52092 3528
rect 51491 3488 52092 3516
rect 51491 3485 51503 3488
rect 51445 3479 51503 3485
rect 52086 3476 52092 3488
rect 52144 3476 52150 3528
rect 52181 3519 52239 3525
rect 52181 3485 52193 3519
rect 52227 3485 52239 3519
rect 52181 3479 52239 3485
rect 52196 3448 52224 3479
rect 52362 3476 52368 3528
rect 52420 3516 52426 3528
rect 52825 3519 52883 3525
rect 52825 3516 52837 3519
rect 52420 3488 52837 3516
rect 52420 3476 52426 3488
rect 52825 3485 52837 3488
rect 52871 3485 52883 3519
rect 52825 3479 52883 3485
rect 54297 3519 54355 3525
rect 54297 3485 54309 3519
rect 54343 3516 54355 3519
rect 54570 3516 54576 3528
rect 54343 3488 54576 3516
rect 54343 3485 54355 3488
rect 54297 3479 54355 3485
rect 54570 3476 54576 3488
rect 54628 3476 54634 3528
rect 55398 3476 55404 3528
rect 55456 3516 55462 3528
rect 55953 3519 56011 3525
rect 55953 3516 55965 3519
rect 55456 3488 55965 3516
rect 55456 3476 55462 3488
rect 55953 3485 55965 3488
rect 55999 3485 56011 3519
rect 55953 3479 56011 3485
rect 56410 3476 56416 3528
rect 56468 3516 56474 3528
rect 57241 3519 57299 3525
rect 57241 3516 57253 3519
rect 56468 3488 57253 3516
rect 56468 3476 56474 3488
rect 57241 3485 57253 3488
rect 57287 3485 57299 3519
rect 67174 3516 67180 3528
rect 67135 3488 67180 3516
rect 57241 3479 57299 3485
rect 67174 3476 67180 3488
rect 67232 3516 67238 3528
rect 67821 3519 67879 3525
rect 67821 3516 67833 3519
rect 67232 3488 67833 3516
rect 67232 3476 67238 3488
rect 67821 3485 67833 3488
rect 67867 3485 67879 3519
rect 67821 3479 67879 3485
rect 53466 3448 53472 3460
rect 51368 3420 52224 3448
rect 53427 3420 53472 3448
rect 53466 3408 53472 3420
rect 53524 3408 53530 3460
rect 50157 3383 50215 3389
rect 50157 3380 50169 3383
rect 48976 3352 50169 3380
rect 50157 3349 50169 3352
rect 50203 3349 50215 3383
rect 50157 3343 50215 3349
rect 53926 3340 53932 3392
rect 53984 3380 53990 3392
rect 54113 3383 54171 3389
rect 54113 3380 54125 3383
rect 53984 3352 54125 3380
rect 53984 3340 53990 3352
rect 54113 3349 54125 3352
rect 54159 3349 54171 3383
rect 54113 3343 54171 3349
rect 1104 3290 68816 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 68816 3290
rect 1104 3216 68816 3238
rect 7929 3179 7987 3185
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 10226 3176 10232 3188
rect 7975 3148 10232 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 10226 3136 10232 3148
rect 10284 3136 10290 3188
rect 10321 3179 10379 3185
rect 10321 3145 10333 3179
rect 10367 3176 10379 3179
rect 10367 3148 12664 3176
rect 10367 3145 10379 3148
rect 10321 3139 10379 3145
rect 8478 3108 8484 3120
rect 8439 3080 8484 3108
rect 8478 3068 8484 3080
rect 8536 3068 8542 3120
rect 12636 3108 12664 3148
rect 12710 3136 12716 3188
rect 12768 3176 12774 3188
rect 13357 3179 13415 3185
rect 12768 3148 12813 3176
rect 13004 3148 13308 3176
rect 12768 3136 12774 3148
rect 13004 3108 13032 3148
rect 12406 3080 12572 3108
rect 12636 3080 13032 3108
rect 13280 3108 13308 3148
rect 13357 3145 13369 3179
rect 13403 3176 13415 3179
rect 14461 3179 14519 3185
rect 13403 3148 14320 3176
rect 13403 3145 13415 3148
rect 13357 3139 13415 3145
rect 14292 3108 14320 3148
rect 14461 3145 14473 3179
rect 14507 3176 14519 3179
rect 15102 3176 15108 3188
rect 14507 3148 15108 3176
rect 14507 3145 14519 3148
rect 14461 3139 14519 3145
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 16482 3176 16488 3188
rect 15620 3148 16488 3176
rect 15620 3136 15626 3148
rect 16482 3136 16488 3148
rect 16540 3136 16546 3188
rect 19978 3176 19984 3188
rect 19939 3148 19984 3176
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 21082 3176 21088 3188
rect 21043 3148 21088 3176
rect 21082 3136 21088 3148
rect 21140 3136 21146 3188
rect 29546 3136 29552 3188
rect 29604 3176 29610 3188
rect 30837 3179 30895 3185
rect 29604 3148 29776 3176
rect 29604 3136 29610 3148
rect 15194 3108 15200 3120
rect 13280 3080 14228 3108
rect 14292 3080 15200 3108
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3040 7435 3043
rect 10134 3040 10140 3052
rect 7423 3012 10140 3040
rect 7423 3009 7435 3012
rect 7377 3003 7435 3009
rect 10134 3000 10140 3012
rect 10192 3000 10198 3052
rect 10226 3000 10232 3052
rect 10284 3040 10290 3052
rect 12406 3040 12434 3080
rect 10284 3012 12434 3040
rect 12544 3040 12572 3080
rect 12621 3043 12679 3049
rect 12621 3040 12633 3043
rect 12544 3012 12633 3040
rect 10284 3000 10290 3012
rect 12621 3009 12633 3012
rect 12667 3040 12679 3043
rect 13096 3040 13216 3044
rect 13354 3040 13360 3052
rect 12667 3016 13360 3040
rect 12667 3012 13124 3016
rect 13188 3012 13360 3016
rect 12667 3009 12679 3012
rect 12621 3003 12679 3009
rect 13354 3000 13360 3012
rect 13412 3000 13418 3052
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 9033 2975 9091 2981
rect 9033 2941 9045 2975
rect 9079 2972 9091 2975
rect 10962 2972 10968 2984
rect 9079 2944 10968 2972
rect 9079 2941 9091 2944
rect 9033 2935 9091 2941
rect 10962 2932 10968 2944
rect 11020 2932 11026 2984
rect 12066 2972 12072 2984
rect 12027 2944 12072 2972
rect 12066 2932 12072 2944
rect 12124 2932 12130 2984
rect 12250 2932 12256 2984
rect 12308 2972 12314 2984
rect 13464 2972 13492 3003
rect 13906 3000 13912 3052
rect 13964 3040 13970 3052
rect 14001 3043 14059 3049
rect 14001 3040 14013 3043
rect 13964 3012 14013 3040
rect 13964 3000 13970 3012
rect 14001 3009 14013 3012
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14090 2972 14096 2984
rect 12308 2944 13492 2972
rect 14051 2944 14096 2972
rect 12308 2932 12314 2944
rect 9677 2907 9735 2913
rect 9677 2873 9689 2907
rect 9723 2904 9735 2907
rect 13464 2904 13492 2944
rect 14090 2932 14096 2944
rect 14148 2932 14154 2984
rect 14200 2972 14228 3080
rect 15194 3068 15200 3080
rect 15252 3068 15258 3120
rect 17313 3111 17371 3117
rect 17313 3077 17325 3111
rect 17359 3108 17371 3111
rect 19058 3108 19064 3120
rect 17359 3080 19064 3108
rect 17359 3077 17371 3080
rect 17313 3071 17371 3077
rect 19058 3068 19064 3080
rect 19116 3068 19122 3120
rect 29365 3111 29423 3117
rect 29365 3077 29377 3111
rect 29411 3108 29423 3111
rect 29638 3108 29644 3120
rect 29411 3080 29644 3108
rect 29411 3077 29423 3080
rect 29365 3071 29423 3077
rect 29638 3068 29644 3080
rect 29696 3068 29702 3120
rect 29748 3108 29776 3148
rect 30837 3145 30849 3179
rect 30883 3145 30895 3179
rect 30837 3139 30895 3145
rect 30852 3108 30880 3139
rect 31018 3136 31024 3188
rect 31076 3176 31082 3188
rect 31389 3179 31447 3185
rect 31389 3176 31401 3179
rect 31076 3148 31401 3176
rect 31076 3136 31082 3148
rect 31389 3145 31401 3148
rect 31435 3145 31447 3179
rect 32122 3176 32128 3188
rect 32083 3148 32128 3176
rect 31389 3139 31447 3145
rect 32122 3136 32128 3148
rect 32180 3136 32186 3188
rect 32582 3176 32588 3188
rect 32543 3148 32588 3176
rect 32582 3136 32588 3148
rect 32640 3136 32646 3188
rect 38289 3179 38347 3185
rect 38289 3145 38301 3179
rect 38335 3176 38347 3179
rect 38838 3176 38844 3188
rect 38335 3148 38844 3176
rect 38335 3145 38347 3148
rect 38289 3139 38347 3145
rect 38838 3136 38844 3148
rect 38896 3136 38902 3188
rect 39850 3136 39856 3188
rect 39908 3176 39914 3188
rect 43714 3176 43720 3188
rect 39908 3148 43720 3176
rect 39908 3136 39914 3148
rect 29748 3080 29854 3108
rect 30852 3080 32536 3108
rect 14274 3000 14280 3052
rect 14332 3040 14338 3052
rect 14332 3012 14377 3040
rect 14332 3000 14338 3012
rect 14734 3000 14740 3052
rect 14792 3040 14798 3052
rect 17129 3043 17187 3049
rect 17129 3040 17141 3043
rect 14792 3012 17141 3040
rect 14792 3000 14798 3012
rect 17129 3009 17141 3012
rect 17175 3009 17187 3043
rect 19794 3040 19800 3052
rect 19755 3012 19800 3040
rect 17129 3003 17187 3009
rect 19794 3000 19800 3012
rect 19852 3000 19858 3052
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3040 21327 3043
rect 21818 3040 21824 3052
rect 21315 3012 21824 3040
rect 21315 3009 21327 3012
rect 21269 3003 21327 3009
rect 21818 3000 21824 3012
rect 21876 3000 21882 3052
rect 29086 3040 29092 3052
rect 29047 3012 29092 3040
rect 29086 3000 29092 3012
rect 29144 3000 29150 3052
rect 31573 3043 31631 3049
rect 31573 3009 31585 3043
rect 31619 3040 31631 3043
rect 32214 3040 32220 3052
rect 31619 3012 32220 3040
rect 31619 3009 31631 3012
rect 31573 3003 31631 3009
rect 32214 3000 32220 3012
rect 32272 3000 32278 3052
rect 32508 3049 32536 3080
rect 39022 3068 39028 3120
rect 39080 3068 39086 3120
rect 39758 3108 39764 3120
rect 39719 3080 39764 3108
rect 39758 3068 39764 3080
rect 39816 3068 39822 3120
rect 40052 3049 40080 3148
rect 43714 3136 43720 3148
rect 43772 3176 43778 3188
rect 45186 3176 45192 3188
rect 43772 3148 45192 3176
rect 43772 3136 43778 3148
rect 45186 3136 45192 3148
rect 45244 3176 45250 3188
rect 45244 3148 45416 3176
rect 45244 3136 45250 3148
rect 41138 3068 41144 3120
rect 41196 3108 41202 3120
rect 41601 3111 41659 3117
rect 41601 3108 41613 3111
rect 41196 3080 41613 3108
rect 41196 3068 41202 3080
rect 41601 3077 41613 3080
rect 41647 3077 41659 3111
rect 41601 3071 41659 3077
rect 42058 3068 42064 3120
rect 42116 3108 42122 3120
rect 42702 3108 42708 3120
rect 42116 3080 42708 3108
rect 42116 3068 42122 3080
rect 42702 3068 42708 3080
rect 42760 3068 42766 3120
rect 43530 3068 43536 3120
rect 43588 3108 43594 3120
rect 43588 3080 43838 3108
rect 43588 3068 43594 3080
rect 32493 3043 32551 3049
rect 32493 3009 32505 3043
rect 32539 3040 32551 3043
rect 40037 3043 40095 3049
rect 32539 3012 38516 3040
rect 32539 3009 32551 3012
rect 32493 3003 32551 3009
rect 15378 2972 15384 2984
rect 14200 2944 15384 2972
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15470 2932 15476 2984
rect 15528 2972 15534 2984
rect 15933 2975 15991 2981
rect 15933 2972 15945 2975
rect 15528 2944 15945 2972
rect 15528 2932 15534 2944
rect 15933 2941 15945 2944
rect 15979 2941 15991 2975
rect 15933 2935 15991 2941
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2972 19395 2975
rect 20898 2972 20904 2984
rect 19383 2944 20904 2972
rect 19383 2941 19395 2944
rect 19337 2935 19395 2941
rect 20898 2932 20904 2944
rect 20956 2932 20962 2984
rect 23201 2975 23259 2981
rect 23201 2941 23213 2975
rect 23247 2972 23259 2975
rect 23842 2972 23848 2984
rect 23247 2944 23848 2972
rect 23247 2941 23259 2944
rect 23201 2935 23259 2941
rect 23842 2932 23848 2944
rect 23900 2932 23906 2984
rect 25133 2975 25191 2981
rect 25133 2941 25145 2975
rect 25179 2972 25191 2975
rect 25774 2972 25780 2984
rect 25179 2944 25780 2972
rect 25179 2941 25191 2944
rect 25133 2935 25191 2941
rect 25774 2932 25780 2944
rect 25832 2932 25838 2984
rect 27985 2975 28043 2981
rect 27985 2941 27997 2975
rect 28031 2972 28043 2975
rect 29362 2972 29368 2984
rect 28031 2944 29368 2972
rect 28031 2941 28043 2944
rect 27985 2935 28043 2941
rect 29362 2932 29368 2944
rect 29420 2932 29426 2984
rect 32766 2972 32772 2984
rect 32679 2944 32772 2972
rect 32766 2932 32772 2944
rect 32824 2972 32830 2984
rect 32950 2972 32956 2984
rect 32824 2944 32956 2972
rect 32824 2932 32830 2944
rect 32950 2932 32956 2944
rect 33008 2932 33014 2984
rect 9723 2876 12848 2904
rect 13464 2876 14136 2904
rect 9723 2873 9735 2876
rect 9677 2867 9735 2873
rect 10870 2796 10876 2848
rect 10928 2836 10934 2848
rect 10965 2839 11023 2845
rect 10965 2836 10977 2839
rect 10928 2808 10977 2836
rect 10928 2796 10934 2808
rect 10965 2805 10977 2808
rect 11011 2805 11023 2839
rect 12820 2836 12848 2876
rect 14108 2848 14136 2876
rect 14458 2864 14464 2916
rect 14516 2904 14522 2916
rect 15105 2907 15163 2913
rect 15105 2904 15117 2907
rect 14516 2876 15117 2904
rect 14516 2864 14522 2876
rect 15105 2873 15117 2876
rect 15151 2873 15163 2907
rect 15105 2867 15163 2873
rect 15194 2864 15200 2916
rect 15252 2904 15258 2916
rect 17310 2904 17316 2916
rect 15252 2876 17316 2904
rect 15252 2864 15258 2876
rect 17310 2864 17316 2876
rect 17368 2864 17374 2916
rect 18049 2907 18107 2913
rect 18049 2873 18061 2907
rect 18095 2904 18107 2907
rect 19426 2904 19432 2916
rect 18095 2876 19432 2904
rect 18095 2873 18107 2876
rect 18049 2867 18107 2873
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 19794 2864 19800 2916
rect 19852 2904 19858 2916
rect 21266 2904 21272 2916
rect 19852 2876 21272 2904
rect 19852 2864 19858 2876
rect 21266 2864 21272 2876
rect 21324 2864 21330 2916
rect 24946 2904 24952 2916
rect 23860 2876 24952 2904
rect 13078 2836 13084 2848
rect 12820 2808 13084 2836
rect 10965 2799 11023 2805
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 14090 2796 14096 2848
rect 14148 2796 14154 2848
rect 14182 2796 14188 2848
rect 14240 2836 14246 2848
rect 14240 2808 14285 2836
rect 14240 2796 14246 2808
rect 15286 2796 15292 2848
rect 15344 2836 15350 2848
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 15344 2808 15485 2836
rect 15344 2796 15350 2808
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 15562 2796 15568 2848
rect 15620 2836 15626 2848
rect 18693 2839 18751 2845
rect 15620 2808 15665 2836
rect 15620 2796 15626 2808
rect 18693 2805 18705 2839
rect 18739 2836 18751 2839
rect 20346 2836 20352 2848
rect 18739 2808 20352 2836
rect 18739 2805 18751 2808
rect 18693 2799 18751 2805
rect 20346 2796 20352 2808
rect 20404 2796 20410 2848
rect 20625 2839 20683 2845
rect 20625 2805 20637 2839
rect 20671 2836 20683 2839
rect 21450 2836 21456 2848
rect 20671 2808 21456 2836
rect 20671 2805 20683 2808
rect 20625 2799 20683 2805
rect 21450 2796 21456 2808
rect 21508 2796 21514 2848
rect 22557 2839 22615 2845
rect 22557 2805 22569 2839
rect 22603 2836 22615 2839
rect 23290 2836 23296 2848
rect 22603 2808 23296 2836
rect 22603 2805 22615 2808
rect 22557 2799 22615 2805
rect 23290 2796 23296 2808
rect 23348 2796 23354 2848
rect 23860 2845 23888 2876
rect 24946 2864 24952 2876
rect 25004 2864 25010 2916
rect 27341 2907 27399 2913
rect 27341 2873 27353 2907
rect 27387 2904 27399 2907
rect 28534 2904 28540 2916
rect 27387 2876 28540 2904
rect 27387 2873 27399 2876
rect 27341 2867 27399 2873
rect 28534 2864 28540 2876
rect 28592 2864 28598 2916
rect 38194 2864 38200 2916
rect 38252 2904 38258 2916
rect 38488 2904 38516 3012
rect 40037 3009 40049 3043
rect 40083 3009 40095 3043
rect 41506 3040 41512 3052
rect 41467 3012 41512 3040
rect 40037 3003 40095 3009
rect 41506 3000 41512 3012
rect 41564 3000 41570 3052
rect 41874 3000 41880 3052
rect 41932 3040 41938 3052
rect 42429 3043 42487 3049
rect 42429 3040 42441 3043
rect 41932 3012 42441 3040
rect 41932 3000 41938 3012
rect 42429 3009 42441 3012
rect 42475 3009 42487 3043
rect 42429 3003 42487 3009
rect 45281 3043 45339 3049
rect 45281 3009 45293 3043
rect 45327 3040 45339 3043
rect 45388 3040 45416 3148
rect 48590 3136 48596 3188
rect 48648 3176 48654 3188
rect 49694 3176 49700 3188
rect 48648 3148 49464 3176
rect 49655 3148 49700 3176
rect 48648 3136 48654 3148
rect 48406 3068 48412 3120
rect 48464 3108 48470 3120
rect 49234 3108 49240 3120
rect 48464 3080 49240 3108
rect 48464 3068 48470 3080
rect 49234 3068 49240 3080
rect 49292 3068 49298 3120
rect 49436 3108 49464 3148
rect 49694 3136 49700 3148
rect 49752 3136 49758 3188
rect 50357 3179 50415 3185
rect 50357 3176 50369 3179
rect 49804 3148 50369 3176
rect 49513 3111 49571 3117
rect 49513 3108 49525 3111
rect 49436 3080 49525 3108
rect 45327 3012 45416 3040
rect 46017 3043 46075 3049
rect 45327 3009 45339 3012
rect 45281 3003 45339 3009
rect 46017 3009 46029 3043
rect 46063 3040 46075 3043
rect 49326 3040 49332 3052
rect 46063 3012 49332 3040
rect 46063 3009 46075 3012
rect 46017 3003 46075 3009
rect 38562 2932 38568 2984
rect 38620 2972 38626 2984
rect 41785 2975 41843 2981
rect 38620 2944 39988 2972
rect 38620 2932 38626 2944
rect 38654 2904 38660 2916
rect 38252 2876 38424 2904
rect 38488 2876 38660 2904
rect 38252 2864 38258 2876
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2805 23903 2839
rect 23845 2799 23903 2805
rect 24489 2839 24547 2845
rect 24489 2805 24501 2839
rect 24535 2836 24547 2839
rect 25498 2836 25504 2848
rect 24535 2808 25504 2836
rect 24535 2805 24547 2808
rect 24489 2799 24547 2805
rect 25498 2796 25504 2808
rect 25556 2796 25562 2848
rect 25777 2839 25835 2845
rect 25777 2805 25789 2839
rect 25823 2836 25835 2839
rect 26326 2836 26332 2848
rect 25823 2808 26332 2836
rect 25823 2805 25835 2808
rect 25777 2799 25835 2805
rect 26326 2796 26332 2808
rect 26384 2796 26390 2848
rect 26421 2839 26479 2845
rect 26421 2805 26433 2839
rect 26467 2836 26479 2839
rect 26878 2836 26884 2848
rect 26467 2808 26884 2836
rect 26467 2805 26479 2808
rect 26421 2799 26479 2805
rect 26878 2796 26884 2808
rect 26936 2796 26942 2848
rect 28629 2839 28687 2845
rect 28629 2805 28641 2839
rect 28675 2836 28687 2839
rect 30466 2836 30472 2848
rect 28675 2808 30472 2836
rect 28675 2805 28687 2808
rect 28629 2799 28687 2805
rect 30466 2796 30472 2808
rect 30524 2796 30530 2848
rect 33778 2836 33784 2848
rect 33739 2808 33784 2836
rect 33778 2796 33784 2808
rect 33836 2796 33842 2848
rect 34241 2839 34299 2845
rect 34241 2805 34253 2839
rect 34287 2836 34299 2839
rect 34330 2836 34336 2848
rect 34287 2808 34336 2836
rect 34287 2805 34299 2808
rect 34241 2799 34299 2805
rect 34330 2796 34336 2808
rect 34388 2796 34394 2848
rect 34790 2796 34796 2848
rect 34848 2836 34854 2848
rect 34885 2839 34943 2845
rect 34885 2836 34897 2839
rect 34848 2808 34897 2836
rect 34848 2796 34854 2808
rect 34885 2805 34897 2808
rect 34931 2805 34943 2839
rect 34885 2799 34943 2805
rect 35434 2796 35440 2848
rect 35492 2836 35498 2848
rect 35529 2839 35587 2845
rect 35529 2836 35541 2839
rect 35492 2808 35541 2836
rect 35492 2796 35498 2808
rect 35529 2805 35541 2808
rect 35575 2805 35587 2839
rect 35529 2799 35587 2805
rect 36262 2796 36268 2848
rect 36320 2836 36326 2848
rect 36357 2839 36415 2845
rect 36357 2836 36369 2839
rect 36320 2808 36369 2836
rect 36320 2796 36326 2808
rect 36357 2805 36369 2808
rect 36403 2805 36415 2839
rect 36357 2799 36415 2805
rect 36814 2796 36820 2848
rect 36872 2836 36878 2848
rect 37277 2839 37335 2845
rect 37277 2836 37289 2839
rect 36872 2808 37289 2836
rect 36872 2796 36878 2808
rect 37277 2805 37289 2808
rect 37323 2805 37335 2839
rect 38396 2836 38424 2876
rect 38654 2864 38660 2876
rect 38712 2864 38718 2916
rect 39960 2904 39988 2944
rect 41785 2941 41797 2975
rect 41831 2972 41843 2975
rect 41966 2972 41972 2984
rect 41831 2944 41972 2972
rect 41831 2941 41843 2944
rect 41785 2935 41843 2941
rect 41966 2932 41972 2944
rect 42024 2932 42030 2984
rect 42334 2932 42340 2984
rect 42392 2972 42398 2984
rect 44266 2972 44272 2984
rect 42392 2944 44272 2972
rect 42392 2932 42398 2944
rect 44266 2932 44272 2944
rect 44324 2932 44330 2984
rect 45005 2975 45063 2981
rect 45005 2941 45017 2975
rect 45051 2972 45063 2975
rect 48222 2972 48228 2984
rect 45051 2944 48228 2972
rect 45051 2941 45063 2944
rect 45005 2935 45063 2941
rect 48222 2932 48228 2944
rect 48280 2932 48286 2984
rect 49160 2981 49188 3012
rect 49326 3000 49332 3012
rect 49384 3000 49390 3052
rect 49145 2975 49203 2981
rect 49145 2941 49157 2975
rect 49191 2941 49203 2975
rect 49436 2972 49464 3080
rect 49513 3077 49525 3080
rect 49559 3077 49571 3111
rect 49513 3071 49571 3077
rect 49602 3068 49608 3120
rect 49660 3108 49666 3120
rect 49804 3108 49832 3148
rect 50357 3145 50369 3148
rect 50403 3145 50415 3179
rect 50357 3139 50415 3145
rect 50525 3179 50583 3185
rect 50525 3145 50537 3179
rect 50571 3176 50583 3179
rect 50706 3176 50712 3188
rect 50571 3148 50712 3176
rect 50571 3145 50583 3148
rect 50525 3139 50583 3145
rect 50706 3136 50712 3148
rect 50764 3136 50770 3188
rect 49660 3080 49832 3108
rect 49660 3068 49666 3080
rect 50062 3068 50068 3120
rect 50120 3108 50126 3120
rect 50157 3111 50215 3117
rect 50157 3108 50169 3111
rect 50120 3080 50169 3108
rect 50120 3068 50126 3080
rect 50157 3077 50169 3080
rect 50203 3077 50215 3111
rect 54662 3108 54668 3120
rect 50157 3071 50215 3077
rect 53760 3080 54668 3108
rect 50080 2972 50108 3068
rect 51810 3040 51816 3052
rect 51771 3012 51816 3040
rect 51810 3000 51816 3012
rect 51868 3000 51874 3052
rect 52730 3040 52736 3052
rect 52691 3012 52736 3040
rect 52730 3000 52736 3012
rect 52788 3000 52794 3052
rect 53760 3049 53788 3080
rect 54662 3068 54668 3080
rect 54720 3068 54726 3120
rect 54754 3068 54760 3120
rect 54812 3108 54818 3120
rect 56778 3108 56784 3120
rect 54812 3080 56784 3108
rect 54812 3068 54818 3080
rect 56778 3068 56784 3080
rect 56836 3068 56842 3120
rect 53745 3043 53803 3049
rect 53745 3009 53757 3043
rect 53791 3009 53803 3043
rect 53745 3003 53803 3009
rect 54481 3043 54539 3049
rect 54481 3009 54493 3043
rect 54527 3040 54539 3043
rect 55122 3040 55128 3052
rect 54527 3012 55128 3040
rect 54527 3009 54539 3012
rect 54481 3003 54539 3009
rect 55122 3000 55128 3012
rect 55180 3000 55186 3052
rect 55217 3043 55275 3049
rect 55217 3009 55229 3043
rect 55263 3040 55275 3043
rect 55306 3040 55312 3052
rect 55263 3012 55312 3040
rect 55263 3009 55275 3012
rect 55217 3003 55275 3009
rect 55306 3000 55312 3012
rect 55364 3000 55370 3052
rect 49436 2944 50108 2972
rect 49145 2935 49203 2941
rect 39960 2876 40632 2904
rect 40497 2839 40555 2845
rect 40497 2836 40509 2839
rect 38396 2808 40509 2836
rect 37277 2799 37335 2805
rect 40497 2805 40509 2808
rect 40543 2805 40555 2839
rect 40604 2836 40632 2876
rect 41046 2864 41052 2916
rect 41104 2904 41110 2916
rect 42613 2907 42671 2913
rect 42613 2904 42625 2907
rect 41104 2876 42625 2904
rect 41104 2864 41110 2876
rect 42613 2873 42625 2876
rect 42659 2873 42671 2907
rect 42613 2867 42671 2873
rect 43162 2864 43168 2916
rect 43220 2904 43226 2916
rect 43220 2876 43668 2904
rect 43220 2864 43226 2876
rect 41141 2839 41199 2845
rect 41141 2836 41153 2839
rect 40604 2808 41153 2836
rect 40497 2799 40555 2805
rect 41141 2805 41153 2808
rect 41187 2805 41199 2839
rect 41141 2799 41199 2805
rect 42242 2796 42248 2848
rect 42300 2836 42306 2848
rect 42518 2836 42524 2848
rect 42300 2808 42524 2836
rect 42300 2796 42306 2808
rect 42518 2796 42524 2808
rect 42576 2796 42582 2848
rect 42794 2796 42800 2848
rect 42852 2836 42858 2848
rect 43530 2836 43536 2848
rect 42852 2808 43536 2836
rect 42852 2796 42858 2808
rect 43530 2796 43536 2808
rect 43588 2796 43594 2848
rect 43640 2836 43668 2876
rect 45278 2864 45284 2916
rect 45336 2904 45342 2916
rect 46477 2907 46535 2913
rect 46477 2904 46489 2907
rect 45336 2876 46489 2904
rect 45336 2864 45342 2876
rect 46477 2873 46489 2876
rect 46523 2873 46535 2907
rect 47578 2904 47584 2916
rect 47539 2876 47584 2904
rect 46477 2867 46535 2873
rect 47578 2864 47584 2876
rect 47636 2864 47642 2916
rect 49160 2904 49188 2935
rect 51718 2932 51724 2984
rect 51776 2972 51782 2984
rect 55677 2975 55735 2981
rect 55677 2972 55689 2975
rect 51776 2944 55689 2972
rect 51776 2932 51782 2944
rect 55677 2941 55689 2944
rect 55723 2941 55735 2975
rect 55677 2935 55735 2941
rect 56962 2932 56968 2984
rect 57020 2972 57026 2984
rect 57885 2975 57943 2981
rect 57885 2972 57897 2975
rect 57020 2944 57897 2972
rect 57020 2932 57026 2944
rect 57885 2941 57897 2944
rect 57931 2941 57943 2975
rect 57885 2935 57943 2941
rect 49160 2876 49648 2904
rect 45833 2839 45891 2845
rect 45833 2836 45845 2839
rect 43640 2808 45845 2836
rect 45833 2805 45845 2808
rect 45879 2805 45891 2839
rect 45833 2799 45891 2805
rect 46014 2796 46020 2848
rect 46072 2836 46078 2848
rect 48225 2839 48283 2845
rect 48225 2836 48237 2839
rect 46072 2808 48237 2836
rect 46072 2796 46078 2808
rect 48225 2805 48237 2808
rect 48271 2805 48283 2839
rect 49510 2836 49516 2848
rect 49471 2808 49516 2836
rect 48225 2799 48283 2805
rect 49510 2796 49516 2808
rect 49568 2796 49574 2848
rect 49620 2836 49648 2876
rect 50614 2864 50620 2916
rect 50672 2904 50678 2916
rect 51166 2904 51172 2916
rect 50672 2876 51172 2904
rect 50672 2864 50678 2876
rect 51166 2864 51172 2876
rect 51224 2864 51230 2916
rect 52822 2864 52828 2916
rect 52880 2904 52886 2916
rect 53561 2907 53619 2913
rect 53561 2904 53573 2907
rect 52880 2876 53573 2904
rect 52880 2864 52886 2876
rect 53561 2873 53573 2876
rect 53607 2873 53619 2907
rect 53561 2867 53619 2873
rect 54202 2864 54208 2916
rect 54260 2904 54266 2916
rect 55033 2907 55091 2913
rect 55033 2904 55045 2907
rect 54260 2876 55045 2904
rect 54260 2864 54266 2876
rect 55033 2873 55045 2876
rect 55079 2873 55091 2907
rect 55033 2867 55091 2873
rect 55122 2864 55128 2916
rect 55180 2904 55186 2916
rect 56321 2907 56379 2913
rect 56321 2904 56333 2907
rect 55180 2876 56333 2904
rect 55180 2864 55186 2876
rect 56321 2873 56333 2876
rect 56367 2873 56379 2907
rect 56321 2867 56379 2873
rect 57514 2864 57520 2916
rect 57572 2904 57578 2916
rect 58529 2907 58587 2913
rect 58529 2904 58541 2907
rect 57572 2876 58541 2904
rect 57572 2864 57578 2876
rect 58529 2873 58541 2876
rect 58575 2873 58587 2907
rect 58529 2867 58587 2873
rect 50341 2839 50399 2845
rect 50341 2836 50353 2839
rect 49620 2808 50353 2836
rect 50341 2805 50353 2808
rect 50387 2805 50399 2839
rect 51074 2836 51080 2848
rect 51035 2808 51080 2836
rect 50341 2799 50399 2805
rect 51074 2796 51080 2808
rect 51132 2796 51138 2848
rect 51442 2796 51448 2848
rect 51500 2836 51506 2848
rect 51629 2839 51687 2845
rect 51629 2836 51641 2839
rect 51500 2808 51641 2836
rect 51500 2796 51506 2808
rect 51629 2805 51641 2808
rect 51675 2805 51687 2839
rect 51629 2799 51687 2805
rect 52270 2796 52276 2848
rect 52328 2836 52334 2848
rect 52917 2839 52975 2845
rect 52917 2836 52929 2839
rect 52328 2808 52929 2836
rect 52328 2796 52334 2808
rect 52917 2805 52929 2808
rect 52963 2805 52975 2839
rect 52917 2799 52975 2805
rect 53374 2796 53380 2848
rect 53432 2836 53438 2848
rect 54297 2839 54355 2845
rect 54297 2836 54309 2839
rect 53432 2808 54309 2836
rect 53432 2796 53438 2808
rect 54297 2805 54309 2808
rect 54343 2805 54355 2839
rect 54297 2799 54355 2805
rect 55582 2796 55588 2848
rect 55640 2836 55646 2848
rect 56965 2839 57023 2845
rect 56965 2836 56977 2839
rect 55640 2808 56977 2836
rect 55640 2796 55646 2808
rect 56965 2805 56977 2808
rect 57011 2805 57023 2839
rect 56965 2799 57023 2805
rect 1104 2746 68816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 65654 2746
rect 65706 2694 65718 2746
rect 65770 2694 65782 2746
rect 65834 2694 65846 2746
rect 65898 2694 65910 2746
rect 65962 2694 68816 2746
rect 1104 2672 68816 2694
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 14461 2635 14519 2641
rect 11020 2604 14044 2632
rect 11020 2592 11026 2604
rect 8389 2567 8447 2573
rect 8389 2533 8401 2567
rect 8435 2564 8447 2567
rect 11330 2564 11336 2576
rect 8435 2536 11336 2564
rect 8435 2533 8447 2536
rect 8389 2527 8447 2533
rect 11330 2524 11336 2536
rect 11388 2524 11394 2576
rect 12342 2524 12348 2576
rect 12400 2564 12406 2576
rect 12526 2564 12532 2576
rect 12400 2536 12532 2564
rect 12400 2524 12406 2536
rect 12526 2524 12532 2536
rect 12584 2524 12590 2576
rect 7745 2499 7803 2505
rect 7745 2465 7757 2499
rect 7791 2496 7803 2499
rect 12434 2496 12440 2508
rect 7791 2468 12440 2496
rect 7791 2465 7803 2468
rect 7745 2459 7803 2465
rect 12434 2456 12440 2468
rect 12492 2496 12498 2508
rect 12710 2496 12716 2508
rect 12492 2468 12572 2496
rect 12671 2468 12716 2496
rect 12492 2456 12498 2468
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 8202 2428 8208 2440
rect 6687 2400 8208 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 9674 2428 9680 2440
rect 9635 2400 9680 2428
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10962 2428 10968 2440
rect 10923 2400 10968 2428
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 12544 2437 12572 2468
rect 12710 2456 12716 2468
rect 12768 2456 12774 2508
rect 12529 2431 12587 2437
rect 12529 2397 12541 2431
rect 12575 2397 12587 2431
rect 14016 2428 14044 2604
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 14642 2632 14648 2644
rect 14507 2604 14648 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 14642 2592 14648 2604
rect 14700 2592 14706 2644
rect 16022 2632 16028 2644
rect 15983 2604 16028 2632
rect 16022 2592 16028 2604
rect 16080 2592 16086 2644
rect 16758 2632 16764 2644
rect 16719 2604 16764 2632
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 19337 2635 19395 2641
rect 19337 2601 19349 2635
rect 19383 2632 19395 2635
rect 19794 2632 19800 2644
rect 19383 2604 19800 2632
rect 19383 2601 19395 2604
rect 19337 2595 19395 2601
rect 19794 2592 19800 2604
rect 19852 2592 19858 2644
rect 19981 2635 20039 2641
rect 19981 2601 19993 2635
rect 20027 2632 20039 2635
rect 20254 2632 20260 2644
rect 20027 2604 20260 2632
rect 20027 2601 20039 2604
rect 19981 2595 20039 2601
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 32217 2635 32275 2641
rect 32217 2601 32229 2635
rect 32263 2632 32275 2635
rect 32766 2632 32772 2644
rect 32263 2604 32772 2632
rect 32263 2601 32275 2604
rect 32217 2595 32275 2601
rect 32766 2592 32772 2604
rect 32824 2592 32830 2644
rect 56137 2635 56195 2641
rect 56137 2632 56149 2635
rect 35866 2604 56149 2632
rect 15102 2564 15108 2576
rect 15063 2536 15108 2564
rect 15102 2524 15108 2536
rect 15160 2524 15166 2576
rect 17494 2564 17500 2576
rect 17455 2536 17500 2564
rect 17494 2524 17500 2536
rect 17552 2524 17558 2576
rect 18693 2567 18751 2573
rect 18693 2533 18705 2567
rect 18739 2564 18751 2567
rect 21174 2564 21180 2576
rect 18739 2536 21180 2564
rect 18739 2533 18751 2536
rect 18693 2527 18751 2533
rect 21174 2524 21180 2536
rect 21232 2524 21238 2576
rect 22557 2567 22615 2573
rect 22557 2533 22569 2567
rect 22603 2564 22615 2567
rect 24118 2564 24124 2576
rect 22603 2536 24124 2564
rect 22603 2533 22615 2536
rect 22557 2527 22615 2533
rect 24118 2524 24124 2536
rect 24176 2524 24182 2576
rect 25777 2567 25835 2573
rect 25777 2533 25789 2567
rect 25823 2564 25835 2567
rect 27154 2564 27160 2576
rect 25823 2536 27160 2564
rect 25823 2533 25835 2536
rect 25777 2527 25835 2533
rect 27154 2524 27160 2536
rect 27212 2524 27218 2576
rect 27709 2567 27767 2573
rect 27709 2533 27721 2567
rect 27755 2564 27767 2567
rect 30190 2564 30196 2576
rect 27755 2536 30196 2564
rect 27755 2533 27767 2536
rect 27709 2527 27767 2533
rect 30190 2524 30196 2536
rect 30248 2524 30254 2576
rect 30285 2567 30343 2573
rect 30285 2533 30297 2567
rect 30331 2564 30343 2567
rect 32398 2564 32404 2576
rect 30331 2536 32404 2564
rect 30331 2533 30343 2536
rect 30285 2527 30343 2533
rect 32398 2524 32404 2536
rect 32456 2524 32462 2576
rect 32861 2567 32919 2573
rect 32861 2533 32873 2567
rect 32907 2564 32919 2567
rect 33502 2564 33508 2576
rect 32907 2536 33508 2564
rect 32907 2533 32919 2536
rect 32861 2527 32919 2533
rect 33502 2524 33508 2536
rect 33560 2524 33566 2576
rect 15286 2456 15292 2508
rect 15344 2456 15350 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 22186 2496 22192 2508
rect 20671 2468 22192 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 22186 2456 22192 2468
rect 22244 2456 22250 2508
rect 23201 2499 23259 2505
rect 23201 2465 23213 2499
rect 23247 2496 23259 2499
rect 24670 2496 24676 2508
rect 23247 2468 24676 2496
rect 23247 2465 23259 2468
rect 23201 2459 23259 2465
rect 24670 2456 24676 2468
rect 24728 2456 24734 2508
rect 25133 2499 25191 2505
rect 25133 2465 25145 2499
rect 25179 2496 25191 2499
rect 26421 2499 26479 2505
rect 25179 2468 25912 2496
rect 25179 2465 25191 2468
rect 25133 2459 25191 2465
rect 14645 2431 14703 2437
rect 14645 2428 14657 2431
rect 14016 2400 14657 2428
rect 12529 2391 12587 2397
rect 14645 2397 14657 2400
rect 14691 2428 14703 2431
rect 15304 2428 15332 2456
rect 17678 2428 17684 2440
rect 14691 2400 15332 2428
rect 17639 2400 17684 2428
rect 14691 2397 14703 2400
rect 14645 2391 14703 2397
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 19797 2431 19855 2437
rect 19797 2397 19809 2431
rect 19843 2397 19855 2431
rect 19797 2391 19855 2397
rect 21269 2431 21327 2437
rect 21269 2397 21281 2431
rect 21315 2428 21327 2431
rect 22738 2428 22744 2440
rect 21315 2400 22744 2428
rect 21315 2397 21327 2400
rect 21269 2391 21327 2397
rect 7193 2363 7251 2369
rect 7193 2329 7205 2363
rect 7239 2360 7251 2363
rect 11698 2360 11704 2372
rect 7239 2332 11704 2360
rect 7239 2329 7251 2332
rect 7193 2323 7251 2329
rect 11698 2320 11704 2332
rect 11756 2360 11762 2372
rect 11885 2363 11943 2369
rect 11885 2360 11897 2363
rect 11756 2332 11897 2360
rect 11756 2320 11762 2332
rect 11885 2329 11897 2332
rect 11931 2329 11943 2363
rect 11885 2323 11943 2329
rect 11974 2320 11980 2372
rect 12032 2360 12038 2372
rect 12069 2363 12127 2369
rect 12069 2360 12081 2363
rect 12032 2332 12081 2360
rect 12032 2320 12038 2332
rect 12069 2329 12081 2332
rect 12115 2329 12127 2363
rect 15289 2363 15347 2369
rect 12069 2323 12127 2329
rect 12360 2332 15240 2360
rect 9033 2295 9091 2301
rect 9033 2261 9045 2295
rect 9079 2292 9091 2295
rect 12360 2292 12388 2332
rect 9079 2264 12388 2292
rect 13541 2295 13599 2301
rect 9079 2261 9091 2264
rect 9033 2255 9091 2261
rect 13541 2261 13553 2295
rect 13587 2292 13599 2295
rect 14734 2292 14740 2304
rect 13587 2264 14740 2292
rect 13587 2261 13599 2264
rect 13541 2255 13599 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 15212 2292 15240 2332
rect 15289 2329 15301 2363
rect 15335 2360 15347 2363
rect 15378 2360 15384 2372
rect 15335 2332 15384 2360
rect 15335 2329 15347 2332
rect 15289 2323 15347 2329
rect 15378 2320 15384 2332
rect 15436 2320 15442 2372
rect 15933 2363 15991 2369
rect 15933 2329 15945 2363
rect 15979 2329 15991 2363
rect 15933 2323 15991 2329
rect 15838 2292 15844 2304
rect 15212 2264 15844 2292
rect 15838 2252 15844 2264
rect 15896 2292 15902 2304
rect 15948 2292 15976 2323
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 16853 2363 16911 2369
rect 16853 2360 16865 2363
rect 16448 2332 16865 2360
rect 16448 2320 16454 2332
rect 16853 2329 16865 2332
rect 16899 2329 16911 2363
rect 19812 2360 19840 2391
rect 22738 2388 22744 2400
rect 22796 2388 22802 2440
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2428 23903 2431
rect 25222 2428 25228 2440
rect 23891 2400 25228 2428
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 25222 2388 25228 2400
rect 25280 2388 25286 2440
rect 25884 2428 25912 2468
rect 26421 2465 26433 2499
rect 26467 2496 26479 2499
rect 27982 2496 27988 2508
rect 26467 2468 27988 2496
rect 26467 2465 26479 2468
rect 26421 2459 26479 2465
rect 27982 2456 27988 2468
rect 28040 2456 28046 2508
rect 28353 2499 28411 2505
rect 28353 2465 28365 2499
rect 28399 2496 28411 2499
rect 30742 2496 30748 2508
rect 28399 2468 30748 2496
rect 28399 2465 28411 2468
rect 28353 2459 28411 2465
rect 30742 2456 30748 2468
rect 30800 2456 30806 2508
rect 30929 2499 30987 2505
rect 30929 2465 30941 2499
rect 30975 2496 30987 2499
rect 32674 2496 32680 2508
rect 30975 2468 32680 2496
rect 30975 2465 30987 2468
rect 30929 2459 30987 2465
rect 32674 2456 32680 2468
rect 32732 2456 32738 2508
rect 28997 2431 29055 2437
rect 25884 2400 26234 2428
rect 19812 2332 21588 2360
rect 16853 2323 16911 2329
rect 21560 2304 21588 2332
rect 21634 2320 21640 2372
rect 21692 2360 21698 2372
rect 24397 2363 24455 2369
rect 24397 2360 24409 2363
rect 21692 2332 24409 2360
rect 21692 2320 21698 2332
rect 24397 2329 24409 2332
rect 24443 2329 24455 2363
rect 26206 2360 26234 2400
rect 28997 2397 29009 2431
rect 29043 2428 29055 2431
rect 31294 2428 31300 2440
rect 29043 2400 31300 2428
rect 29043 2397 29055 2400
rect 28997 2391 29055 2397
rect 31294 2388 31300 2400
rect 31352 2388 31358 2440
rect 31573 2431 31631 2437
rect 31573 2397 31585 2431
rect 31619 2428 31631 2431
rect 32950 2428 32956 2440
rect 31619 2400 32956 2428
rect 31619 2397 31631 2400
rect 31573 2391 31631 2397
rect 32950 2388 32956 2400
rect 33008 2388 33014 2440
rect 33505 2431 33563 2437
rect 33505 2397 33517 2431
rect 33551 2428 33563 2431
rect 34054 2428 34060 2440
rect 33551 2400 34060 2428
rect 33551 2397 33563 2400
rect 33505 2391 33563 2397
rect 34054 2388 34060 2400
rect 34112 2388 34118 2440
rect 34149 2431 34207 2437
rect 34149 2397 34161 2431
rect 34195 2428 34207 2431
rect 34606 2428 34612 2440
rect 34195 2400 34612 2428
rect 34195 2397 34207 2400
rect 34149 2391 34207 2397
rect 34606 2388 34612 2400
rect 34664 2388 34670 2440
rect 34977 2431 35035 2437
rect 34977 2397 34989 2431
rect 35023 2428 35035 2431
rect 35158 2428 35164 2440
rect 35023 2400 35164 2428
rect 35023 2397 35035 2400
rect 34977 2391 35035 2397
rect 35158 2388 35164 2400
rect 35216 2388 35222 2440
rect 35621 2431 35679 2437
rect 35621 2397 35633 2431
rect 35667 2428 35679 2431
rect 35710 2428 35716 2440
rect 35667 2400 35716 2428
rect 35667 2397 35679 2400
rect 35621 2391 35679 2397
rect 35710 2388 35716 2400
rect 35768 2388 35774 2440
rect 26602 2360 26608 2372
rect 26206 2332 26608 2360
rect 24397 2323 24455 2329
rect 26602 2320 26608 2332
rect 26660 2320 26666 2372
rect 30650 2320 30656 2372
rect 30708 2360 30714 2372
rect 35866 2360 35894 2604
rect 56137 2601 56149 2604
rect 56183 2601 56195 2635
rect 56778 2632 56784 2644
rect 56739 2604 56784 2632
rect 56137 2595 56195 2601
rect 56778 2592 56784 2604
rect 56836 2592 56842 2644
rect 40402 2524 40408 2576
rect 40460 2564 40466 2576
rect 41509 2567 41567 2573
rect 41509 2564 41521 2567
rect 40460 2536 41521 2564
rect 40460 2524 40466 2536
rect 41509 2533 41521 2536
rect 41555 2533 41567 2567
rect 41509 2527 41567 2533
rect 41598 2524 41604 2576
rect 41656 2564 41662 2576
rect 44085 2567 44143 2573
rect 44085 2564 44097 2567
rect 41656 2536 44097 2564
rect 41656 2524 41662 2536
rect 44085 2533 44097 2536
rect 44131 2533 44143 2567
rect 44085 2527 44143 2533
rect 44266 2524 44272 2576
rect 44324 2564 44330 2576
rect 45189 2567 45247 2573
rect 45189 2564 45201 2567
rect 44324 2536 45201 2564
rect 44324 2524 44330 2536
rect 45189 2533 45201 2536
rect 45235 2533 45247 2567
rect 45189 2527 45247 2533
rect 45833 2567 45891 2573
rect 45833 2533 45845 2567
rect 45879 2533 45891 2567
rect 45833 2527 45891 2533
rect 37090 2456 37096 2508
rect 37148 2496 37154 2508
rect 37921 2499 37979 2505
rect 37921 2496 37933 2499
rect 37148 2468 37933 2496
rect 37148 2456 37154 2468
rect 37921 2465 37933 2468
rect 37967 2465 37979 2499
rect 37921 2459 37979 2465
rect 39301 2499 39359 2505
rect 39301 2465 39313 2499
rect 39347 2496 39359 2499
rect 39942 2496 39948 2508
rect 39347 2468 39948 2496
rect 39347 2465 39359 2468
rect 39301 2459 39359 2465
rect 39942 2456 39948 2468
rect 40000 2496 40006 2508
rect 42794 2496 42800 2508
rect 40000 2468 42800 2496
rect 40000 2456 40006 2468
rect 35986 2388 35992 2440
rect 36044 2428 36050 2440
rect 36081 2431 36139 2437
rect 36081 2428 36093 2431
rect 36044 2400 36093 2428
rect 36044 2388 36050 2400
rect 36081 2397 36093 2400
rect 36127 2397 36139 2431
rect 36081 2391 36139 2397
rect 36538 2388 36544 2440
rect 36596 2428 36602 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36596 2400 37289 2428
rect 36596 2388 36602 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 37366 2388 37372 2440
rect 37424 2428 37430 2440
rect 38565 2431 38623 2437
rect 38565 2428 38577 2431
rect 37424 2400 38577 2428
rect 37424 2388 37430 2400
rect 38565 2397 38577 2400
rect 38611 2397 38623 2431
rect 40218 2428 40224 2440
rect 40179 2400 40224 2428
rect 38565 2391 38623 2397
rect 40218 2388 40224 2400
rect 40276 2388 40282 2440
rect 40954 2428 40960 2440
rect 40915 2400 40960 2428
rect 40954 2388 40960 2400
rect 41012 2388 41018 2440
rect 41708 2437 41736 2468
rect 42794 2456 42800 2468
rect 42852 2456 42858 2508
rect 42886 2456 42892 2508
rect 42944 2496 42950 2508
rect 45848 2496 45876 2527
rect 46290 2524 46296 2576
rect 46348 2564 46354 2576
rect 46477 2567 46535 2573
rect 46477 2564 46489 2567
rect 46348 2536 46489 2564
rect 46348 2524 46354 2536
rect 46477 2533 46489 2536
rect 46523 2533 46535 2567
rect 46477 2527 46535 2533
rect 46658 2524 46664 2576
rect 46716 2564 46722 2576
rect 49329 2567 49387 2573
rect 49329 2564 49341 2567
rect 46716 2536 49341 2564
rect 46716 2524 46722 2536
rect 49329 2533 49341 2536
rect 49375 2533 49387 2567
rect 49329 2527 49387 2533
rect 52546 2524 52552 2576
rect 52604 2564 52610 2576
rect 53653 2567 53711 2573
rect 53653 2564 53665 2567
rect 52604 2536 53665 2564
rect 52604 2524 52610 2536
rect 53653 2533 53665 2536
rect 53699 2533 53711 2567
rect 53653 2527 53711 2533
rect 56686 2524 56692 2576
rect 56744 2564 56750 2576
rect 58529 2567 58587 2573
rect 58529 2564 58541 2567
rect 56744 2536 58541 2564
rect 56744 2524 56750 2536
rect 58529 2533 58541 2536
rect 58575 2533 58587 2567
rect 58529 2527 58587 2533
rect 42944 2468 45876 2496
rect 42944 2456 42950 2468
rect 47486 2456 47492 2508
rect 47544 2496 47550 2508
rect 47949 2499 48007 2505
rect 47949 2496 47961 2499
rect 47544 2468 47961 2496
rect 47544 2456 47550 2468
rect 47949 2465 47961 2468
rect 47995 2465 48007 2499
rect 47949 2459 48007 2465
rect 49878 2456 49884 2508
rect 49936 2496 49942 2508
rect 51074 2496 51080 2508
rect 49936 2468 51080 2496
rect 49936 2456 49942 2468
rect 51074 2456 51080 2468
rect 51132 2456 51138 2508
rect 54018 2496 54024 2508
rect 53024 2468 54024 2496
rect 41693 2431 41751 2437
rect 41693 2397 41705 2431
rect 41739 2428 41751 2431
rect 41739 2400 41773 2428
rect 41739 2397 41751 2400
rect 41693 2391 41751 2397
rect 42150 2388 42156 2440
rect 42208 2428 42214 2440
rect 42429 2431 42487 2437
rect 42429 2428 42441 2431
rect 42208 2400 42441 2428
rect 42208 2388 42214 2400
rect 42429 2397 42441 2400
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 42518 2388 42524 2440
rect 42576 2428 42582 2440
rect 43165 2431 43223 2437
rect 43165 2428 43177 2431
rect 42576 2400 43177 2428
rect 42576 2388 42582 2400
rect 43165 2397 43177 2400
rect 43211 2397 43223 2431
rect 43898 2428 43904 2440
rect 43859 2400 43904 2428
rect 43165 2391 43223 2397
rect 43898 2388 43904 2400
rect 43956 2388 43962 2440
rect 45005 2431 45063 2437
rect 45005 2397 45017 2431
rect 45051 2397 45063 2431
rect 45005 2391 45063 2397
rect 46017 2431 46075 2437
rect 46017 2397 46029 2431
rect 46063 2428 46075 2431
rect 48590 2428 48596 2440
rect 46063 2400 48596 2428
rect 46063 2397 46075 2400
rect 46017 2391 46075 2397
rect 30708 2332 35894 2360
rect 41386 2332 42656 2360
rect 30708 2320 30714 2332
rect 15896 2264 15976 2292
rect 15896 2252 15902 2264
rect 21542 2252 21548 2304
rect 21600 2292 21606 2304
rect 21821 2295 21879 2301
rect 21821 2292 21833 2295
rect 21600 2264 21833 2292
rect 21600 2252 21606 2264
rect 21821 2261 21833 2264
rect 21867 2261 21879 2295
rect 21821 2255 21879 2261
rect 39850 2252 39856 2304
rect 39908 2292 39914 2304
rect 40037 2295 40095 2301
rect 40037 2292 40049 2295
rect 39908 2264 40049 2292
rect 39908 2252 39914 2264
rect 40037 2261 40049 2264
rect 40083 2261 40095 2295
rect 40037 2255 40095 2261
rect 40126 2252 40132 2304
rect 40184 2292 40190 2304
rect 40773 2295 40831 2301
rect 40773 2292 40785 2295
rect 40184 2264 40785 2292
rect 40184 2252 40190 2264
rect 40773 2261 40785 2264
rect 40819 2261 40831 2295
rect 40773 2255 40831 2261
rect 40862 2252 40868 2304
rect 40920 2292 40926 2304
rect 41386 2292 41414 2332
rect 42628 2301 42656 2332
rect 42794 2320 42800 2372
rect 42852 2360 42858 2372
rect 45020 2360 45048 2391
rect 48590 2388 48596 2400
rect 48648 2388 48654 2440
rect 48685 2431 48743 2437
rect 48685 2397 48697 2431
rect 48731 2397 48743 2431
rect 48685 2391 48743 2397
rect 46658 2360 46664 2372
rect 42852 2332 45048 2360
rect 46492 2332 46664 2360
rect 42852 2320 42858 2332
rect 40920 2264 41414 2292
rect 42613 2295 42671 2301
rect 40920 2252 40926 2264
rect 42613 2261 42625 2295
rect 42659 2261 42671 2295
rect 42613 2255 42671 2261
rect 42702 2252 42708 2304
rect 42760 2292 42766 2304
rect 43349 2295 43407 2301
rect 43349 2292 43361 2295
rect 42760 2264 43361 2292
rect 42760 2252 42766 2264
rect 43349 2261 43361 2264
rect 43395 2261 43407 2295
rect 43349 2255 43407 2261
rect 45002 2252 45008 2304
rect 45060 2292 45066 2304
rect 46492 2292 46520 2332
rect 46658 2320 46664 2332
rect 46716 2320 46722 2372
rect 47854 2320 47860 2372
rect 47912 2360 47918 2372
rect 48133 2363 48191 2369
rect 48133 2360 48145 2363
rect 47912 2332 48145 2360
rect 47912 2320 47918 2332
rect 48133 2329 48145 2332
rect 48179 2329 48191 2363
rect 48133 2323 48191 2329
rect 48222 2320 48228 2372
rect 48280 2360 48286 2372
rect 48700 2360 48728 2391
rect 48958 2388 48964 2440
rect 49016 2428 49022 2440
rect 49513 2431 49571 2437
rect 49513 2428 49525 2431
rect 49016 2400 49525 2428
rect 49016 2388 49022 2400
rect 49513 2397 49525 2400
rect 49559 2397 49571 2431
rect 49513 2391 49571 2397
rect 48280 2332 48728 2360
rect 49528 2360 49556 2391
rect 49602 2388 49608 2440
rect 49660 2428 49666 2440
rect 50341 2431 50399 2437
rect 50341 2428 50353 2431
rect 49660 2400 50353 2428
rect 49660 2388 49666 2400
rect 50341 2397 50353 2400
rect 50387 2397 50399 2431
rect 51258 2428 51264 2440
rect 51219 2400 51264 2428
rect 50341 2391 50399 2397
rect 51258 2388 51264 2400
rect 51316 2388 51322 2440
rect 51626 2388 51632 2440
rect 51684 2428 51690 2440
rect 53024 2437 53052 2468
rect 54018 2456 54024 2468
rect 54076 2456 54082 2508
rect 55766 2496 55772 2508
rect 55186 2468 55772 2496
rect 51721 2431 51779 2437
rect 51721 2428 51733 2431
rect 51684 2400 51733 2428
rect 51684 2388 51690 2400
rect 51721 2397 51733 2400
rect 51767 2397 51779 2431
rect 51721 2391 51779 2397
rect 53009 2431 53067 2437
rect 53009 2397 53021 2431
rect 53055 2397 53067 2431
rect 53009 2391 53067 2397
rect 53282 2388 53288 2440
rect 53340 2428 53346 2440
rect 53469 2431 53527 2437
rect 53469 2428 53481 2431
rect 53340 2400 53481 2428
rect 53340 2388 53346 2400
rect 53469 2397 53481 2400
rect 53515 2397 53527 2431
rect 53469 2391 53527 2397
rect 54481 2431 54539 2437
rect 54481 2397 54493 2431
rect 54527 2428 54539 2431
rect 55186 2428 55214 2468
rect 55766 2456 55772 2468
rect 55824 2456 55830 2508
rect 57422 2456 57428 2508
rect 57480 2496 57486 2508
rect 59173 2499 59231 2505
rect 59173 2496 59185 2499
rect 57480 2468 59185 2496
rect 57480 2456 57486 2468
rect 59173 2465 59185 2468
rect 59219 2465 59231 2499
rect 59173 2459 59231 2465
rect 54527 2400 55214 2428
rect 55585 2431 55643 2437
rect 54527 2397 54539 2400
rect 54481 2391 54539 2397
rect 55585 2397 55597 2431
rect 55631 2428 55643 2431
rect 56318 2428 56324 2440
rect 55631 2400 56324 2428
rect 55631 2397 55643 2400
rect 55585 2391 55643 2397
rect 56318 2388 56324 2400
rect 56376 2388 56382 2440
rect 57885 2431 57943 2437
rect 57885 2397 57897 2431
rect 57931 2397 57943 2431
rect 57885 2391 57943 2397
rect 51350 2360 51356 2372
rect 49528 2332 51356 2360
rect 48280 2320 48286 2332
rect 51350 2320 51356 2332
rect 51408 2320 51414 2372
rect 53650 2320 53656 2372
rect 53708 2360 53714 2372
rect 53708 2332 55214 2360
rect 53708 2320 53714 2332
rect 45060 2264 46520 2292
rect 45060 2252 45066 2264
rect 46566 2252 46572 2304
rect 46624 2292 46630 2304
rect 50157 2295 50215 2301
rect 50157 2292 50169 2295
rect 46624 2264 50169 2292
rect 46624 2252 46630 2264
rect 50157 2261 50169 2264
rect 50203 2261 50215 2295
rect 50157 2255 50215 2261
rect 50890 2252 50896 2304
rect 50948 2292 50954 2304
rect 51077 2295 51135 2301
rect 51077 2292 51089 2295
rect 50948 2264 51089 2292
rect 50948 2252 50954 2264
rect 51077 2261 51089 2264
rect 51123 2261 51135 2295
rect 51077 2255 51135 2261
rect 51166 2252 51172 2304
rect 51224 2292 51230 2304
rect 51905 2295 51963 2301
rect 51905 2292 51917 2295
rect 51224 2264 51917 2292
rect 51224 2252 51230 2264
rect 51905 2261 51917 2264
rect 51951 2261 51963 2295
rect 51905 2255 51963 2261
rect 51994 2252 52000 2304
rect 52052 2292 52058 2304
rect 52825 2295 52883 2301
rect 52825 2292 52837 2295
rect 52052 2264 52837 2292
rect 52052 2252 52058 2264
rect 52825 2261 52837 2264
rect 52871 2261 52883 2295
rect 52825 2255 52883 2261
rect 53098 2252 53104 2304
rect 53156 2292 53162 2304
rect 54297 2295 54355 2301
rect 54297 2292 54309 2295
rect 53156 2264 54309 2292
rect 53156 2252 53162 2264
rect 54297 2261 54309 2264
rect 54343 2261 54355 2295
rect 55186 2292 55214 2332
rect 55490 2320 55496 2372
rect 55548 2360 55554 2372
rect 55950 2360 55956 2372
rect 55548 2332 55956 2360
rect 55548 2320 55554 2332
rect 55950 2320 55956 2332
rect 56008 2360 56014 2372
rect 56229 2363 56287 2369
rect 56229 2360 56241 2363
rect 56008 2332 56241 2360
rect 56008 2320 56014 2332
rect 56229 2329 56241 2332
rect 56275 2329 56287 2363
rect 56229 2323 56287 2329
rect 55401 2295 55459 2301
rect 55401 2292 55413 2295
rect 55186 2264 55413 2292
rect 54297 2255 54355 2261
rect 55401 2261 55413 2264
rect 55447 2261 55459 2295
rect 55401 2255 55459 2261
rect 56134 2252 56140 2304
rect 56192 2292 56198 2304
rect 57900 2292 57928 2391
rect 56192 2264 57928 2292
rect 56192 2252 56198 2264
rect 1104 2202 68816 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 68816 2202
rect 1104 2128 68816 2150
rect 8202 2048 8208 2100
rect 8260 2088 8266 2100
rect 12710 2088 12716 2100
rect 8260 2060 12716 2088
rect 8260 2048 8266 2060
rect 12710 2048 12716 2060
rect 12768 2048 12774 2100
rect 17678 2048 17684 2100
rect 17736 2088 17742 2100
rect 21634 2088 21640 2100
rect 17736 2060 21640 2088
rect 17736 2048 17742 2060
rect 21634 2048 21640 2060
rect 21692 2048 21698 2100
rect 40218 2048 40224 2100
rect 40276 2088 40282 2100
rect 44358 2088 44364 2100
rect 40276 2060 44364 2088
rect 40276 2048 40282 2060
rect 44358 2048 44364 2060
rect 44416 2048 44422 2100
rect 46658 2048 46664 2100
rect 46716 2088 46722 2100
rect 49878 2088 49884 2100
rect 46716 2060 49884 2088
rect 46716 2048 46722 2060
rect 49878 2048 49884 2060
rect 49936 2048 49942 2100
rect 9674 1980 9680 2032
rect 9732 2020 9738 2032
rect 14826 2020 14832 2032
rect 9732 1992 14832 2020
rect 9732 1980 9738 1992
rect 14826 1980 14832 1992
rect 14884 1980 14890 2032
rect 41322 1980 41328 2032
rect 41380 2020 41386 2032
rect 43898 2020 43904 2032
rect 41380 1992 43904 2020
rect 41380 1980 41386 1992
rect 43898 1980 43904 1992
rect 43956 1980 43962 2032
rect 44266 1980 44272 2032
rect 44324 2020 44330 2032
rect 48222 2020 48228 2032
rect 44324 1992 48228 2020
rect 44324 1980 44330 1992
rect 48222 1980 48228 1992
rect 48280 1980 48286 2032
rect 10318 1912 10324 1964
rect 10376 1952 10382 1964
rect 15378 1952 15384 1964
rect 10376 1924 15384 1952
rect 10376 1912 10382 1924
rect 15378 1912 15384 1924
rect 15436 1912 15442 1964
rect 40954 1912 40960 1964
rect 41012 1952 41018 1964
rect 48498 1952 48504 1964
rect 41012 1924 48504 1952
rect 41012 1912 41018 1924
rect 48498 1912 48504 1924
rect 48556 1912 48562 1964
rect 12158 1844 12164 1896
rect 12216 1884 12222 1896
rect 16298 1884 16304 1896
rect 12216 1856 16304 1884
rect 12216 1844 12222 1856
rect 16298 1844 16304 1856
rect 16356 1844 16362 1896
rect 45094 1844 45100 1896
rect 45152 1884 45158 1896
rect 47394 1884 47400 1896
rect 45152 1856 47400 1884
rect 45152 1844 45158 1856
rect 47394 1844 47400 1856
rect 47452 1844 47458 1896
rect 11698 1776 11704 1828
rect 11756 1816 11762 1828
rect 12986 1816 12992 1828
rect 11756 1788 12992 1816
rect 11756 1776 11762 1788
rect 12986 1776 12992 1788
rect 13044 1776 13050 1828
rect 41230 1776 41236 1828
rect 41288 1816 41294 1828
rect 42702 1816 42708 1828
rect 41288 1788 42708 1816
rect 41288 1776 41294 1788
rect 42702 1776 42708 1788
rect 42760 1776 42766 1828
rect 45554 1776 45560 1828
rect 45612 1816 45618 1828
rect 49142 1816 49148 1828
rect 45612 1788 49148 1816
rect 45612 1776 45618 1788
rect 49142 1776 49148 1788
rect 49200 1816 49206 1828
rect 49602 1816 49608 1828
rect 49200 1788 49608 1816
rect 49200 1776 49206 1788
rect 49602 1776 49608 1788
rect 49660 1776 49666 1828
rect 11422 1708 11428 1760
rect 11480 1748 11486 1760
rect 12894 1748 12900 1760
rect 11480 1720 12900 1748
rect 11480 1708 11486 1720
rect 12894 1708 12900 1720
rect 12952 1708 12958 1760
rect 16114 1708 16120 1760
rect 16172 1748 16178 1760
rect 16390 1748 16396 1760
rect 16172 1720 16396 1748
rect 16172 1708 16178 1720
rect 16390 1708 16396 1720
rect 16448 1708 16454 1760
rect 47210 1708 47216 1760
rect 47268 1748 47274 1760
rect 47854 1748 47860 1760
rect 47268 1720 47860 1748
rect 47268 1708 47274 1720
rect 47854 1708 47860 1720
rect 47912 1708 47918 1760
rect 10686 1640 10692 1692
rect 10744 1680 10750 1692
rect 12802 1680 12808 1692
rect 10744 1652 12808 1680
rect 10744 1640 10750 1652
rect 12802 1640 12808 1652
rect 12860 1640 12866 1692
rect 48958 1572 48964 1624
rect 49016 1612 49022 1624
rect 52362 1612 52368 1624
rect 49016 1584 52368 1612
rect 49016 1572 49022 1584
rect 52362 1572 52368 1584
rect 52420 1572 52426 1624
rect 13906 1368 13912 1420
rect 13964 1408 13970 1420
rect 14642 1408 14648 1420
rect 13964 1380 14648 1408
rect 13964 1368 13970 1380
rect 14642 1368 14648 1380
rect 14700 1368 14706 1420
rect 17678 1408 17684 1420
rect 14752 1380 17684 1408
rect 14752 1340 14780 1380
rect 17678 1368 17684 1380
rect 17736 1368 17742 1420
rect 14660 1312 14780 1340
rect 11606 1164 11612 1216
rect 11664 1204 11670 1216
rect 14182 1204 14188 1216
rect 11664 1176 14188 1204
rect 11664 1164 11670 1176
rect 14182 1164 14188 1176
rect 14240 1164 14246 1216
rect 14660 1068 14688 1312
rect 15010 1164 15016 1216
rect 15068 1204 15074 1216
rect 15068 1176 15148 1204
rect 15068 1164 15074 1176
rect 14734 1096 14740 1148
rect 14792 1136 14798 1148
rect 14792 1108 15056 1136
rect 14792 1096 14798 1108
rect 14660 1040 14780 1068
rect 14752 944 14780 1040
rect 15028 944 15056 1108
rect 15120 944 15148 1176
rect 14734 892 14740 944
rect 14792 892 14798 944
rect 15010 892 15016 944
rect 15068 892 15074 944
rect 15102 892 15108 944
rect 15160 892 15166 944
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 4344 57443 4396 57452
rect 4344 57409 4353 57443
rect 4353 57409 4387 57443
rect 4387 57409 4396 57443
rect 4344 57400 4396 57409
rect 4896 57400 4948 57452
rect 6000 57400 6052 57452
rect 6552 57400 6604 57452
rect 7656 57400 7708 57452
rect 8208 57443 8260 57452
rect 8208 57409 8217 57443
rect 8217 57409 8251 57443
rect 8251 57409 8260 57443
rect 8208 57400 8260 57409
rect 9312 57443 9364 57452
rect 9312 57409 9321 57443
rect 9321 57409 9355 57443
rect 9355 57409 9364 57443
rect 9312 57400 9364 57409
rect 9864 57400 9916 57452
rect 10968 57443 11020 57452
rect 10968 57409 10977 57443
rect 10977 57409 11011 57443
rect 11011 57409 11020 57443
rect 10968 57400 11020 57409
rect 11520 57400 11572 57452
rect 12624 57443 12676 57452
rect 12624 57409 12633 57443
rect 12633 57409 12667 57443
rect 12667 57409 12676 57443
rect 12624 57400 12676 57409
rect 13176 57400 13228 57452
rect 14280 57443 14332 57452
rect 14280 57409 14289 57443
rect 14289 57409 14323 57443
rect 14323 57409 14332 57443
rect 14280 57400 14332 57409
rect 14832 57400 14884 57452
rect 15936 57443 15988 57452
rect 15936 57409 15945 57443
rect 15945 57409 15979 57443
rect 15979 57409 15988 57443
rect 15936 57400 15988 57409
rect 17592 57443 17644 57452
rect 17592 57409 17601 57443
rect 17601 57409 17635 57443
rect 17635 57409 17644 57443
rect 17592 57400 17644 57409
rect 18144 57400 18196 57452
rect 19248 57443 19300 57452
rect 19248 57409 19257 57443
rect 19257 57409 19291 57443
rect 19291 57409 19300 57443
rect 19248 57400 19300 57409
rect 19984 57400 20036 57452
rect 20904 57400 20956 57452
rect 21456 57400 21508 57452
rect 22560 57443 22612 57452
rect 22560 57409 22569 57443
rect 22569 57409 22603 57443
rect 22603 57409 22612 57443
rect 22560 57400 22612 57409
rect 23112 57400 23164 57452
rect 24860 57443 24912 57452
rect 24860 57409 24869 57443
rect 24869 57409 24903 57443
rect 24903 57409 24912 57443
rect 24860 57400 24912 57409
rect 25872 57400 25924 57452
rect 26424 57443 26476 57452
rect 26424 57409 26433 57443
rect 26433 57409 26467 57443
rect 26467 57409 26476 57443
rect 26424 57400 26476 57409
rect 27528 57443 27580 57452
rect 27528 57409 27537 57443
rect 27537 57409 27571 57443
rect 27571 57409 27580 57443
rect 27528 57400 27580 57409
rect 28080 57400 28132 57452
rect 29184 57400 29236 57452
rect 29736 57400 29788 57452
rect 30840 57400 30892 57452
rect 31392 57443 31444 57452
rect 31392 57409 31401 57443
rect 31401 57409 31435 57443
rect 31435 57409 31444 57443
rect 31392 57400 31444 57409
rect 32496 57443 32548 57452
rect 32496 57409 32505 57443
rect 32505 57409 32539 57443
rect 32539 57409 32548 57443
rect 32496 57400 32548 57409
rect 33140 57443 33192 57452
rect 33140 57409 33149 57443
rect 33149 57409 33183 57443
rect 33183 57409 33192 57443
rect 33140 57400 33192 57409
rect 34152 57443 34204 57452
rect 34152 57409 34161 57443
rect 34161 57409 34195 57443
rect 34195 57409 34204 57443
rect 34152 57400 34204 57409
rect 34704 57400 34756 57452
rect 36360 57400 36412 57452
rect 37464 57400 37516 57452
rect 38016 57400 38068 57452
rect 39120 57400 39172 57452
rect 40040 57400 40092 57452
rect 40776 57400 40828 57452
rect 42432 57400 42484 57452
rect 42984 57400 43036 57452
rect 44180 57443 44232 57452
rect 44180 57409 44189 57443
rect 44189 57409 44223 57443
rect 44223 57409 44232 57443
rect 44180 57400 44232 57409
rect 44640 57400 44692 57452
rect 45744 57400 45796 57452
rect 46296 57400 46348 57452
rect 47400 57400 47452 57452
rect 47952 57400 48004 57452
rect 49056 57400 49108 57452
rect 49700 57400 49752 57452
rect 50712 57400 50764 57452
rect 51264 57400 51316 57452
rect 52460 57400 52512 57452
rect 52920 57400 52972 57452
rect 54024 57400 54076 57452
rect 55680 57400 55732 57452
rect 56600 57443 56652 57452
rect 56600 57409 56609 57443
rect 56609 57409 56643 57443
rect 56643 57409 56652 57443
rect 56600 57400 56652 57409
rect 57336 57400 57388 57452
rect 57980 57400 58032 57452
rect 58992 57400 59044 57452
rect 59544 57400 59596 57452
rect 60740 57400 60792 57452
rect 61200 57400 61252 57452
rect 62304 57400 62356 57452
rect 63960 57400 64012 57452
rect 65616 57400 65668 57452
rect 66260 57400 66312 57452
rect 16488 57332 16540 57384
rect 35808 57332 35860 57384
rect 62856 57332 62908 57384
rect 54576 57264 54628 57316
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 65654 57094 65706 57146
rect 65718 57094 65770 57146
rect 65782 57094 65834 57146
rect 65846 57094 65898 57146
rect 65910 57094 65962 57146
rect 24216 56992 24268 57044
rect 41420 57035 41472 57044
rect 41420 57001 41429 57035
rect 41429 57001 41463 57035
rect 41463 57001 41472 57035
rect 41420 56992 41472 57001
rect 64512 56992 64564 57044
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 67364 56355 67416 56364
rect 67364 56321 67373 56355
rect 67373 56321 67407 56355
rect 67407 56321 67416 56355
rect 67364 56312 67416 56321
rect 67548 56151 67600 56160
rect 67548 56117 67557 56151
rect 67557 56117 67591 56151
rect 67591 56117 67600 56151
rect 67548 56108 67600 56117
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 65654 56006 65706 56058
rect 65718 56006 65770 56058
rect 65782 56006 65834 56058
rect 65846 56006 65898 56058
rect 65910 56006 65962 56058
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 65654 54918 65706 54970
rect 65718 54918 65770 54970
rect 65782 54918 65834 54970
rect 65846 54918 65898 54970
rect 65910 54918 65962 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 65654 53830 65706 53882
rect 65718 53830 65770 53882
rect 65782 53830 65834 53882
rect 65846 53830 65898 53882
rect 65910 53830 65962 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 65654 52742 65706 52794
rect 65718 52742 65770 52794
rect 65782 52742 65834 52794
rect 65846 52742 65898 52794
rect 65910 52742 65962 52794
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 65654 51654 65706 51706
rect 65718 51654 65770 51706
rect 65782 51654 65834 51706
rect 65846 51654 65898 51706
rect 65910 51654 65962 51706
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 65654 50566 65706 50618
rect 65718 50566 65770 50618
rect 65782 50566 65834 50618
rect 65846 50566 65898 50618
rect 65910 50566 65962 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 65654 49478 65706 49530
rect 65718 49478 65770 49530
rect 65782 49478 65834 49530
rect 65846 49478 65898 49530
rect 65910 49478 65962 49530
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 67456 48696 67508 48748
rect 67548 48603 67600 48612
rect 67548 48569 67557 48603
rect 67557 48569 67591 48603
rect 67591 48569 67600 48603
rect 67548 48560 67600 48569
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 65654 48390 65706 48442
rect 65718 48390 65770 48442
rect 65782 48390 65834 48442
rect 65846 48390 65898 48442
rect 65910 48390 65962 48442
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 65654 47302 65706 47354
rect 65718 47302 65770 47354
rect 65782 47302 65834 47354
rect 65846 47302 65898 47354
rect 65910 47302 65962 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 65654 46214 65706 46266
rect 65718 46214 65770 46266
rect 65782 46214 65834 46266
rect 65846 46214 65898 46266
rect 65910 46214 65962 46266
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 43996 45432 44048 45484
rect 67364 45339 67416 45348
rect 67364 45305 67373 45339
rect 67373 45305 67407 45339
rect 67407 45305 67416 45339
rect 67364 45296 67416 45305
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 65654 45126 65706 45178
rect 65718 45126 65770 45178
rect 65782 45126 65834 45178
rect 65846 45126 65898 45178
rect 65910 45126 65962 45178
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 65654 44038 65706 44090
rect 65718 44038 65770 44090
rect 65782 44038 65834 44090
rect 65846 44038 65898 44090
rect 65910 44038 65962 44090
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 65654 42950 65706 43002
rect 65718 42950 65770 43002
rect 65782 42950 65834 43002
rect 65846 42950 65898 43002
rect 65910 42950 65962 43002
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 65654 41862 65706 41914
rect 65718 41862 65770 41914
rect 65782 41862 65834 41914
rect 65846 41862 65898 41914
rect 65910 41862 65962 41914
rect 67272 41463 67324 41472
rect 67272 41429 67281 41463
rect 67281 41429 67315 41463
rect 67315 41429 67324 41463
rect 67272 41420 67324 41429
rect 68008 41463 68060 41472
rect 68008 41429 68017 41463
rect 68017 41429 68051 41463
rect 68051 41429 68060 41463
rect 68008 41420 68060 41429
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 65654 40774 65706 40826
rect 65718 40774 65770 40826
rect 65782 40774 65834 40826
rect 65846 40774 65898 40826
rect 65910 40774 65962 40826
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 65654 39686 65706 39738
rect 65718 39686 65770 39738
rect 65782 39686 65834 39738
rect 65846 39686 65898 39738
rect 65910 39686 65962 39738
rect 67456 39584 67508 39636
rect 67180 39423 67232 39432
rect 67180 39389 67189 39423
rect 67189 39389 67223 39423
rect 67223 39389 67232 39423
rect 67180 39380 67232 39389
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 65654 38598 65706 38650
rect 65718 38598 65770 38650
rect 65782 38598 65834 38650
rect 65846 38598 65898 38650
rect 65910 38598 65962 38650
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 65654 37510 65706 37562
rect 65718 37510 65770 37562
rect 65782 37510 65834 37562
rect 65846 37510 65898 37562
rect 65910 37510 65962 37562
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 65654 36422 65706 36474
rect 65718 36422 65770 36474
rect 65782 36422 65834 36474
rect 65846 36422 65898 36474
rect 65910 36422 65962 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 65654 35334 65706 35386
rect 65718 35334 65770 35386
rect 65782 35334 65834 35386
rect 65846 35334 65898 35386
rect 65910 35334 65962 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 27620 34391 27672 34400
rect 27620 34357 27629 34391
rect 27629 34357 27663 34391
rect 27663 34357 27672 34391
rect 27620 34348 27672 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 65654 34246 65706 34298
rect 65718 34246 65770 34298
rect 65782 34246 65834 34298
rect 65846 34246 65898 34298
rect 65910 34246 65962 34298
rect 26884 34076 26936 34128
rect 29092 34076 29144 34128
rect 27252 34008 27304 34060
rect 27896 34008 27948 34060
rect 29000 34008 29052 34060
rect 26884 33940 26936 33992
rect 27068 33872 27120 33924
rect 67364 33940 67416 33992
rect 12900 33804 12952 33856
rect 27436 33804 27488 33856
rect 27620 33804 27672 33856
rect 28172 33804 28224 33856
rect 28816 33847 28868 33856
rect 28816 33813 28825 33847
rect 28825 33813 28859 33847
rect 28859 33813 28868 33847
rect 28816 33804 28868 33813
rect 68008 33847 68060 33856
rect 68008 33813 68017 33847
rect 68017 33813 68051 33847
rect 68051 33813 68060 33847
rect 68008 33804 68060 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 13176 33643 13228 33652
rect 13176 33609 13185 33643
rect 13185 33609 13219 33643
rect 13219 33609 13228 33643
rect 13176 33600 13228 33609
rect 7472 33464 7524 33516
rect 14280 33532 14332 33584
rect 13268 33507 13320 33516
rect 13268 33473 13277 33507
rect 13277 33473 13311 33507
rect 13311 33473 13320 33507
rect 13268 33464 13320 33473
rect 12532 33396 12584 33448
rect 16212 33464 16264 33516
rect 22192 33464 22244 33516
rect 31208 33600 31260 33652
rect 28172 33575 28224 33584
rect 28172 33541 28181 33575
rect 28181 33541 28215 33575
rect 28215 33541 28224 33575
rect 28908 33575 28960 33584
rect 28172 33532 28224 33541
rect 28908 33541 28917 33575
rect 28917 33541 28951 33575
rect 28951 33541 28960 33575
rect 28908 33532 28960 33541
rect 25964 33507 26016 33516
rect 25964 33473 25973 33507
rect 25973 33473 26007 33507
rect 26007 33473 26016 33507
rect 25964 33464 26016 33473
rect 9772 33328 9824 33380
rect 13176 33328 13228 33380
rect 23664 33396 23716 33448
rect 27712 33464 27764 33516
rect 27897 33464 27949 33516
rect 28080 33507 28132 33516
rect 28080 33473 28089 33507
rect 28089 33473 28123 33507
rect 28123 33473 28132 33507
rect 28080 33464 28132 33473
rect 27068 33396 27120 33448
rect 28448 33464 28500 33516
rect 29092 33507 29144 33516
rect 29092 33473 29101 33507
rect 29101 33473 29135 33507
rect 29135 33473 29144 33507
rect 32404 33600 32456 33652
rect 29092 33464 29144 33473
rect 34520 33464 34572 33516
rect 35348 33507 35400 33516
rect 35348 33473 35357 33507
rect 35357 33473 35391 33507
rect 35391 33473 35400 33507
rect 35348 33464 35400 33473
rect 26332 33371 26384 33380
rect 26332 33337 26341 33371
rect 26341 33337 26375 33371
rect 26375 33337 26384 33371
rect 26332 33328 26384 33337
rect 28080 33328 28132 33380
rect 28264 33328 28316 33380
rect 11152 33260 11204 33312
rect 14096 33303 14148 33312
rect 14096 33269 14105 33303
rect 14105 33269 14139 33303
rect 14139 33269 14148 33303
rect 14096 33260 14148 33269
rect 16028 33260 16080 33312
rect 26056 33260 26108 33312
rect 28816 33396 28868 33448
rect 37740 33396 37792 33448
rect 31116 33328 31168 33380
rect 31208 33328 31260 33380
rect 35900 33371 35952 33380
rect 35900 33337 35909 33371
rect 35909 33337 35943 33371
rect 35943 33337 35952 33371
rect 35900 33328 35952 33337
rect 34520 33260 34572 33312
rect 37188 33260 37240 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 65654 33158 65706 33210
rect 65718 33158 65770 33210
rect 65782 33158 65834 33210
rect 65846 33158 65898 33210
rect 65910 33158 65962 33210
rect 16212 33099 16264 33108
rect 16212 33065 16221 33099
rect 16221 33065 16255 33099
rect 16255 33065 16264 33099
rect 16212 33056 16264 33065
rect 26056 33099 26108 33108
rect 26056 33065 26065 33099
rect 26065 33065 26099 33099
rect 26099 33065 26108 33099
rect 26056 33056 26108 33065
rect 27068 33056 27120 33108
rect 12532 33031 12584 33040
rect 12532 32997 12541 33031
rect 12541 32997 12575 33031
rect 12575 32997 12584 33031
rect 12532 32988 12584 32997
rect 12900 32988 12952 33040
rect 19340 33031 19392 33040
rect 9772 32963 9824 32972
rect 9772 32929 9781 32963
rect 9781 32929 9815 32963
rect 9815 32929 9824 32963
rect 9772 32920 9824 32929
rect 12992 32963 13044 32972
rect 12992 32929 13001 32963
rect 13001 32929 13035 32963
rect 13035 32929 13044 32963
rect 12992 32920 13044 32929
rect 11152 32852 11204 32904
rect 12900 32895 12952 32904
rect 12900 32861 12909 32895
rect 12909 32861 12943 32895
rect 12943 32861 12952 32895
rect 12900 32852 12952 32861
rect 14280 32895 14332 32904
rect 14280 32861 14289 32895
rect 14289 32861 14323 32895
rect 14323 32861 14332 32895
rect 14280 32852 14332 32861
rect 14464 32895 14516 32904
rect 14464 32861 14473 32895
rect 14473 32861 14507 32895
rect 14507 32861 14516 32895
rect 14464 32852 14516 32861
rect 15016 32895 15068 32904
rect 15016 32861 15025 32895
rect 15025 32861 15059 32895
rect 15059 32861 15068 32895
rect 15016 32852 15068 32861
rect 16396 32895 16448 32904
rect 16396 32861 16405 32895
rect 16405 32861 16439 32895
rect 16439 32861 16448 32895
rect 16396 32852 16448 32861
rect 16028 32784 16080 32836
rect 19340 32997 19349 33031
rect 19349 32997 19383 33031
rect 19383 32997 19392 33031
rect 19340 32988 19392 32997
rect 19340 32852 19392 32904
rect 22192 32895 22244 32904
rect 22192 32861 22201 32895
rect 22201 32861 22235 32895
rect 22235 32861 22244 32895
rect 22192 32852 22244 32861
rect 10232 32716 10284 32768
rect 13820 32716 13872 32768
rect 15016 32716 15068 32768
rect 18236 32759 18288 32768
rect 18236 32725 18245 32759
rect 18245 32725 18279 32759
rect 18279 32725 18288 32759
rect 18236 32716 18288 32725
rect 20168 32716 20220 32768
rect 26332 32920 26384 32972
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 23664 32784 23716 32836
rect 26792 32895 26844 32904
rect 26792 32861 26801 32895
rect 26801 32861 26835 32895
rect 26835 32861 26844 32895
rect 26792 32852 26844 32861
rect 27436 32895 27488 32904
rect 27436 32861 27445 32895
rect 27445 32861 27479 32895
rect 27479 32861 27488 32895
rect 27436 32852 27488 32861
rect 33140 32920 33192 32972
rect 36544 32920 36596 32972
rect 38660 32920 38712 32972
rect 28356 32895 28408 32904
rect 28356 32861 28365 32895
rect 28365 32861 28399 32895
rect 28399 32861 28408 32895
rect 28356 32852 28408 32861
rect 28632 32895 28684 32904
rect 28632 32861 28641 32895
rect 28641 32861 28675 32895
rect 28675 32861 28684 32895
rect 28632 32852 28684 32861
rect 29000 32852 29052 32904
rect 29736 32895 29788 32904
rect 29736 32861 29745 32895
rect 29745 32861 29779 32895
rect 29779 32861 29788 32895
rect 29736 32852 29788 32861
rect 32404 32895 32456 32904
rect 32404 32861 32413 32895
rect 32413 32861 32447 32895
rect 32447 32861 32456 32895
rect 32404 32852 32456 32861
rect 35348 32852 35400 32904
rect 35900 32852 35952 32904
rect 37188 32895 37240 32904
rect 37188 32861 37197 32895
rect 37197 32861 37231 32895
rect 37231 32861 37240 32895
rect 37188 32852 37240 32861
rect 38292 32895 38344 32904
rect 26424 32716 26476 32768
rect 33324 32716 33376 32768
rect 38292 32861 38301 32895
rect 38301 32861 38335 32895
rect 38335 32861 38344 32895
rect 38292 32852 38344 32861
rect 38752 32716 38804 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 18236 32512 18288 32564
rect 26792 32512 26844 32564
rect 28632 32555 28684 32564
rect 28632 32521 28641 32555
rect 28641 32521 28675 32555
rect 28675 32521 28684 32555
rect 28632 32512 28684 32521
rect 34520 32512 34572 32564
rect 38660 32555 38712 32564
rect 38660 32521 38669 32555
rect 38669 32521 38703 32555
rect 38703 32521 38712 32555
rect 38660 32512 38712 32521
rect 7104 32376 7156 32428
rect 9036 32419 9088 32428
rect 9036 32385 9045 32419
rect 9045 32385 9079 32419
rect 9079 32385 9088 32419
rect 9036 32376 9088 32385
rect 13176 32376 13228 32428
rect 13820 32419 13872 32428
rect 13820 32385 13829 32419
rect 13829 32385 13863 32419
rect 13863 32385 13872 32419
rect 13820 32376 13872 32385
rect 12808 32351 12860 32360
rect 12808 32317 12817 32351
rect 12817 32317 12851 32351
rect 12851 32317 12860 32351
rect 12808 32308 12860 32317
rect 13268 32308 13320 32360
rect 14096 32419 14148 32428
rect 14096 32385 14105 32419
rect 14105 32385 14139 32419
rect 14139 32385 14148 32419
rect 14096 32376 14148 32385
rect 14464 32376 14516 32428
rect 15476 32419 15528 32428
rect 15476 32385 15485 32419
rect 15485 32385 15519 32419
rect 15519 32385 15528 32419
rect 15476 32376 15528 32385
rect 16028 32419 16080 32428
rect 16028 32385 16037 32419
rect 16037 32385 16071 32419
rect 16071 32385 16080 32419
rect 16028 32376 16080 32385
rect 14740 32308 14792 32360
rect 17408 32308 17460 32360
rect 18696 32376 18748 32428
rect 23204 32419 23256 32428
rect 23204 32385 23213 32419
rect 23213 32385 23247 32419
rect 23247 32385 23256 32419
rect 23204 32376 23256 32385
rect 23388 32376 23440 32428
rect 25320 32419 25372 32428
rect 25320 32385 25329 32419
rect 25329 32385 25363 32419
rect 25363 32385 25372 32419
rect 25320 32376 25372 32385
rect 35348 32444 35400 32496
rect 26424 32419 26476 32428
rect 26424 32385 26433 32419
rect 26433 32385 26467 32419
rect 26467 32385 26476 32419
rect 26424 32376 26476 32385
rect 27896 32376 27948 32428
rect 29000 32419 29052 32428
rect 28724 32308 28776 32360
rect 29000 32385 29009 32419
rect 29009 32385 29043 32419
rect 29043 32385 29052 32419
rect 29000 32376 29052 32385
rect 34520 32419 34572 32428
rect 29736 32308 29788 32360
rect 27620 32283 27672 32292
rect 27620 32249 27629 32283
rect 27629 32249 27663 32283
rect 27663 32249 27672 32283
rect 27620 32240 27672 32249
rect 34520 32385 34529 32419
rect 34529 32385 34563 32419
rect 34563 32385 34572 32419
rect 34520 32376 34572 32385
rect 35808 32376 35860 32428
rect 36544 32419 36596 32428
rect 36544 32385 36553 32419
rect 36553 32385 36587 32419
rect 36587 32385 36596 32419
rect 36544 32376 36596 32385
rect 37188 32376 37240 32428
rect 37740 32419 37792 32428
rect 37740 32385 37749 32419
rect 37749 32385 37783 32419
rect 37783 32385 37792 32419
rect 37740 32376 37792 32385
rect 35532 32351 35584 32360
rect 35532 32317 35541 32351
rect 35541 32317 35575 32351
rect 35575 32317 35584 32351
rect 35532 32308 35584 32317
rect 37648 32283 37700 32292
rect 37648 32249 37657 32283
rect 37657 32249 37691 32283
rect 37691 32249 37700 32283
rect 37648 32240 37700 32249
rect 40500 32308 40552 32360
rect 6368 32215 6420 32224
rect 6368 32181 6377 32215
rect 6377 32181 6411 32215
rect 6411 32181 6420 32215
rect 6368 32172 6420 32181
rect 9680 32172 9732 32224
rect 14280 32172 14332 32224
rect 15292 32215 15344 32224
rect 15292 32181 15301 32215
rect 15301 32181 15335 32215
rect 15335 32181 15344 32215
rect 15292 32172 15344 32181
rect 17592 32172 17644 32224
rect 22744 32172 22796 32224
rect 33968 32172 34020 32224
rect 35900 32172 35952 32224
rect 37280 32215 37332 32224
rect 37280 32181 37289 32215
rect 37289 32181 37323 32215
rect 37323 32181 37332 32215
rect 37280 32172 37332 32181
rect 37464 32172 37516 32224
rect 40040 32172 40092 32224
rect 41144 32172 41196 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 65654 32070 65706 32122
rect 65718 32070 65770 32122
rect 65782 32070 65834 32122
rect 65846 32070 65898 32122
rect 65910 32070 65962 32122
rect 7104 32011 7156 32020
rect 7104 31977 7113 32011
rect 7113 31977 7147 32011
rect 7147 31977 7156 32011
rect 7104 31968 7156 31977
rect 7012 31832 7064 31884
rect 5264 31807 5316 31816
rect 5264 31773 5273 31807
rect 5273 31773 5307 31807
rect 5307 31773 5316 31807
rect 5264 31764 5316 31773
rect 7288 31764 7340 31816
rect 12992 31968 13044 32020
rect 13636 31968 13688 32020
rect 14464 31968 14516 32020
rect 16396 32011 16448 32020
rect 16396 31977 16405 32011
rect 16405 31977 16439 32011
rect 16439 31977 16448 32011
rect 16396 31968 16448 31977
rect 19340 32011 19392 32020
rect 19340 31977 19349 32011
rect 19349 31977 19383 32011
rect 19383 31977 19392 32011
rect 19340 31968 19392 31977
rect 22284 31968 22336 32020
rect 23388 31968 23440 32020
rect 25964 31968 26016 32020
rect 27620 31968 27672 32020
rect 16580 31900 16632 31952
rect 12072 31764 12124 31816
rect 13636 31764 13688 31816
rect 18144 31764 18196 31816
rect 23664 31900 23716 31952
rect 36544 31968 36596 32020
rect 27896 31875 27948 31884
rect 19156 31764 19208 31816
rect 20628 31807 20680 31816
rect 20628 31773 20637 31807
rect 20637 31773 20671 31807
rect 20671 31773 20680 31807
rect 20628 31764 20680 31773
rect 5540 31739 5592 31748
rect 5540 31705 5574 31739
rect 5574 31705 5592 31739
rect 5540 31696 5592 31705
rect 12624 31696 12676 31748
rect 15292 31739 15344 31748
rect 15292 31705 15326 31739
rect 15326 31705 15344 31739
rect 15292 31696 15344 31705
rect 15384 31696 15436 31748
rect 17592 31739 17644 31748
rect 17592 31705 17626 31739
rect 17626 31705 17644 31739
rect 17592 31696 17644 31705
rect 20996 31696 21048 31748
rect 22744 31739 22796 31748
rect 22744 31705 22778 31739
rect 22778 31705 22796 31739
rect 22744 31696 22796 31705
rect 24308 31696 24360 31748
rect 24492 31696 24544 31748
rect 27436 31696 27488 31748
rect 27896 31841 27905 31875
rect 27905 31841 27939 31875
rect 27939 31841 27948 31875
rect 27896 31832 27948 31841
rect 36452 31900 36504 31952
rect 34704 31807 34756 31816
rect 34704 31773 34713 31807
rect 34713 31773 34747 31807
rect 34747 31773 34756 31807
rect 34704 31764 34756 31773
rect 37280 31807 37332 31816
rect 37280 31773 37289 31807
rect 37289 31773 37323 31807
rect 37323 31773 37332 31807
rect 37280 31764 37332 31773
rect 37464 31807 37516 31816
rect 37464 31773 37471 31807
rect 37471 31773 37516 31807
rect 37464 31764 37516 31773
rect 38660 31968 38712 32020
rect 38200 31900 38252 31952
rect 37648 31832 37700 31884
rect 38292 31832 38344 31884
rect 67272 31900 67324 31952
rect 41144 31875 41196 31884
rect 41144 31841 41153 31875
rect 41153 31841 41187 31875
rect 41187 31841 41196 31875
rect 41144 31832 41196 31841
rect 38568 31807 38620 31816
rect 38568 31773 38577 31807
rect 38577 31773 38611 31807
rect 38611 31773 38620 31807
rect 38568 31764 38620 31773
rect 40040 31807 40092 31816
rect 40040 31773 40049 31807
rect 40049 31773 40083 31807
rect 40083 31773 40092 31807
rect 40040 31764 40092 31773
rect 41236 31807 41288 31816
rect 41236 31773 41245 31807
rect 41245 31773 41279 31807
rect 41279 31773 41288 31807
rect 41236 31764 41288 31773
rect 41880 31807 41932 31816
rect 41880 31773 41889 31807
rect 41889 31773 41923 31807
rect 41923 31773 41932 31807
rect 41880 31764 41932 31773
rect 57704 31807 57756 31816
rect 57704 31773 57713 31807
rect 57713 31773 57747 31807
rect 57747 31773 57756 31807
rect 57704 31764 57756 31773
rect 31484 31739 31536 31748
rect 31484 31705 31518 31739
rect 31518 31705 31536 31739
rect 31484 31696 31536 31705
rect 35716 31696 35768 31748
rect 36452 31696 36504 31748
rect 5632 31628 5684 31680
rect 6460 31628 6512 31680
rect 7472 31671 7524 31680
rect 7472 31637 7481 31671
rect 7481 31637 7515 31671
rect 7515 31637 7524 31671
rect 7472 31628 7524 31637
rect 19984 31671 20036 31680
rect 19984 31637 19993 31671
rect 19993 31637 20027 31671
rect 20027 31637 20036 31671
rect 19984 31628 20036 31637
rect 22192 31628 22244 31680
rect 28448 31628 28500 31680
rect 28816 31671 28868 31680
rect 28816 31637 28825 31671
rect 28825 31637 28859 31671
rect 28859 31637 28868 31671
rect 28816 31628 28868 31637
rect 32312 31628 32364 31680
rect 34520 31628 34572 31680
rect 35808 31628 35860 31680
rect 40408 31671 40460 31680
rect 40408 31637 40417 31671
rect 40417 31637 40451 31671
rect 40451 31637 40460 31671
rect 40408 31628 40460 31637
rect 40868 31671 40920 31680
rect 40868 31637 40877 31671
rect 40877 31637 40911 31671
rect 40911 31637 40920 31671
rect 40868 31628 40920 31637
rect 42064 31671 42116 31680
rect 42064 31637 42073 31671
rect 42073 31637 42107 31671
rect 42107 31637 42116 31671
rect 42064 31628 42116 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 5632 31424 5684 31476
rect 7104 31424 7156 31476
rect 12624 31467 12676 31476
rect 12624 31433 12633 31467
rect 12633 31433 12667 31467
rect 12667 31433 12676 31467
rect 12624 31424 12676 31433
rect 13636 31467 13688 31476
rect 6460 31288 6512 31340
rect 8392 31331 8444 31340
rect 8392 31297 8401 31331
rect 8401 31297 8435 31331
rect 8435 31297 8444 31331
rect 8392 31288 8444 31297
rect 9772 31288 9824 31340
rect 9956 31331 10008 31340
rect 9956 31297 9965 31331
rect 9965 31297 9999 31331
rect 9999 31297 10008 31331
rect 9956 31288 10008 31297
rect 10232 31331 10284 31340
rect 10232 31297 10241 31331
rect 10241 31297 10275 31331
rect 10275 31297 10284 31331
rect 10232 31288 10284 31297
rect 13636 31433 13645 31467
rect 13645 31433 13679 31467
rect 13679 31433 13688 31467
rect 13636 31424 13688 31433
rect 15476 31424 15528 31476
rect 16396 31424 16448 31476
rect 17224 31424 17276 31476
rect 17408 31424 17460 31476
rect 20168 31424 20220 31476
rect 20996 31467 21048 31476
rect 20996 31433 21005 31467
rect 21005 31433 21039 31467
rect 21039 31433 21048 31467
rect 20996 31424 21048 31433
rect 22284 31467 22336 31476
rect 5172 31084 5224 31136
rect 5448 31152 5500 31204
rect 8300 31152 8352 31204
rect 9036 31152 9088 31204
rect 13728 31263 13780 31272
rect 13728 31229 13737 31263
rect 13737 31229 13771 31263
rect 13771 31229 13780 31263
rect 13728 31220 13780 31229
rect 13820 31263 13872 31272
rect 13820 31229 13829 31263
rect 13829 31229 13863 31263
rect 13863 31229 13872 31263
rect 13820 31220 13872 31229
rect 14924 31220 14976 31272
rect 17040 31288 17092 31340
rect 18236 31288 18288 31340
rect 18420 31331 18472 31340
rect 18420 31297 18454 31331
rect 18454 31297 18472 31331
rect 18420 31288 18472 31297
rect 18972 31288 19024 31340
rect 19984 31288 20036 31340
rect 22284 31433 22293 31467
rect 22293 31433 22327 31467
rect 22327 31433 22336 31467
rect 22284 31424 22336 31433
rect 23204 31467 23256 31476
rect 23204 31433 23213 31467
rect 23213 31433 23247 31467
rect 23247 31433 23256 31467
rect 23204 31424 23256 31433
rect 23664 31467 23716 31476
rect 23664 31433 23673 31467
rect 23673 31433 23707 31467
rect 23707 31433 23716 31467
rect 23664 31424 23716 31433
rect 24492 31467 24544 31476
rect 24492 31433 24501 31467
rect 24501 31433 24535 31467
rect 24535 31433 24544 31467
rect 24492 31424 24544 31433
rect 22192 31399 22244 31408
rect 17132 31263 17184 31272
rect 17132 31229 17141 31263
rect 17141 31229 17175 31263
rect 17175 31229 17184 31263
rect 17132 31220 17184 31229
rect 16948 31152 17000 31204
rect 22192 31365 22201 31399
rect 22201 31365 22235 31399
rect 22235 31365 22244 31399
rect 22192 31356 22244 31365
rect 22744 31220 22796 31272
rect 25964 31424 26016 31476
rect 28356 31424 28408 31476
rect 28448 31424 28500 31476
rect 29736 31467 29788 31476
rect 28816 31356 28868 31408
rect 29736 31433 29745 31467
rect 29745 31433 29779 31467
rect 29779 31433 29788 31467
rect 29736 31424 29788 31433
rect 31484 31424 31536 31476
rect 34520 31424 34572 31476
rect 25504 31331 25556 31340
rect 25504 31297 25513 31331
rect 25513 31297 25547 31331
rect 25547 31297 25556 31331
rect 25504 31288 25556 31297
rect 27160 31331 27212 31340
rect 27160 31297 27169 31331
rect 27169 31297 27203 31331
rect 27203 31297 27212 31331
rect 27160 31288 27212 31297
rect 25780 31220 25832 31272
rect 28356 31263 28408 31272
rect 28356 31229 28365 31263
rect 28365 31229 28399 31263
rect 28399 31229 28408 31263
rect 28356 31220 28408 31229
rect 27436 31152 27488 31204
rect 8484 31084 8536 31136
rect 9680 31084 9732 31136
rect 14188 31084 14240 31136
rect 14924 31127 14976 31136
rect 14924 31093 14933 31127
rect 14933 31093 14967 31127
rect 14967 31093 14976 31127
rect 14924 31084 14976 31093
rect 17316 31084 17368 31136
rect 32312 31220 32364 31272
rect 32680 31263 32732 31272
rect 32680 31229 32689 31263
rect 32689 31229 32723 31263
rect 32723 31229 32732 31263
rect 34704 31356 34756 31408
rect 35348 31424 35400 31476
rect 35716 31467 35768 31476
rect 35716 31433 35725 31467
rect 35725 31433 35759 31467
rect 35759 31433 35768 31467
rect 35716 31424 35768 31433
rect 41236 31424 41288 31476
rect 41880 31424 41932 31476
rect 33968 31288 34020 31340
rect 35900 31331 35952 31340
rect 35900 31297 35909 31331
rect 35909 31297 35943 31331
rect 35943 31297 35952 31331
rect 35900 31288 35952 31297
rect 37004 31288 37056 31340
rect 32680 31220 32732 31229
rect 31944 31152 31996 31204
rect 35992 31220 36044 31272
rect 42432 31331 42484 31340
rect 42432 31297 42441 31331
rect 42441 31297 42475 31331
rect 42475 31297 42484 31331
rect 42432 31288 42484 31297
rect 41512 31152 41564 31204
rect 37464 31084 37516 31136
rect 38568 31084 38620 31136
rect 43536 31084 43588 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 65654 30982 65706 31034
rect 65718 30982 65770 31034
rect 65782 30982 65834 31034
rect 65846 30982 65898 31034
rect 65910 30982 65962 31034
rect 5540 30880 5592 30932
rect 7472 30880 7524 30932
rect 8392 30923 8444 30932
rect 8392 30889 8401 30923
rect 8401 30889 8435 30923
rect 8435 30889 8444 30923
rect 8392 30880 8444 30889
rect 8484 30880 8536 30932
rect 15936 30880 15988 30932
rect 16580 30923 16632 30932
rect 16580 30889 16589 30923
rect 16589 30889 16623 30923
rect 16623 30889 16632 30923
rect 16580 30880 16632 30889
rect 18420 30880 18472 30932
rect 18696 30923 18748 30932
rect 18696 30889 18705 30923
rect 18705 30889 18739 30923
rect 18739 30889 18748 30923
rect 18696 30880 18748 30889
rect 17960 30812 18012 30864
rect 5080 30744 5132 30796
rect 5448 30744 5500 30796
rect 7104 30744 7156 30796
rect 5172 30719 5224 30728
rect 5172 30685 5181 30719
rect 5181 30685 5215 30719
rect 5215 30685 5224 30719
rect 5172 30676 5224 30685
rect 6368 30676 6420 30728
rect 8300 30676 8352 30728
rect 7932 30651 7984 30660
rect 7932 30617 7941 30651
rect 7941 30617 7975 30651
rect 7975 30617 7984 30651
rect 7932 30608 7984 30617
rect 11704 30608 11756 30660
rect 12072 30676 12124 30728
rect 15476 30719 15528 30728
rect 15476 30685 15485 30719
rect 15485 30685 15519 30719
rect 15519 30685 15528 30719
rect 15476 30676 15528 30685
rect 13728 30608 13780 30660
rect 16948 30608 17000 30660
rect 17132 30744 17184 30796
rect 20260 30744 20312 30796
rect 17316 30719 17368 30728
rect 17316 30685 17325 30719
rect 17325 30685 17359 30719
rect 17359 30685 17368 30719
rect 17316 30676 17368 30685
rect 20628 30719 20680 30728
rect 20628 30685 20637 30719
rect 20637 30685 20671 30719
rect 20671 30685 20680 30719
rect 20628 30676 20680 30685
rect 18052 30608 18104 30660
rect 19432 30608 19484 30660
rect 21088 30608 21140 30660
rect 22192 30880 22244 30932
rect 24400 30744 24452 30796
rect 27160 30812 27212 30864
rect 31300 30880 31352 30932
rect 32680 30880 32732 30932
rect 36452 30923 36504 30932
rect 36452 30889 36461 30923
rect 36461 30889 36495 30923
rect 36495 30889 36504 30923
rect 36452 30880 36504 30889
rect 37004 30923 37056 30932
rect 37004 30889 37013 30923
rect 37013 30889 37047 30923
rect 37047 30889 37056 30923
rect 37004 30880 37056 30889
rect 41236 30923 41288 30932
rect 41236 30889 41245 30923
rect 41245 30889 41279 30923
rect 41279 30889 41288 30923
rect 41236 30880 41288 30889
rect 37464 30787 37516 30796
rect 24676 30719 24728 30728
rect 24676 30685 24685 30719
rect 24685 30685 24719 30719
rect 24719 30685 24728 30719
rect 24676 30676 24728 30685
rect 25504 30676 25556 30728
rect 25964 30651 26016 30660
rect 25964 30617 25998 30651
rect 25998 30617 26016 30651
rect 27436 30676 27488 30728
rect 25964 30608 26016 30617
rect 29644 30608 29696 30660
rect 12164 30540 12216 30592
rect 15568 30540 15620 30592
rect 18144 30540 18196 30592
rect 19340 30540 19392 30592
rect 21916 30540 21968 30592
rect 24492 30583 24544 30592
rect 24492 30549 24501 30583
rect 24501 30549 24535 30583
rect 24535 30549 24544 30583
rect 24492 30540 24544 30549
rect 27528 30583 27580 30592
rect 27528 30549 27537 30583
rect 27537 30549 27571 30583
rect 27571 30549 27580 30583
rect 27528 30540 27580 30549
rect 27896 30583 27948 30592
rect 27896 30549 27905 30583
rect 27905 30549 27939 30583
rect 27939 30549 27948 30583
rect 27896 30540 27948 30549
rect 29000 30540 29052 30592
rect 31944 30719 31996 30728
rect 31944 30685 31953 30719
rect 31953 30685 31987 30719
rect 31987 30685 31996 30719
rect 31944 30676 31996 30685
rect 37464 30753 37473 30787
rect 37473 30753 37507 30787
rect 37507 30753 37516 30787
rect 37464 30744 37516 30753
rect 37280 30676 37332 30728
rect 42064 30676 42116 30728
rect 43812 30676 43864 30728
rect 32036 30608 32088 30660
rect 35808 30608 35860 30660
rect 32588 30540 32640 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 9772 30336 9824 30388
rect 11704 30379 11756 30388
rect 11704 30345 11713 30379
rect 11713 30345 11747 30379
rect 11747 30345 11756 30379
rect 11704 30336 11756 30345
rect 15476 30336 15528 30388
rect 18052 30379 18104 30388
rect 18052 30345 18061 30379
rect 18061 30345 18095 30379
rect 18095 30345 18104 30379
rect 21088 30379 21140 30388
rect 18052 30336 18104 30345
rect 17040 30268 17092 30320
rect 18144 30268 18196 30320
rect 18972 30268 19024 30320
rect 21088 30345 21097 30379
rect 21097 30345 21131 30379
rect 21131 30345 21140 30379
rect 21088 30336 21140 30345
rect 25964 30379 26016 30388
rect 25964 30345 25973 30379
rect 25973 30345 26007 30379
rect 26007 30345 26016 30379
rect 25964 30336 26016 30345
rect 32036 30336 32088 30388
rect 42432 30336 42484 30388
rect 20536 30268 20588 30320
rect 24492 30268 24544 30320
rect 27896 30268 27948 30320
rect 32588 30311 32640 30320
rect 11152 30200 11204 30252
rect 11796 30200 11848 30252
rect 16672 30200 16724 30252
rect 22192 30243 22244 30252
rect 11060 30132 11112 30184
rect 15844 30175 15896 30184
rect 15844 30141 15853 30175
rect 15853 30141 15887 30175
rect 15887 30141 15896 30175
rect 15844 30132 15896 30141
rect 13820 30064 13872 30116
rect 19432 30107 19484 30116
rect 19432 30073 19441 30107
rect 19441 30073 19475 30107
rect 19475 30073 19484 30107
rect 19432 30064 19484 30073
rect 22192 30209 22201 30243
rect 22201 30209 22235 30243
rect 22235 30209 22244 30243
rect 22192 30200 22244 30209
rect 21916 30132 21968 30184
rect 22744 30132 22796 30184
rect 27528 30200 27580 30252
rect 28356 30200 28408 30252
rect 28816 30200 28868 30252
rect 30840 30243 30892 30252
rect 30840 30209 30849 30243
rect 30849 30209 30883 30243
rect 30883 30209 30892 30243
rect 30840 30200 30892 30209
rect 32588 30277 32597 30311
rect 32597 30277 32631 30311
rect 32631 30277 32640 30311
rect 32588 30268 32640 30277
rect 43536 30311 43588 30320
rect 43536 30277 43554 30311
rect 43554 30277 43588 30311
rect 43536 30268 43588 30277
rect 32496 30243 32548 30252
rect 32496 30209 32505 30243
rect 32505 30209 32539 30243
rect 32539 30209 32548 30243
rect 32496 30200 32548 30209
rect 37280 30200 37332 30252
rect 40408 30243 40460 30252
rect 40408 30209 40417 30243
rect 40417 30209 40451 30243
rect 40451 30209 40460 30243
rect 40408 30200 40460 30209
rect 40684 30243 40736 30252
rect 40684 30209 40693 30243
rect 40693 30209 40727 30243
rect 40727 30209 40736 30243
rect 40684 30200 40736 30209
rect 40776 30200 40828 30252
rect 43812 30243 43864 30252
rect 43812 30209 43821 30243
rect 43821 30209 43855 30243
rect 43855 30209 43864 30243
rect 43812 30200 43864 30209
rect 16948 29996 17000 30048
rect 20076 30039 20128 30048
rect 20076 30005 20085 30039
rect 20085 30005 20119 30039
rect 20119 30005 20128 30039
rect 20076 29996 20128 30005
rect 27896 30132 27948 30184
rect 32680 30175 32732 30184
rect 32680 30141 32689 30175
rect 32689 30141 32723 30175
rect 32723 30141 32732 30175
rect 32680 30132 32732 30141
rect 40592 30175 40644 30184
rect 40592 30141 40601 30175
rect 40601 30141 40635 30175
rect 40635 30141 40644 30175
rect 40592 30132 40644 30141
rect 24400 29996 24452 30048
rect 24768 29996 24820 30048
rect 29644 30039 29696 30048
rect 29644 30005 29653 30039
rect 29653 30005 29687 30039
rect 29687 30005 29696 30039
rect 29644 29996 29696 30005
rect 30656 30039 30708 30048
rect 30656 30005 30665 30039
rect 30665 30005 30699 30039
rect 30699 30005 30708 30039
rect 30656 29996 30708 30005
rect 36360 29996 36412 30048
rect 40132 29996 40184 30048
rect 40868 29996 40920 30048
rect 41604 30064 41656 30116
rect 41512 29996 41564 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 65654 29894 65706 29946
rect 65718 29894 65770 29946
rect 65782 29894 65834 29946
rect 65846 29894 65898 29946
rect 65910 29894 65962 29946
rect 11796 29835 11848 29844
rect 11796 29801 11805 29835
rect 11805 29801 11839 29835
rect 11839 29801 11848 29835
rect 11796 29792 11848 29801
rect 16672 29835 16724 29844
rect 16672 29801 16681 29835
rect 16681 29801 16715 29835
rect 16715 29801 16724 29835
rect 16672 29792 16724 29801
rect 24676 29792 24728 29844
rect 28816 29835 28868 29844
rect 28816 29801 28825 29835
rect 28825 29801 28859 29835
rect 28859 29801 28868 29835
rect 28816 29792 28868 29801
rect 32496 29792 32548 29844
rect 37648 29792 37700 29844
rect 4988 29588 5040 29640
rect 7012 29699 7064 29708
rect 7012 29665 7021 29699
rect 7021 29665 7055 29699
rect 7055 29665 7064 29699
rect 7012 29656 7064 29665
rect 9956 29724 10008 29776
rect 40592 29792 40644 29844
rect 67364 29835 67416 29844
rect 67364 29801 67373 29835
rect 67373 29801 67407 29835
rect 67407 29801 67416 29835
rect 67364 29792 67416 29801
rect 40776 29724 40828 29776
rect 13820 29656 13872 29708
rect 27528 29656 27580 29708
rect 28356 29656 28408 29708
rect 30472 29699 30524 29708
rect 30472 29665 30481 29699
rect 30481 29665 30515 29699
rect 30515 29665 30524 29699
rect 30472 29656 30524 29665
rect 35992 29699 36044 29708
rect 35992 29665 36001 29699
rect 36001 29665 36035 29699
rect 36035 29665 36044 29699
rect 35992 29656 36044 29665
rect 41052 29656 41104 29708
rect 6736 29588 6788 29640
rect 9128 29631 9180 29640
rect 9128 29597 9137 29631
rect 9137 29597 9171 29631
rect 9171 29597 9180 29631
rect 9128 29588 9180 29597
rect 10968 29631 11020 29640
rect 10968 29597 10977 29631
rect 10977 29597 11011 29631
rect 11011 29597 11020 29631
rect 10968 29588 11020 29597
rect 11152 29631 11204 29640
rect 11152 29597 11161 29631
rect 11161 29597 11195 29631
rect 11195 29597 11204 29631
rect 11152 29588 11204 29597
rect 11796 29588 11848 29640
rect 5264 29520 5316 29572
rect 12164 29563 12216 29572
rect 12164 29529 12173 29563
rect 12173 29529 12207 29563
rect 12207 29529 12216 29563
rect 12164 29520 12216 29529
rect 15384 29588 15436 29640
rect 15568 29631 15620 29640
rect 15568 29597 15602 29631
rect 15602 29597 15620 29631
rect 15568 29588 15620 29597
rect 16672 29588 16724 29640
rect 18328 29588 18380 29640
rect 19248 29588 19300 29640
rect 22192 29588 22244 29640
rect 29000 29631 29052 29640
rect 29000 29597 29009 29631
rect 29009 29597 29043 29631
rect 29043 29597 29052 29631
rect 29000 29588 29052 29597
rect 20076 29520 20128 29572
rect 24768 29520 24820 29572
rect 30656 29520 30708 29572
rect 35900 29588 35952 29640
rect 41604 29631 41656 29640
rect 41604 29597 41613 29631
rect 41613 29597 41647 29631
rect 41647 29597 41656 29631
rect 41604 29588 41656 29597
rect 61384 29588 61436 29640
rect 11704 29452 11756 29504
rect 13912 29452 13964 29504
rect 15108 29452 15160 29504
rect 19432 29452 19484 29504
rect 23848 29495 23900 29504
rect 23848 29461 23857 29495
rect 23857 29461 23891 29495
rect 23891 29461 23900 29495
rect 23848 29452 23900 29461
rect 25412 29452 25464 29504
rect 31392 29452 31444 29504
rect 37372 29495 37424 29504
rect 37372 29461 37381 29495
rect 37381 29461 37415 29495
rect 37415 29461 37424 29495
rect 37372 29452 37424 29461
rect 38660 29452 38712 29504
rect 40960 29452 41012 29504
rect 42800 29452 42852 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 5264 29291 5316 29300
rect 5264 29257 5273 29291
rect 5273 29257 5307 29291
rect 5307 29257 5316 29291
rect 5264 29248 5316 29257
rect 6736 29291 6788 29300
rect 6736 29257 6745 29291
rect 6745 29257 6779 29291
rect 6779 29257 6788 29291
rect 6736 29248 6788 29257
rect 14004 29248 14056 29300
rect 14556 29248 14608 29300
rect 37280 29291 37332 29300
rect 6184 29180 6236 29232
rect 15936 29223 15988 29232
rect 7012 29112 7064 29164
rect 10324 29155 10376 29164
rect 10324 29121 10333 29155
rect 10333 29121 10367 29155
rect 10367 29121 10376 29155
rect 10324 29112 10376 29121
rect 11152 29112 11204 29164
rect 15936 29189 15945 29223
rect 15945 29189 15979 29223
rect 15979 29189 15988 29223
rect 15936 29180 15988 29189
rect 11704 29155 11756 29164
rect 11704 29121 11713 29155
rect 11713 29121 11747 29155
rect 11747 29121 11756 29155
rect 11704 29112 11756 29121
rect 12532 29155 12584 29164
rect 12532 29121 12541 29155
rect 12541 29121 12575 29155
rect 12575 29121 12584 29155
rect 12532 29112 12584 29121
rect 15108 29112 15160 29164
rect 15844 29112 15896 29164
rect 16672 29155 16724 29164
rect 16672 29121 16681 29155
rect 16681 29121 16715 29155
rect 16715 29121 16724 29155
rect 16672 29112 16724 29121
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 18236 29180 18288 29232
rect 16856 29112 16908 29121
rect 7104 29044 7156 29096
rect 9588 29044 9640 29096
rect 14280 29087 14332 29096
rect 11060 28976 11112 29028
rect 12440 28976 12492 29028
rect 14280 29053 14289 29087
rect 14289 29053 14323 29087
rect 14323 29053 14332 29087
rect 14280 29044 14332 29053
rect 19064 29112 19116 29164
rect 19432 29155 19484 29164
rect 30472 29180 30524 29232
rect 19432 29121 19450 29155
rect 19450 29121 19484 29155
rect 19432 29112 19484 29121
rect 20720 29112 20772 29164
rect 21732 29112 21784 29164
rect 22100 29155 22152 29164
rect 22100 29121 22109 29155
rect 22109 29121 22143 29155
rect 22143 29121 22152 29155
rect 24584 29155 24636 29164
rect 22100 29112 22152 29121
rect 24584 29121 24593 29155
rect 24593 29121 24627 29155
rect 24627 29121 24636 29155
rect 24584 29112 24636 29121
rect 31944 29180 31996 29232
rect 35348 29180 35400 29232
rect 37280 29257 37289 29291
rect 37289 29257 37323 29291
rect 37323 29257 37332 29291
rect 37280 29248 37332 29257
rect 37648 29291 37700 29300
rect 37648 29257 37657 29291
rect 37657 29257 37691 29291
rect 37691 29257 37700 29291
rect 37648 29248 37700 29257
rect 40684 29248 40736 29300
rect 41052 29291 41104 29300
rect 41052 29257 41061 29291
rect 41061 29257 41095 29291
rect 41095 29257 41104 29291
rect 41052 29248 41104 29257
rect 35532 29112 35584 29164
rect 31668 29044 31720 29096
rect 34704 29044 34756 29096
rect 37464 29044 37516 29096
rect 39672 29155 39724 29164
rect 16672 28951 16724 28960
rect 16672 28917 16681 28951
rect 16681 28917 16715 28951
rect 16715 28917 16724 28951
rect 16672 28908 16724 28917
rect 18328 28951 18380 28960
rect 18328 28917 18337 28951
rect 18337 28917 18371 28951
rect 18371 28917 18380 28951
rect 18328 28908 18380 28917
rect 36176 28976 36228 29028
rect 39672 29121 39681 29155
rect 39681 29121 39715 29155
rect 39715 29121 39724 29155
rect 39672 29112 39724 29121
rect 40684 29155 40736 29164
rect 40684 29121 40693 29155
rect 40693 29121 40727 29155
rect 40727 29121 40736 29155
rect 40684 29112 40736 29121
rect 45284 29248 45336 29300
rect 43352 29155 43404 29164
rect 43352 29121 43361 29155
rect 43361 29121 43395 29155
rect 43395 29121 43404 29155
rect 43352 29112 43404 29121
rect 38752 29087 38804 29096
rect 38752 29053 38761 29087
rect 38761 29053 38795 29087
rect 38795 29053 38804 29087
rect 38752 29044 38804 29053
rect 40316 29044 40368 29096
rect 42800 29044 42852 29096
rect 45008 29112 45060 29164
rect 45928 29044 45980 29096
rect 43628 28976 43680 29028
rect 19984 28908 20036 28960
rect 22008 28908 22060 28960
rect 24676 28908 24728 28960
rect 30196 28951 30248 28960
rect 30196 28917 30205 28951
rect 30205 28917 30239 28951
rect 30239 28917 30248 28951
rect 30196 28908 30248 28917
rect 43444 28908 43496 28960
rect 44272 28951 44324 28960
rect 44272 28917 44281 28951
rect 44281 28917 44315 28951
rect 44315 28917 44324 28951
rect 44272 28908 44324 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 65654 28806 65706 28858
rect 65718 28806 65770 28858
rect 65782 28806 65834 28858
rect 65846 28806 65898 28858
rect 65910 28806 65962 28858
rect 9128 28704 9180 28756
rect 9680 28568 9732 28620
rect 10324 28704 10376 28756
rect 12624 28704 12676 28756
rect 12808 28704 12860 28756
rect 14096 28747 14148 28756
rect 14096 28713 14105 28747
rect 14105 28713 14139 28747
rect 14139 28713 14148 28747
rect 14096 28704 14148 28713
rect 14556 28747 14608 28756
rect 14556 28713 14565 28747
rect 14565 28713 14599 28747
rect 14599 28713 14608 28747
rect 14556 28704 14608 28713
rect 19248 28747 19300 28756
rect 19248 28713 19257 28747
rect 19257 28713 19291 28747
rect 19291 28713 19300 28747
rect 19248 28704 19300 28713
rect 30840 28747 30892 28756
rect 30840 28713 30849 28747
rect 30849 28713 30883 28747
rect 30883 28713 30892 28747
rect 30840 28704 30892 28713
rect 11704 28636 11756 28688
rect 9588 28500 9640 28552
rect 11612 28543 11664 28552
rect 11612 28509 11621 28543
rect 11621 28509 11655 28543
rect 11655 28509 11664 28543
rect 11612 28500 11664 28509
rect 11152 28432 11204 28484
rect 12072 28543 12124 28552
rect 12072 28509 12086 28543
rect 12086 28509 12120 28543
rect 12120 28509 12124 28543
rect 16672 28636 16724 28688
rect 25412 28636 25464 28688
rect 12624 28568 12676 28620
rect 14188 28611 14240 28620
rect 14188 28577 14197 28611
rect 14197 28577 14231 28611
rect 14231 28577 14240 28611
rect 14188 28568 14240 28577
rect 14740 28568 14792 28620
rect 20260 28568 20312 28620
rect 21732 28611 21784 28620
rect 21732 28577 21741 28611
rect 21741 28577 21775 28611
rect 21775 28577 21784 28611
rect 21732 28568 21784 28577
rect 12072 28500 12124 28509
rect 11980 28475 12032 28484
rect 11980 28441 11989 28475
rect 11989 28441 12023 28475
rect 12023 28441 12032 28475
rect 11980 28432 12032 28441
rect 9312 28364 9364 28416
rect 13544 28500 13596 28552
rect 14004 28500 14056 28552
rect 14372 28543 14424 28552
rect 14372 28509 14381 28543
rect 14381 28509 14415 28543
rect 14415 28509 14424 28543
rect 14372 28500 14424 28509
rect 15200 28543 15252 28552
rect 15200 28509 15209 28543
rect 15209 28509 15243 28543
rect 15243 28509 15252 28543
rect 15200 28500 15252 28509
rect 16764 28543 16816 28552
rect 16764 28509 16773 28543
rect 16773 28509 16807 28543
rect 16807 28509 16816 28543
rect 16764 28500 16816 28509
rect 18328 28500 18380 28552
rect 19064 28500 19116 28552
rect 20076 28500 20128 28552
rect 22008 28543 22060 28552
rect 22008 28509 22042 28543
rect 22042 28509 22060 28543
rect 22008 28500 22060 28509
rect 24400 28543 24452 28552
rect 24400 28509 24409 28543
rect 24409 28509 24443 28543
rect 24443 28509 24452 28543
rect 24400 28500 24452 28509
rect 24676 28543 24728 28552
rect 24676 28509 24710 28543
rect 24710 28509 24728 28543
rect 24676 28500 24728 28509
rect 12440 28432 12492 28484
rect 17040 28475 17092 28484
rect 17040 28441 17049 28475
rect 17049 28441 17083 28475
rect 17083 28441 17092 28475
rect 17040 28432 17092 28441
rect 17132 28364 17184 28416
rect 17500 28364 17552 28416
rect 18328 28364 18380 28416
rect 19248 28364 19300 28416
rect 21088 28475 21140 28484
rect 21088 28441 21097 28475
rect 21097 28441 21131 28475
rect 21131 28441 21140 28475
rect 21088 28432 21140 28441
rect 21272 28432 21324 28484
rect 29644 28500 29696 28552
rect 28816 28432 28868 28484
rect 30932 28568 30984 28620
rect 31300 28568 31352 28620
rect 31484 28568 31536 28620
rect 36452 28704 36504 28756
rect 37188 28704 37240 28756
rect 40684 28636 40736 28688
rect 35992 28568 36044 28620
rect 37464 28568 37516 28620
rect 32588 28500 32640 28552
rect 36176 28500 36228 28552
rect 36360 28543 36412 28552
rect 36360 28509 36394 28543
rect 36394 28509 36412 28543
rect 36360 28500 36412 28509
rect 38108 28543 38160 28552
rect 38108 28509 38117 28543
rect 38117 28509 38151 28543
rect 38151 28509 38160 28543
rect 38108 28500 38160 28509
rect 42248 28543 42300 28552
rect 42248 28509 42257 28543
rect 42257 28509 42291 28543
rect 42291 28509 42300 28543
rect 42800 28543 42852 28552
rect 42248 28500 42300 28509
rect 42800 28509 42809 28543
rect 42809 28509 42843 28543
rect 42843 28509 42852 28543
rect 42800 28500 42852 28509
rect 43352 28568 43404 28620
rect 44272 28568 44324 28620
rect 43444 28543 43496 28552
rect 43444 28509 43453 28543
rect 43453 28509 43487 28543
rect 43487 28509 43496 28543
rect 43444 28500 43496 28509
rect 45284 28543 45336 28552
rect 36084 28432 36136 28484
rect 45284 28509 45293 28543
rect 45293 28509 45327 28543
rect 45327 28509 45336 28543
rect 45284 28500 45336 28509
rect 54576 28500 54628 28552
rect 67180 28500 67232 28552
rect 20904 28364 20956 28416
rect 22468 28364 22520 28416
rect 23112 28407 23164 28416
rect 23112 28373 23121 28407
rect 23121 28373 23155 28407
rect 23155 28373 23164 28407
rect 23112 28364 23164 28373
rect 25044 28364 25096 28416
rect 28264 28407 28316 28416
rect 28264 28373 28273 28407
rect 28273 28373 28307 28407
rect 28307 28373 28316 28407
rect 28264 28364 28316 28373
rect 31392 28364 31444 28416
rect 33416 28364 33468 28416
rect 34796 28364 34848 28416
rect 35624 28407 35676 28416
rect 35624 28373 35633 28407
rect 35633 28373 35667 28407
rect 35667 28373 35676 28407
rect 35624 28364 35676 28373
rect 37464 28407 37516 28416
rect 37464 28373 37473 28407
rect 37473 28373 37507 28407
rect 37507 28373 37516 28407
rect 37464 28364 37516 28373
rect 43996 28364 44048 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 7012 28160 7064 28212
rect 9956 28160 10008 28212
rect 10968 28160 11020 28212
rect 11796 28160 11848 28212
rect 11980 28160 12032 28212
rect 14372 28160 14424 28212
rect 15200 28160 15252 28212
rect 20168 28203 20220 28212
rect 14280 28092 14332 28144
rect 20168 28169 20177 28203
rect 20177 28169 20211 28203
rect 20211 28169 20220 28203
rect 20168 28160 20220 28169
rect 21272 28203 21324 28212
rect 21272 28169 21281 28203
rect 21281 28169 21315 28203
rect 21315 28169 21324 28203
rect 21272 28160 21324 28169
rect 22100 28203 22152 28212
rect 22100 28169 22109 28203
rect 22109 28169 22143 28203
rect 22143 28169 22152 28203
rect 22100 28160 22152 28169
rect 23112 28160 23164 28212
rect 23848 28160 23900 28212
rect 24584 28160 24636 28212
rect 24860 28160 24912 28212
rect 31300 28160 31352 28212
rect 31668 28160 31720 28212
rect 35348 28160 35400 28212
rect 35900 28160 35952 28212
rect 37372 28160 37424 28212
rect 37832 28203 37884 28212
rect 37832 28169 37841 28203
rect 37841 28169 37875 28203
rect 37875 28169 37884 28203
rect 37832 28160 37884 28169
rect 45468 28203 45520 28212
rect 45468 28169 45477 28203
rect 45477 28169 45511 28203
rect 45511 28169 45520 28203
rect 45468 28160 45520 28169
rect 45928 28203 45980 28212
rect 45928 28169 45937 28203
rect 45937 28169 45971 28203
rect 45971 28169 45980 28203
rect 45928 28160 45980 28169
rect 5908 28024 5960 28076
rect 6460 27999 6512 28008
rect 6460 27965 6469 27999
rect 6469 27965 6503 27999
rect 6503 27965 6512 27999
rect 6460 27956 6512 27965
rect 11060 28024 11112 28076
rect 12072 28024 12124 28076
rect 12164 28024 12216 28076
rect 12992 28024 13044 28076
rect 11244 27956 11296 28008
rect 11704 27888 11756 27940
rect 12164 27888 12216 27940
rect 15292 28024 15344 28076
rect 19248 28024 19300 28076
rect 20168 28024 20220 28076
rect 22468 28067 22520 28076
rect 22468 28033 22477 28067
rect 22477 28033 22511 28067
rect 22511 28033 22520 28067
rect 22468 28024 22520 28033
rect 23848 28024 23900 28076
rect 25044 28024 25096 28076
rect 28356 28067 28408 28076
rect 19432 27956 19484 28008
rect 22744 27999 22796 28008
rect 22744 27965 22753 27999
rect 22753 27965 22787 27999
rect 22787 27965 22796 27999
rect 22744 27956 22796 27965
rect 24216 27956 24268 28008
rect 15568 27888 15620 27940
rect 19984 27888 20036 27940
rect 28356 28033 28365 28067
rect 28365 28033 28399 28067
rect 28399 28033 28408 28067
rect 28356 28024 28408 28033
rect 30196 28024 30248 28076
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 43996 28135 44048 28144
rect 33416 28067 33468 28076
rect 33416 28033 33425 28067
rect 33425 28033 33459 28067
rect 33459 28033 33468 28067
rect 33416 28024 33468 28033
rect 35624 28024 35676 28076
rect 36084 28024 36136 28076
rect 27344 27956 27396 28008
rect 27528 27999 27580 28008
rect 27528 27965 27537 27999
rect 27537 27965 27571 27999
rect 27571 27965 27580 27999
rect 28264 27999 28316 28008
rect 27528 27956 27580 27965
rect 28264 27965 28273 27999
rect 28273 27965 28307 27999
rect 28307 27965 28316 27999
rect 28264 27956 28316 27965
rect 29644 27956 29696 28008
rect 30932 27999 30984 28008
rect 30932 27965 30941 27999
rect 30941 27965 30975 27999
rect 30975 27965 30984 27999
rect 30932 27956 30984 27965
rect 31024 27956 31076 28008
rect 8300 27820 8352 27872
rect 12808 27820 12860 27872
rect 13544 27820 13596 27872
rect 17132 27820 17184 27872
rect 17684 27820 17736 27872
rect 19064 27820 19116 27872
rect 26240 27820 26292 27872
rect 30288 27888 30340 27940
rect 31208 27888 31260 27940
rect 35532 27956 35584 28008
rect 37372 27956 37424 28008
rect 39304 27956 39356 28008
rect 37924 27888 37976 27940
rect 43996 28101 44005 28135
rect 44005 28101 44039 28135
rect 44039 28101 44048 28135
rect 43996 28092 44048 28101
rect 45836 28092 45888 28144
rect 43720 28067 43772 28076
rect 43720 28033 43729 28067
rect 43729 28033 43763 28067
rect 43763 28033 43772 28067
rect 43720 28024 43772 28033
rect 45468 28024 45520 28076
rect 45192 27956 45244 28008
rect 32404 27820 32456 27872
rect 33600 27863 33652 27872
rect 33600 27829 33609 27863
rect 33609 27829 33643 27863
rect 33643 27829 33652 27863
rect 33600 27820 33652 27829
rect 41420 27820 41472 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 65654 27718 65706 27770
rect 65718 27718 65770 27770
rect 65782 27718 65834 27770
rect 65846 27718 65898 27770
rect 65910 27718 65962 27770
rect 6460 27659 6512 27668
rect 6460 27625 6469 27659
rect 6469 27625 6503 27659
rect 6503 27625 6512 27659
rect 6460 27616 6512 27625
rect 11612 27616 11664 27668
rect 19248 27616 19300 27668
rect 22560 27616 22612 27668
rect 28356 27616 28408 27668
rect 31300 27616 31352 27668
rect 34612 27616 34664 27668
rect 34796 27616 34848 27668
rect 36084 27616 36136 27668
rect 37924 27659 37976 27668
rect 37924 27625 37933 27659
rect 37933 27625 37967 27659
rect 37967 27625 37976 27659
rect 37924 27616 37976 27625
rect 11152 27548 11204 27600
rect 19432 27548 19484 27600
rect 20352 27548 20404 27600
rect 9956 27523 10008 27532
rect 9956 27489 9965 27523
rect 9965 27489 9999 27523
rect 9999 27489 10008 27523
rect 9956 27480 10008 27489
rect 15108 27480 15160 27532
rect 4804 27412 4856 27464
rect 5080 27455 5132 27464
rect 5080 27421 5089 27455
rect 5089 27421 5123 27455
rect 5123 27421 5132 27455
rect 5080 27412 5132 27421
rect 7380 27412 7432 27464
rect 8760 27412 8812 27464
rect 6000 27344 6052 27396
rect 7748 27344 7800 27396
rect 11060 27412 11112 27464
rect 11704 27455 11756 27464
rect 9220 27387 9272 27396
rect 9220 27353 9229 27387
rect 9229 27353 9263 27387
rect 9263 27353 9272 27387
rect 9220 27344 9272 27353
rect 11704 27421 11713 27455
rect 11713 27421 11747 27455
rect 11747 27421 11756 27455
rect 11704 27412 11756 27421
rect 14740 27455 14792 27464
rect 14740 27421 14749 27455
rect 14749 27421 14783 27455
rect 14783 27421 14792 27455
rect 14740 27412 14792 27421
rect 15200 27412 15252 27464
rect 18236 27412 18288 27464
rect 20444 27480 20496 27532
rect 22008 27480 22060 27532
rect 20904 27412 20956 27464
rect 24400 27548 24452 27600
rect 23204 27480 23256 27532
rect 31024 27548 31076 27600
rect 32404 27548 32456 27600
rect 36452 27548 36504 27600
rect 40316 27591 40368 27600
rect 22652 27455 22704 27464
rect 22652 27421 22661 27455
rect 22661 27421 22695 27455
rect 22695 27421 22704 27455
rect 24768 27455 24820 27464
rect 22652 27412 22704 27421
rect 24768 27421 24797 27455
rect 24797 27421 24820 27455
rect 24768 27412 24820 27421
rect 29368 27480 29420 27532
rect 31208 27523 31260 27532
rect 31208 27489 31217 27523
rect 31217 27489 31251 27523
rect 31251 27489 31260 27523
rect 31208 27480 31260 27489
rect 39212 27480 39264 27532
rect 40316 27557 40325 27591
rect 40325 27557 40359 27591
rect 40359 27557 40368 27591
rect 40316 27548 40368 27557
rect 45008 27591 45060 27600
rect 45008 27557 45017 27591
rect 45017 27557 45051 27591
rect 45051 27557 45060 27591
rect 45008 27548 45060 27557
rect 45192 27591 45244 27600
rect 45192 27557 45201 27591
rect 45201 27557 45235 27591
rect 45235 27557 45244 27591
rect 45192 27548 45244 27557
rect 28816 27455 28868 27464
rect 28816 27421 28825 27455
rect 28825 27421 28859 27455
rect 28859 27421 28868 27455
rect 28816 27412 28868 27421
rect 31300 27455 31352 27464
rect 17040 27344 17092 27396
rect 17316 27344 17368 27396
rect 19340 27387 19392 27396
rect 19340 27353 19349 27387
rect 19349 27353 19383 27387
rect 19383 27353 19392 27387
rect 19340 27344 19392 27353
rect 19524 27344 19576 27396
rect 20168 27344 20220 27396
rect 20812 27344 20864 27396
rect 4712 27276 4764 27328
rect 6920 27319 6972 27328
rect 6920 27285 6929 27319
rect 6929 27285 6963 27319
rect 6963 27285 6972 27319
rect 6920 27276 6972 27285
rect 9312 27276 9364 27328
rect 10232 27319 10284 27328
rect 10232 27285 10241 27319
rect 10241 27285 10275 27319
rect 10275 27285 10284 27319
rect 10232 27276 10284 27285
rect 11244 27276 11296 27328
rect 12992 27276 13044 27328
rect 15568 27319 15620 27328
rect 15568 27285 15577 27319
rect 15577 27285 15611 27319
rect 15611 27285 15620 27319
rect 15568 27276 15620 27285
rect 18420 27276 18472 27328
rect 19984 27319 20036 27328
rect 19984 27285 19993 27319
rect 19993 27285 20027 27319
rect 20027 27285 20036 27319
rect 19984 27276 20036 27285
rect 23296 27276 23348 27328
rect 23664 27276 23716 27328
rect 25412 27276 25464 27328
rect 26240 27387 26292 27396
rect 26240 27353 26274 27387
rect 26274 27353 26292 27387
rect 26240 27344 26292 27353
rect 31300 27421 31309 27455
rect 31309 27421 31343 27455
rect 31343 27421 31352 27455
rect 31300 27412 31352 27421
rect 30288 27344 30340 27396
rect 37464 27412 37516 27464
rect 39304 27455 39356 27464
rect 39304 27421 39313 27455
rect 39313 27421 39347 27455
rect 39347 27421 39356 27455
rect 39304 27412 39356 27421
rect 41512 27480 41564 27532
rect 43444 27523 43496 27532
rect 43444 27489 43453 27523
rect 43453 27489 43487 27523
rect 43487 27489 43496 27523
rect 43444 27480 43496 27489
rect 45468 27523 45520 27532
rect 45468 27489 45477 27523
rect 45477 27489 45511 27523
rect 45511 27489 45520 27523
rect 45468 27480 45520 27489
rect 41420 27455 41472 27464
rect 39764 27344 39816 27396
rect 41420 27421 41429 27455
rect 41429 27421 41463 27455
rect 41463 27421 41472 27455
rect 41420 27412 41472 27421
rect 27344 27319 27396 27328
rect 27344 27285 27353 27319
rect 27353 27285 27387 27319
rect 27387 27285 27396 27319
rect 27344 27276 27396 27285
rect 29000 27319 29052 27328
rect 29000 27285 29009 27319
rect 29009 27285 29043 27319
rect 29043 27285 29052 27319
rect 29000 27276 29052 27285
rect 35532 27276 35584 27328
rect 36728 27319 36780 27328
rect 36728 27285 36737 27319
rect 36737 27285 36771 27319
rect 36771 27285 36780 27319
rect 36728 27276 36780 27285
rect 38660 27319 38712 27328
rect 38660 27285 38669 27319
rect 38669 27285 38703 27319
rect 38703 27285 38712 27319
rect 38660 27276 38712 27285
rect 39580 27276 39632 27328
rect 40224 27276 40276 27328
rect 41328 27319 41380 27328
rect 41328 27285 41337 27319
rect 41337 27285 41371 27319
rect 41371 27285 41380 27319
rect 41328 27276 41380 27285
rect 43628 27412 43680 27464
rect 42432 27319 42484 27328
rect 42432 27285 42441 27319
rect 42441 27285 42475 27319
rect 42475 27285 42484 27319
rect 42432 27276 42484 27285
rect 43904 27276 43956 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 7748 27115 7800 27124
rect 7748 27081 7757 27115
rect 7757 27081 7791 27115
rect 7791 27081 7800 27115
rect 7748 27072 7800 27081
rect 8760 27115 8812 27124
rect 8760 27081 8769 27115
rect 8769 27081 8803 27115
rect 8803 27081 8812 27115
rect 8760 27072 8812 27081
rect 4620 27004 4672 27056
rect 6920 27004 6972 27056
rect 4712 26979 4764 26988
rect 4712 26945 4746 26979
rect 4746 26945 4764 26979
rect 4712 26936 4764 26945
rect 5080 26936 5132 26988
rect 8300 26979 8352 26988
rect 8300 26945 8309 26979
rect 8309 26945 8343 26979
rect 8343 26945 8352 26979
rect 8300 26936 8352 26945
rect 6368 26911 6420 26920
rect 6368 26877 6377 26911
rect 6377 26877 6411 26911
rect 6411 26877 6420 26911
rect 6368 26868 6420 26877
rect 9680 27004 9732 27056
rect 10232 27004 10284 27056
rect 9588 26936 9640 26988
rect 10692 26911 10744 26920
rect 10692 26877 10701 26911
rect 10701 26877 10735 26911
rect 10735 26877 10744 26911
rect 10692 26868 10744 26877
rect 5172 26732 5224 26784
rect 6552 26732 6604 26784
rect 9128 26732 9180 26784
rect 9772 26775 9824 26784
rect 9772 26741 9781 26775
rect 9781 26741 9815 26775
rect 9815 26741 9824 26775
rect 9772 26732 9824 26741
rect 10232 26775 10284 26784
rect 10232 26741 10241 26775
rect 10241 26741 10275 26775
rect 10275 26741 10284 26775
rect 10232 26732 10284 26741
rect 12256 26868 12308 26920
rect 14096 27072 14148 27124
rect 17316 27115 17368 27124
rect 17316 27081 17325 27115
rect 17325 27081 17359 27115
rect 17359 27081 17368 27115
rect 17316 27072 17368 27081
rect 20352 27115 20404 27124
rect 20352 27081 20361 27115
rect 20361 27081 20395 27115
rect 20395 27081 20404 27115
rect 20352 27072 20404 27081
rect 23204 27115 23256 27124
rect 23204 27081 23213 27115
rect 23213 27081 23247 27115
rect 23247 27081 23256 27115
rect 23204 27072 23256 27081
rect 24216 27115 24268 27124
rect 24216 27081 24225 27115
rect 24225 27081 24259 27115
rect 24259 27081 24268 27115
rect 24216 27072 24268 27081
rect 25780 27072 25832 27124
rect 27528 27072 27580 27124
rect 12808 27004 12860 27056
rect 13176 26979 13228 26988
rect 13176 26945 13185 26979
rect 13185 26945 13219 26979
rect 13219 26945 13228 26979
rect 17040 27004 17092 27056
rect 13176 26936 13228 26945
rect 17132 26979 17184 26988
rect 17132 26945 17141 26979
rect 17141 26945 17175 26979
rect 17175 26945 17184 26979
rect 17132 26936 17184 26945
rect 18328 26979 18380 26988
rect 18328 26945 18362 26979
rect 18362 26945 18380 26979
rect 18328 26936 18380 26945
rect 12348 26800 12400 26852
rect 17868 26868 17920 26920
rect 12808 26800 12860 26852
rect 19984 27004 20036 27056
rect 29552 27004 29604 27056
rect 30932 27004 30984 27056
rect 40224 27072 40276 27124
rect 40500 27072 40552 27124
rect 45192 27072 45244 27124
rect 45836 27072 45888 27124
rect 38752 27004 38804 27056
rect 20628 26936 20680 26988
rect 23664 26936 23716 26988
rect 20720 26868 20772 26920
rect 23112 26868 23164 26920
rect 22744 26800 22796 26852
rect 25136 26936 25188 26988
rect 27436 26936 27488 26988
rect 32128 26979 32180 26988
rect 24952 26911 25004 26920
rect 24952 26877 24961 26911
rect 24961 26877 24995 26911
rect 24995 26877 25004 26911
rect 24952 26868 25004 26877
rect 32128 26945 32137 26979
rect 32137 26945 32171 26979
rect 32171 26945 32180 26979
rect 32128 26936 32180 26945
rect 34520 26979 34572 26988
rect 34520 26945 34529 26979
rect 34529 26945 34563 26979
rect 34563 26945 34572 26979
rect 34520 26936 34572 26945
rect 35624 26936 35676 26988
rect 38844 26979 38896 26988
rect 38844 26945 38853 26979
rect 38853 26945 38887 26979
rect 38887 26945 38896 26979
rect 38844 26936 38896 26945
rect 40776 27004 40828 27056
rect 43904 27047 43956 27056
rect 43904 27013 43913 27047
rect 43913 27013 43947 27047
rect 43947 27013 43956 27047
rect 43904 27004 43956 27013
rect 39580 26979 39632 26988
rect 39580 26945 39589 26979
rect 39589 26945 39623 26979
rect 39623 26945 39632 26979
rect 39580 26936 39632 26945
rect 34428 26868 34480 26920
rect 36084 26868 36136 26920
rect 38200 26868 38252 26920
rect 39764 26936 39816 26988
rect 39856 26868 39908 26920
rect 25872 26843 25924 26852
rect 25872 26809 25881 26843
rect 25881 26809 25915 26843
rect 25915 26809 25924 26843
rect 25872 26800 25924 26809
rect 36728 26800 36780 26852
rect 40040 26800 40092 26852
rect 41052 26979 41104 26988
rect 41052 26945 41061 26979
rect 41061 26945 41095 26979
rect 41095 26945 41104 26979
rect 41052 26936 41104 26945
rect 43628 26979 43680 26988
rect 43628 26945 43637 26979
rect 43637 26945 43671 26979
rect 43671 26945 43680 26979
rect 43628 26936 43680 26945
rect 45008 26936 45060 26988
rect 45284 26936 45336 26988
rect 13820 26732 13872 26784
rect 14004 26732 14056 26784
rect 14280 26775 14332 26784
rect 14280 26741 14289 26775
rect 14289 26741 14323 26775
rect 14323 26741 14332 26775
rect 14280 26732 14332 26741
rect 15568 26775 15620 26784
rect 15568 26741 15577 26775
rect 15577 26741 15611 26775
rect 15611 26741 15620 26775
rect 15568 26732 15620 26741
rect 19984 26732 20036 26784
rect 33232 26732 33284 26784
rect 34796 26732 34848 26784
rect 35624 26732 35676 26784
rect 39212 26732 39264 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 65654 26630 65706 26682
rect 65718 26630 65770 26682
rect 65782 26630 65834 26682
rect 65846 26630 65898 26682
rect 65910 26630 65962 26682
rect 4804 26571 4856 26580
rect 4804 26537 4813 26571
rect 4813 26537 4847 26571
rect 4847 26537 4856 26571
rect 4804 26528 4856 26537
rect 6000 26571 6052 26580
rect 6000 26537 6009 26571
rect 6009 26537 6043 26571
rect 6043 26537 6052 26571
rect 6000 26528 6052 26537
rect 7380 26571 7432 26580
rect 7380 26537 7389 26571
rect 7389 26537 7423 26571
rect 7423 26537 7432 26571
rect 7380 26528 7432 26537
rect 9220 26528 9272 26580
rect 9680 26528 9732 26580
rect 10692 26528 10744 26580
rect 11980 26528 12032 26580
rect 12256 26571 12308 26580
rect 12256 26537 12265 26571
rect 12265 26537 12299 26571
rect 12299 26537 12308 26571
rect 12256 26528 12308 26537
rect 12348 26528 12400 26580
rect 12992 26528 13044 26580
rect 5724 26460 5776 26512
rect 7288 26460 7340 26512
rect 9128 26503 9180 26512
rect 9128 26469 9137 26503
rect 9137 26469 9171 26503
rect 9171 26469 9180 26503
rect 9128 26460 9180 26469
rect 14280 26460 14332 26512
rect 15200 26528 15252 26580
rect 17960 26503 18012 26512
rect 17960 26469 17969 26503
rect 17969 26469 18003 26503
rect 18003 26469 18012 26503
rect 17960 26460 18012 26469
rect 20812 26503 20864 26512
rect 20812 26469 20821 26503
rect 20821 26469 20855 26503
rect 20855 26469 20864 26503
rect 20812 26460 20864 26469
rect 22652 26528 22704 26580
rect 27436 26528 27488 26580
rect 31852 26528 31904 26580
rect 36452 26528 36504 26580
rect 38200 26571 38252 26580
rect 38200 26537 38209 26571
rect 38209 26537 38243 26571
rect 38243 26537 38252 26571
rect 38200 26528 38252 26537
rect 39672 26528 39724 26580
rect 40776 26571 40828 26580
rect 40776 26537 40785 26571
rect 40785 26537 40819 26571
rect 40819 26537 40828 26571
rect 40776 26528 40828 26537
rect 45008 26528 45060 26580
rect 23572 26460 23624 26512
rect 29368 26460 29420 26512
rect 5448 26435 5500 26444
rect 5448 26401 5457 26435
rect 5457 26401 5491 26435
rect 5491 26401 5500 26435
rect 5448 26392 5500 26401
rect 7104 26392 7156 26444
rect 7564 26392 7616 26444
rect 9772 26392 9824 26444
rect 15384 26435 15436 26444
rect 5172 26367 5224 26376
rect 5172 26333 5181 26367
rect 5181 26333 5215 26367
rect 5215 26333 5224 26367
rect 5172 26324 5224 26333
rect 10232 26324 10284 26376
rect 11980 26324 12032 26376
rect 6920 26299 6972 26308
rect 6920 26265 6929 26299
rect 6929 26265 6963 26299
rect 6963 26265 6972 26299
rect 6920 26256 6972 26265
rect 7748 26256 7800 26308
rect 8300 26256 8352 26308
rect 10600 26299 10652 26308
rect 10600 26265 10609 26299
rect 10609 26265 10643 26299
rect 10643 26265 10652 26299
rect 10600 26256 10652 26265
rect 12072 26299 12124 26308
rect 12072 26265 12081 26299
rect 12081 26265 12115 26299
rect 12115 26265 12124 26299
rect 12072 26256 12124 26265
rect 12256 26324 12308 26376
rect 15384 26401 15393 26435
rect 15393 26401 15427 26435
rect 15427 26401 15436 26435
rect 15384 26392 15436 26401
rect 19156 26392 19208 26444
rect 20352 26392 20404 26444
rect 17960 26324 18012 26376
rect 18880 26324 18932 26376
rect 23204 26392 23256 26444
rect 24860 26392 24912 26444
rect 23296 26324 23348 26376
rect 25136 26392 25188 26444
rect 25228 26367 25280 26376
rect 25228 26333 25237 26367
rect 25237 26333 25271 26367
rect 25271 26333 25280 26367
rect 25228 26324 25280 26333
rect 29000 26367 29052 26376
rect 29000 26333 29009 26367
rect 29009 26333 29043 26367
rect 29043 26333 29052 26367
rect 29000 26324 29052 26333
rect 29552 26367 29604 26376
rect 29552 26333 29561 26367
rect 29561 26333 29595 26367
rect 29595 26333 29604 26367
rect 29552 26324 29604 26333
rect 31116 26392 31168 26444
rect 40408 26460 40460 26512
rect 40592 26460 40644 26512
rect 41328 26460 41380 26512
rect 68008 26503 68060 26512
rect 68008 26469 68017 26503
rect 68017 26469 68051 26503
rect 68051 26469 68060 26503
rect 68008 26460 68060 26469
rect 43628 26392 43680 26444
rect 32312 26367 32364 26376
rect 13084 26256 13136 26308
rect 13176 26256 13228 26308
rect 13636 26256 13688 26308
rect 13820 26256 13872 26308
rect 15660 26299 15712 26308
rect 15660 26265 15669 26299
rect 15669 26265 15703 26299
rect 15703 26265 15712 26299
rect 15660 26256 15712 26265
rect 15568 26188 15620 26240
rect 20076 26256 20128 26308
rect 30748 26256 30800 26308
rect 31944 26256 31996 26308
rect 32312 26333 32321 26367
rect 32321 26333 32355 26367
rect 32355 26333 32364 26367
rect 32312 26324 32364 26333
rect 34704 26367 34756 26376
rect 34704 26333 34713 26367
rect 34713 26333 34747 26367
rect 34747 26333 34756 26367
rect 34704 26324 34756 26333
rect 34796 26324 34848 26376
rect 37924 26367 37976 26376
rect 37924 26333 37933 26367
rect 37933 26333 37967 26367
rect 37967 26333 37976 26367
rect 37924 26324 37976 26333
rect 38844 26324 38896 26376
rect 39212 26324 39264 26376
rect 40040 26367 40092 26376
rect 40040 26333 40049 26367
rect 40049 26333 40083 26367
rect 40083 26333 40092 26367
rect 40040 26324 40092 26333
rect 40316 26367 40368 26376
rect 40316 26333 40325 26367
rect 40325 26333 40359 26367
rect 40359 26333 40368 26367
rect 40316 26324 40368 26333
rect 40684 26324 40736 26376
rect 41144 26367 41196 26376
rect 41144 26333 41153 26367
rect 41153 26333 41187 26367
rect 41187 26333 41196 26367
rect 41144 26324 41196 26333
rect 42432 26324 42484 26376
rect 45284 26324 45336 26376
rect 67824 26367 67876 26376
rect 67824 26333 67833 26367
rect 67833 26333 67867 26367
rect 67867 26333 67876 26367
rect 67824 26324 67876 26333
rect 32588 26256 32640 26308
rect 36452 26256 36504 26308
rect 38016 26299 38068 26308
rect 38016 26265 38025 26299
rect 38025 26265 38059 26299
rect 38059 26265 38068 26299
rect 38016 26256 38068 26265
rect 38200 26299 38252 26308
rect 38200 26265 38209 26299
rect 38209 26265 38243 26299
rect 38243 26265 38252 26299
rect 38200 26256 38252 26265
rect 24492 26188 24544 26240
rect 32680 26231 32732 26240
rect 32680 26197 32689 26231
rect 32689 26197 32723 26231
rect 32723 26197 32732 26231
rect 32680 26188 32732 26197
rect 36084 26231 36136 26240
rect 36084 26197 36093 26231
rect 36093 26197 36127 26231
rect 36127 26197 36136 26231
rect 36084 26188 36136 26197
rect 37464 26188 37516 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 5724 26027 5776 26036
rect 5724 25993 5733 26027
rect 5733 25993 5767 26027
rect 5767 25993 5776 26027
rect 5724 25984 5776 25993
rect 7932 25984 7984 26036
rect 10508 25984 10560 26036
rect 12440 25984 12492 26036
rect 6368 25916 6420 25968
rect 15384 25984 15436 26036
rect 15660 25984 15712 26036
rect 17132 25984 17184 26036
rect 19432 25984 19484 26036
rect 19800 25984 19852 26036
rect 4896 25891 4948 25900
rect 4896 25857 4905 25891
rect 4905 25857 4939 25891
rect 4939 25857 4948 25891
rect 4896 25848 4948 25857
rect 17040 25916 17092 25968
rect 18052 25916 18104 25968
rect 18236 25959 18288 25968
rect 18236 25925 18245 25959
rect 18245 25925 18279 25959
rect 18279 25925 18288 25959
rect 18236 25916 18288 25925
rect 20352 25916 20404 25968
rect 22744 25959 22796 25968
rect 22744 25925 22753 25959
rect 22753 25925 22787 25959
rect 22787 25925 22796 25959
rect 22744 25916 22796 25925
rect 32312 25984 32364 26036
rect 34520 25984 34572 26036
rect 38200 25984 38252 26036
rect 39856 25984 39908 26036
rect 41052 25984 41104 26036
rect 33232 25959 33284 25968
rect 33232 25925 33250 25959
rect 33250 25925 33284 25959
rect 33232 25916 33284 25925
rect 34612 25916 34664 25968
rect 9496 25891 9548 25900
rect 9496 25857 9530 25891
rect 9530 25857 9548 25891
rect 9496 25848 9548 25857
rect 10600 25848 10652 25900
rect 13176 25848 13228 25900
rect 14096 25848 14148 25900
rect 15568 25848 15620 25900
rect 16580 25848 16632 25900
rect 14280 25823 14332 25832
rect 14280 25789 14289 25823
rect 14289 25789 14323 25823
rect 14323 25789 14332 25823
rect 14280 25780 14332 25789
rect 14740 25823 14792 25832
rect 14740 25789 14749 25823
rect 14749 25789 14783 25823
rect 14783 25789 14792 25823
rect 14740 25780 14792 25789
rect 16488 25780 16540 25832
rect 19432 25848 19484 25900
rect 19800 25891 19852 25900
rect 19800 25857 19809 25891
rect 19809 25857 19843 25891
rect 19843 25857 19852 25891
rect 19800 25848 19852 25857
rect 20536 25848 20588 25900
rect 22008 25891 22060 25900
rect 22008 25857 22017 25891
rect 22017 25857 22051 25891
rect 22051 25857 22060 25891
rect 22008 25848 22060 25857
rect 23112 25848 23164 25900
rect 24216 25891 24268 25900
rect 13820 25712 13872 25764
rect 19340 25712 19392 25764
rect 4712 25687 4764 25696
rect 4712 25653 4721 25687
rect 4721 25653 4755 25687
rect 4755 25653 4764 25687
rect 4712 25644 4764 25653
rect 14924 25644 14976 25696
rect 22744 25780 22796 25832
rect 24216 25857 24225 25891
rect 24225 25857 24259 25891
rect 24259 25857 24268 25891
rect 24216 25848 24268 25857
rect 24492 25891 24544 25900
rect 24492 25857 24501 25891
rect 24501 25857 24535 25891
rect 24535 25857 24544 25891
rect 24492 25848 24544 25857
rect 24676 25891 24728 25900
rect 24676 25857 24690 25891
rect 24690 25857 24724 25891
rect 24724 25857 24728 25891
rect 25504 25891 25556 25900
rect 24676 25848 24728 25857
rect 25504 25857 25513 25891
rect 25513 25857 25547 25891
rect 25547 25857 25556 25891
rect 25504 25848 25556 25857
rect 32772 25848 32824 25900
rect 39304 25891 39356 25900
rect 39304 25857 39313 25891
rect 39313 25857 39347 25891
rect 39347 25857 39356 25891
rect 39304 25848 39356 25857
rect 40224 25891 40276 25900
rect 25412 25823 25464 25832
rect 25412 25789 25421 25823
rect 25421 25789 25455 25823
rect 25455 25789 25464 25823
rect 25412 25780 25464 25789
rect 32036 25780 32088 25832
rect 33508 25823 33560 25832
rect 33508 25789 33517 25823
rect 33517 25789 33551 25823
rect 33551 25789 33560 25823
rect 33508 25780 33560 25789
rect 25596 25712 25648 25764
rect 27528 25712 27580 25764
rect 35440 25780 35492 25832
rect 37464 25823 37516 25832
rect 37464 25789 37473 25823
rect 37473 25789 37507 25823
rect 37507 25789 37516 25823
rect 37464 25780 37516 25789
rect 40224 25857 40233 25891
rect 40233 25857 40267 25891
rect 40267 25857 40276 25891
rect 40224 25848 40276 25857
rect 40776 25848 40828 25900
rect 36084 25712 36136 25764
rect 37740 25755 37792 25764
rect 37740 25721 37749 25755
rect 37749 25721 37783 25755
rect 37783 25721 37792 25755
rect 37740 25712 37792 25721
rect 20444 25644 20496 25696
rect 24860 25687 24912 25696
rect 24860 25653 24869 25687
rect 24869 25653 24903 25687
rect 24903 25653 24912 25687
rect 24860 25644 24912 25653
rect 33232 25644 33284 25696
rect 36452 25687 36504 25696
rect 36452 25653 36461 25687
rect 36461 25653 36495 25687
rect 36495 25653 36504 25687
rect 36452 25644 36504 25653
rect 38752 25687 38804 25696
rect 38752 25653 38761 25687
rect 38761 25653 38795 25687
rect 38795 25653 38804 25687
rect 38752 25644 38804 25653
rect 41052 25644 41104 25696
rect 41512 25644 41564 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 65654 25542 65706 25594
rect 65718 25542 65770 25594
rect 65782 25542 65834 25594
rect 65846 25542 65898 25594
rect 65910 25542 65962 25594
rect 4896 25440 4948 25492
rect 9496 25440 9548 25492
rect 12900 25440 12952 25492
rect 14004 25440 14056 25492
rect 16856 25440 16908 25492
rect 18328 25440 18380 25492
rect 22744 25483 22796 25492
rect 22744 25449 22753 25483
rect 22753 25449 22787 25483
rect 22787 25449 22796 25483
rect 22744 25440 22796 25449
rect 24216 25440 24268 25492
rect 25504 25440 25556 25492
rect 27252 25440 27304 25492
rect 32128 25440 32180 25492
rect 32956 25483 33008 25492
rect 32956 25449 32965 25483
rect 32965 25449 32999 25483
rect 32999 25449 33008 25483
rect 32956 25440 33008 25449
rect 37740 25483 37792 25492
rect 37740 25449 37749 25483
rect 37749 25449 37783 25483
rect 37783 25449 37792 25483
rect 37740 25440 37792 25449
rect 37924 25483 37976 25492
rect 37924 25449 37933 25483
rect 37933 25449 37967 25483
rect 37967 25449 37976 25483
rect 37924 25440 37976 25449
rect 7564 25415 7616 25424
rect 7564 25381 7573 25415
rect 7573 25381 7607 25415
rect 7607 25381 7616 25415
rect 7564 25372 7616 25381
rect 13176 25372 13228 25424
rect 5540 25304 5592 25356
rect 16488 25304 16540 25356
rect 4620 25236 4672 25288
rect 4712 25168 4764 25220
rect 7932 25236 7984 25288
rect 9864 25279 9916 25288
rect 9864 25245 9873 25279
rect 9873 25245 9907 25279
rect 9907 25245 9916 25279
rect 9864 25236 9916 25245
rect 16856 25236 16908 25288
rect 19984 25304 20036 25356
rect 18696 25236 18748 25288
rect 20076 25236 20128 25288
rect 31484 25372 31536 25424
rect 22836 25304 22888 25356
rect 23020 25236 23072 25288
rect 23112 25236 23164 25288
rect 24860 25304 24912 25356
rect 24676 25279 24728 25288
rect 24676 25245 24685 25279
rect 24685 25245 24719 25279
rect 24719 25245 24728 25279
rect 24676 25236 24728 25245
rect 24952 25279 25004 25288
rect 24952 25245 24961 25279
rect 24961 25245 24995 25279
rect 24995 25245 25004 25279
rect 24952 25236 25004 25245
rect 25596 25279 25648 25288
rect 25596 25245 25605 25279
rect 25605 25245 25639 25279
rect 25639 25245 25648 25279
rect 25596 25236 25648 25245
rect 26700 25279 26752 25288
rect 26700 25245 26709 25279
rect 26709 25245 26743 25279
rect 26743 25245 26752 25279
rect 26700 25236 26752 25245
rect 30012 25304 30064 25356
rect 31852 25347 31904 25356
rect 31852 25313 31861 25347
rect 31861 25313 31895 25347
rect 31895 25313 31904 25347
rect 31852 25304 31904 25313
rect 32312 25304 32364 25356
rect 33140 25347 33192 25356
rect 33140 25313 33149 25347
rect 33149 25313 33183 25347
rect 33183 25313 33192 25347
rect 33140 25304 33192 25313
rect 29920 25236 29972 25288
rect 32680 25236 32732 25288
rect 33232 25279 33284 25288
rect 33232 25245 33241 25279
rect 33241 25245 33275 25279
rect 33275 25245 33284 25279
rect 33232 25236 33284 25245
rect 37464 25279 37516 25288
rect 14464 25211 14516 25220
rect 5632 25100 5684 25152
rect 14464 25177 14473 25211
rect 14473 25177 14507 25211
rect 14507 25177 14516 25211
rect 14464 25168 14516 25177
rect 20536 25168 20588 25220
rect 25136 25168 25188 25220
rect 34520 25168 34572 25220
rect 11612 25100 11664 25152
rect 11888 25100 11940 25152
rect 14096 25100 14148 25152
rect 15292 25143 15344 25152
rect 15292 25109 15301 25143
rect 15301 25109 15335 25143
rect 15335 25109 15344 25143
rect 15292 25100 15344 25109
rect 15384 25143 15436 25152
rect 15384 25109 15393 25143
rect 15393 25109 15427 25143
rect 15427 25109 15436 25143
rect 15384 25100 15436 25109
rect 15936 25100 15988 25152
rect 16856 25100 16908 25152
rect 19432 25100 19484 25152
rect 25688 25100 25740 25152
rect 27712 25100 27764 25152
rect 31208 25143 31260 25152
rect 31208 25109 31217 25143
rect 31217 25109 31251 25143
rect 31251 25109 31260 25143
rect 31208 25100 31260 25109
rect 33416 25143 33468 25152
rect 33416 25109 33425 25143
rect 33425 25109 33459 25143
rect 33459 25109 33468 25143
rect 33416 25100 33468 25109
rect 35900 25100 35952 25152
rect 37464 25245 37473 25279
rect 37473 25245 37507 25279
rect 37507 25245 37516 25279
rect 37464 25236 37516 25245
rect 60556 25279 60608 25288
rect 60556 25245 60565 25279
rect 60565 25245 60599 25279
rect 60599 25245 60608 25279
rect 60556 25236 60608 25245
rect 67824 25168 67876 25220
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 9864 24896 9916 24948
rect 10508 24939 10560 24948
rect 10508 24905 10517 24939
rect 10517 24905 10551 24939
rect 10551 24905 10560 24939
rect 10508 24896 10560 24905
rect 16488 24896 16540 24948
rect 20720 24896 20772 24948
rect 21456 24896 21508 24948
rect 29000 24896 29052 24948
rect 10692 24828 10744 24880
rect 5172 24760 5224 24812
rect 7380 24760 7432 24812
rect 7932 24760 7984 24812
rect 11888 24760 11940 24812
rect 12900 24828 12952 24880
rect 12808 24760 12860 24812
rect 6644 24735 6696 24744
rect 4712 24556 4764 24608
rect 6644 24701 6653 24735
rect 6653 24701 6687 24735
rect 6687 24701 6696 24735
rect 6644 24692 6696 24701
rect 11428 24692 11480 24744
rect 12900 24692 12952 24744
rect 13728 24828 13780 24880
rect 17040 24828 17092 24880
rect 19432 24828 19484 24880
rect 15936 24803 15988 24812
rect 13912 24735 13964 24744
rect 9772 24624 9824 24676
rect 9128 24556 9180 24608
rect 13084 24599 13136 24608
rect 13084 24565 13093 24599
rect 13093 24565 13127 24599
rect 13127 24565 13136 24599
rect 13084 24556 13136 24565
rect 13912 24701 13921 24735
rect 13921 24701 13955 24735
rect 13955 24701 13964 24735
rect 13912 24692 13964 24701
rect 15936 24769 15945 24803
rect 15945 24769 15979 24803
rect 15979 24769 15988 24803
rect 15936 24760 15988 24769
rect 17224 24803 17276 24812
rect 17224 24769 17233 24803
rect 17233 24769 17267 24803
rect 17267 24769 17276 24803
rect 17224 24760 17276 24769
rect 17592 24760 17644 24812
rect 20076 24760 20128 24812
rect 21916 24760 21968 24812
rect 24492 24760 24544 24812
rect 17868 24735 17920 24744
rect 17868 24701 17877 24735
rect 17877 24701 17911 24735
rect 17911 24701 17920 24735
rect 17868 24692 17920 24701
rect 18604 24692 18656 24744
rect 19156 24692 19208 24744
rect 22560 24692 22612 24744
rect 25688 24692 25740 24744
rect 29184 24828 29236 24880
rect 33416 24896 33468 24948
rect 45192 24896 45244 24948
rect 29092 24803 29144 24812
rect 29092 24769 29101 24803
rect 29101 24769 29135 24803
rect 29135 24769 29144 24803
rect 29092 24760 29144 24769
rect 29276 24803 29328 24812
rect 29276 24769 29285 24803
rect 29285 24769 29319 24803
rect 29319 24769 29328 24803
rect 29736 24803 29788 24812
rect 29276 24760 29328 24769
rect 29736 24769 29745 24803
rect 29745 24769 29779 24803
rect 29779 24769 29788 24803
rect 29736 24760 29788 24769
rect 32036 24760 32088 24812
rect 32312 24803 32364 24812
rect 32312 24769 32321 24803
rect 32321 24769 32355 24803
rect 32355 24769 32364 24803
rect 32312 24760 32364 24769
rect 28172 24735 28224 24744
rect 28172 24701 28181 24735
rect 28181 24701 28215 24735
rect 28215 24701 28224 24735
rect 28172 24692 28224 24701
rect 28724 24692 28776 24744
rect 27712 24624 27764 24676
rect 29920 24624 29972 24676
rect 31944 24692 31996 24744
rect 32588 24803 32640 24812
rect 32588 24769 32597 24803
rect 32597 24769 32631 24803
rect 32631 24769 32640 24803
rect 32588 24760 32640 24769
rect 34520 24760 34572 24812
rect 35716 24760 35768 24812
rect 34612 24692 34664 24744
rect 35440 24735 35492 24744
rect 35440 24701 35449 24735
rect 35449 24701 35483 24735
rect 35483 24701 35492 24735
rect 35440 24692 35492 24701
rect 39304 24760 39356 24812
rect 40592 24803 40644 24812
rect 40592 24769 40601 24803
rect 40601 24769 40635 24803
rect 40635 24769 40644 24803
rect 40592 24760 40644 24769
rect 45008 24760 45060 24812
rect 45284 24760 45336 24812
rect 14924 24556 14976 24608
rect 15292 24599 15344 24608
rect 15292 24565 15301 24599
rect 15301 24565 15335 24599
rect 15335 24565 15344 24599
rect 15292 24556 15344 24565
rect 16764 24556 16816 24608
rect 18512 24556 18564 24608
rect 20168 24556 20220 24608
rect 20444 24599 20496 24608
rect 20444 24565 20453 24599
rect 20453 24565 20487 24599
rect 20487 24565 20496 24599
rect 20444 24556 20496 24565
rect 21824 24556 21876 24608
rect 23296 24556 23348 24608
rect 24768 24556 24820 24608
rect 29000 24556 29052 24608
rect 29552 24556 29604 24608
rect 29736 24556 29788 24608
rect 38752 24624 38804 24676
rect 41144 24692 41196 24744
rect 45836 24692 45888 24744
rect 36360 24599 36412 24608
rect 36360 24565 36369 24599
rect 36369 24565 36403 24599
rect 36403 24565 36412 24599
rect 36360 24556 36412 24565
rect 40408 24556 40460 24608
rect 44180 24556 44232 24608
rect 45468 24599 45520 24608
rect 45468 24565 45477 24599
rect 45477 24565 45511 24599
rect 45511 24565 45520 24599
rect 45468 24556 45520 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 65654 24454 65706 24506
rect 65718 24454 65770 24506
rect 65782 24454 65834 24506
rect 65846 24454 65898 24506
rect 65910 24454 65962 24506
rect 9128 24352 9180 24404
rect 12808 24352 12860 24404
rect 16580 24395 16632 24404
rect 16580 24361 16589 24395
rect 16589 24361 16623 24395
rect 16623 24361 16632 24395
rect 16580 24352 16632 24361
rect 17960 24395 18012 24404
rect 17960 24361 17969 24395
rect 17969 24361 18003 24395
rect 18003 24361 18012 24395
rect 17960 24352 18012 24361
rect 15292 24284 15344 24336
rect 18144 24284 18196 24336
rect 18696 24284 18748 24336
rect 23572 24327 23624 24336
rect 23572 24293 23581 24327
rect 23581 24293 23615 24327
rect 23615 24293 23624 24327
rect 23572 24284 23624 24293
rect 24768 24284 24820 24336
rect 4712 24259 4764 24268
rect 4712 24225 4721 24259
rect 4721 24225 4755 24259
rect 4755 24225 4764 24259
rect 4712 24216 4764 24225
rect 7840 24216 7892 24268
rect 11704 24216 11756 24268
rect 14924 24259 14976 24268
rect 14924 24225 14933 24259
rect 14933 24225 14967 24259
rect 14967 24225 14976 24259
rect 14924 24216 14976 24225
rect 17868 24216 17920 24268
rect 22100 24216 22152 24268
rect 22560 24216 22612 24268
rect 25044 24216 25096 24268
rect 25780 24259 25832 24268
rect 25780 24225 25789 24259
rect 25789 24225 25823 24259
rect 25823 24225 25832 24259
rect 25780 24216 25832 24225
rect 29092 24352 29144 24404
rect 29184 24352 29236 24404
rect 30380 24284 30432 24336
rect 30840 24352 30892 24404
rect 34520 24284 34572 24336
rect 34612 24284 34664 24336
rect 35440 24352 35492 24404
rect 37648 24352 37700 24404
rect 40500 24352 40552 24404
rect 43628 24352 43680 24404
rect 45008 24395 45060 24404
rect 45008 24361 45017 24395
rect 45017 24361 45051 24395
rect 45051 24361 45060 24395
rect 45008 24352 45060 24361
rect 35808 24284 35860 24336
rect 28816 24216 28868 24268
rect 32036 24216 32088 24268
rect 34704 24216 34756 24268
rect 35992 24216 36044 24268
rect 6552 24191 6604 24200
rect 6552 24157 6561 24191
rect 6561 24157 6595 24191
rect 6595 24157 6604 24191
rect 6552 24148 6604 24157
rect 8024 24148 8076 24200
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 9128 24148 9180 24157
rect 11152 24191 11204 24200
rect 8116 24080 8168 24132
rect 8300 24080 8352 24132
rect 11152 24157 11161 24191
rect 11161 24157 11195 24191
rect 11195 24157 11204 24191
rect 11152 24148 11204 24157
rect 11520 24148 11572 24200
rect 13912 24148 13964 24200
rect 14648 24191 14700 24200
rect 14648 24157 14657 24191
rect 14657 24157 14691 24191
rect 14691 24157 14700 24191
rect 14648 24148 14700 24157
rect 5356 24012 5408 24064
rect 6736 24012 6788 24064
rect 7564 24012 7616 24064
rect 8852 24012 8904 24064
rect 9772 24012 9824 24064
rect 10692 24012 10744 24064
rect 11336 24055 11388 24064
rect 11336 24021 11345 24055
rect 11345 24021 11379 24055
rect 11379 24021 11388 24055
rect 11336 24012 11388 24021
rect 13360 24080 13412 24132
rect 15016 24080 15068 24132
rect 16120 24148 16172 24200
rect 16764 24191 16816 24200
rect 16764 24157 16773 24191
rect 16773 24157 16807 24191
rect 16807 24157 16816 24191
rect 16764 24148 16816 24157
rect 17500 24148 17552 24200
rect 18144 24148 18196 24200
rect 18512 24191 18564 24200
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 19432 24191 19484 24200
rect 16396 24080 16448 24132
rect 19432 24157 19441 24191
rect 19441 24157 19475 24191
rect 19475 24157 19484 24191
rect 19432 24148 19484 24157
rect 20444 24148 20496 24200
rect 19340 24080 19392 24132
rect 21088 24123 21140 24132
rect 21088 24089 21097 24123
rect 21097 24089 21131 24123
rect 21131 24089 21140 24123
rect 21088 24080 21140 24089
rect 21824 24080 21876 24132
rect 23388 24123 23440 24132
rect 23388 24089 23397 24123
rect 23397 24089 23431 24123
rect 23431 24089 23440 24123
rect 23388 24080 23440 24089
rect 24584 24080 24636 24132
rect 27344 24148 27396 24200
rect 28724 24191 28776 24200
rect 28724 24157 28753 24191
rect 28753 24157 28776 24191
rect 13820 24012 13872 24064
rect 15660 24055 15712 24064
rect 15660 24021 15669 24055
rect 15669 24021 15703 24055
rect 15703 24021 15712 24055
rect 15660 24012 15712 24021
rect 18512 24012 18564 24064
rect 27068 24012 27120 24064
rect 27252 24080 27304 24132
rect 28724 24148 28776 24157
rect 28172 24080 28224 24132
rect 30288 24191 30340 24200
rect 30288 24157 30297 24191
rect 30297 24157 30331 24191
rect 30331 24157 30340 24191
rect 30288 24148 30340 24157
rect 35900 24148 35952 24200
rect 39764 24216 39816 24268
rect 45284 24284 45336 24336
rect 45836 24284 45888 24336
rect 46848 24284 46900 24336
rect 45192 24259 45244 24268
rect 45192 24225 45201 24259
rect 45201 24225 45235 24259
rect 45235 24225 45244 24259
rect 45192 24216 45244 24225
rect 46020 24216 46072 24268
rect 38568 24148 38620 24200
rect 40500 24191 40552 24200
rect 40500 24157 40509 24191
rect 40509 24157 40543 24191
rect 40543 24157 40552 24191
rect 40500 24148 40552 24157
rect 44272 24191 44324 24200
rect 36360 24123 36412 24132
rect 36360 24089 36394 24123
rect 36394 24089 36412 24123
rect 30104 24012 30156 24064
rect 32864 24012 32916 24064
rect 36360 24080 36412 24089
rect 40776 24123 40828 24132
rect 40776 24089 40785 24123
rect 40785 24089 40819 24123
rect 40819 24089 40828 24123
rect 40776 24080 40828 24089
rect 42524 24080 42576 24132
rect 34520 24012 34572 24064
rect 38108 24012 38160 24064
rect 42248 24055 42300 24064
rect 42248 24021 42257 24055
rect 42257 24021 42291 24055
rect 42291 24021 42300 24055
rect 42248 24012 42300 24021
rect 42340 24012 42392 24064
rect 44272 24157 44281 24191
rect 44281 24157 44315 24191
rect 44315 24157 44324 24191
rect 44272 24148 44324 24157
rect 45284 24191 45336 24200
rect 45284 24157 45293 24191
rect 45293 24157 45327 24191
rect 45327 24157 45336 24191
rect 45284 24148 45336 24157
rect 44088 24080 44140 24132
rect 44732 24080 44784 24132
rect 44640 24012 44692 24064
rect 45652 24055 45704 24064
rect 45652 24021 45661 24055
rect 45661 24021 45695 24055
rect 45695 24021 45704 24055
rect 45652 24012 45704 24021
rect 46940 24012 46992 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 7380 23851 7432 23860
rect 7380 23817 7389 23851
rect 7389 23817 7423 23851
rect 7423 23817 7432 23851
rect 7380 23808 7432 23817
rect 8116 23851 8168 23860
rect 8116 23817 8125 23851
rect 8125 23817 8159 23851
rect 8159 23817 8168 23851
rect 8116 23808 8168 23817
rect 10876 23808 10928 23860
rect 12900 23851 12952 23860
rect 12900 23817 12909 23851
rect 12909 23817 12943 23851
rect 12943 23817 12952 23851
rect 12900 23808 12952 23817
rect 13360 23851 13412 23860
rect 13360 23817 13369 23851
rect 13369 23817 13403 23851
rect 13403 23817 13412 23851
rect 13360 23808 13412 23817
rect 14096 23851 14148 23860
rect 14096 23817 14105 23851
rect 14105 23817 14139 23851
rect 14139 23817 14148 23851
rect 14096 23808 14148 23817
rect 19432 23808 19484 23860
rect 21088 23808 21140 23860
rect 22836 23851 22888 23860
rect 22836 23817 22845 23851
rect 22845 23817 22879 23851
rect 22879 23817 22888 23851
rect 22836 23808 22888 23817
rect 23020 23808 23072 23860
rect 23756 23808 23808 23860
rect 24584 23851 24636 23860
rect 24584 23817 24593 23851
rect 24593 23817 24627 23851
rect 24627 23817 24636 23851
rect 24584 23808 24636 23817
rect 25688 23851 25740 23860
rect 25688 23817 25697 23851
rect 25697 23817 25731 23851
rect 25731 23817 25740 23851
rect 25688 23808 25740 23817
rect 26608 23808 26660 23860
rect 5632 23783 5684 23792
rect 5632 23749 5641 23783
rect 5641 23749 5675 23783
rect 5675 23749 5684 23783
rect 5632 23740 5684 23749
rect 6736 23715 6788 23724
rect 6736 23681 6745 23715
rect 6745 23681 6779 23715
rect 6779 23681 6788 23715
rect 6736 23672 6788 23681
rect 7564 23715 7616 23724
rect 7564 23681 7573 23715
rect 7573 23681 7607 23715
rect 7607 23681 7616 23715
rect 7564 23672 7616 23681
rect 8024 23715 8076 23724
rect 8024 23681 8033 23715
rect 8033 23681 8067 23715
rect 8067 23681 8076 23715
rect 8024 23672 8076 23681
rect 8300 23672 8352 23724
rect 10140 23740 10192 23792
rect 8852 23715 8904 23724
rect 8852 23681 8861 23715
rect 8861 23681 8895 23715
rect 8895 23681 8904 23715
rect 8852 23672 8904 23681
rect 9772 23715 9824 23724
rect 9772 23681 9781 23715
rect 9781 23681 9815 23715
rect 9815 23681 9824 23715
rect 9772 23672 9824 23681
rect 10692 23715 10744 23724
rect 6552 23604 6604 23656
rect 5724 23536 5776 23588
rect 10692 23681 10701 23715
rect 10701 23681 10735 23715
rect 10735 23681 10744 23715
rect 10692 23672 10744 23681
rect 11336 23740 11388 23792
rect 11888 23740 11940 23792
rect 17132 23740 17184 23792
rect 17500 23783 17552 23792
rect 17500 23749 17509 23783
rect 17509 23749 17543 23783
rect 17543 23749 17552 23783
rect 17500 23740 17552 23749
rect 18604 23783 18656 23792
rect 18604 23749 18613 23783
rect 18613 23749 18647 23783
rect 18647 23749 18656 23783
rect 18604 23740 18656 23749
rect 23388 23740 23440 23792
rect 12532 23672 12584 23724
rect 14004 23672 14056 23724
rect 15200 23672 15252 23724
rect 15844 23672 15896 23724
rect 17224 23672 17276 23724
rect 17592 23715 17644 23724
rect 17592 23681 17601 23715
rect 17601 23681 17635 23715
rect 17635 23681 17644 23715
rect 17592 23672 17644 23681
rect 18512 23715 18564 23724
rect 18512 23681 18521 23715
rect 18521 23681 18555 23715
rect 18555 23681 18564 23715
rect 18512 23672 18564 23681
rect 11520 23647 11572 23656
rect 10140 23536 10192 23588
rect 11520 23613 11529 23647
rect 11529 23613 11563 23647
rect 11563 23613 11572 23647
rect 11520 23604 11572 23613
rect 5816 23511 5868 23520
rect 5816 23477 5825 23511
rect 5825 23477 5859 23511
rect 5859 23477 5868 23511
rect 5816 23468 5868 23477
rect 9128 23468 9180 23520
rect 10416 23511 10468 23520
rect 10416 23477 10425 23511
rect 10425 23477 10459 23511
rect 10459 23477 10468 23511
rect 10416 23468 10468 23477
rect 16764 23604 16816 23656
rect 18052 23604 18104 23656
rect 19984 23672 20036 23724
rect 20536 23715 20588 23724
rect 20536 23681 20545 23715
rect 20545 23681 20579 23715
rect 20579 23681 20588 23715
rect 20536 23672 20588 23681
rect 27252 23740 27304 23792
rect 27528 23740 27580 23792
rect 25780 23672 25832 23724
rect 27160 23715 27212 23724
rect 27160 23681 27169 23715
rect 27169 23681 27203 23715
rect 27203 23681 27212 23715
rect 27160 23672 27212 23681
rect 19248 23604 19300 23656
rect 16120 23579 16172 23588
rect 16120 23545 16129 23579
rect 16129 23545 16163 23579
rect 16163 23545 16172 23579
rect 16120 23536 16172 23545
rect 16396 23536 16448 23588
rect 19156 23536 19208 23588
rect 23388 23604 23440 23656
rect 26056 23647 26108 23656
rect 26056 23613 26065 23647
rect 26065 23613 26099 23647
rect 26099 23613 26108 23647
rect 26056 23604 26108 23613
rect 27068 23647 27120 23656
rect 27068 23613 27077 23647
rect 27077 23613 27111 23647
rect 27111 23613 27120 23647
rect 27068 23604 27120 23613
rect 20536 23536 20588 23588
rect 32956 23808 33008 23860
rect 29092 23672 29144 23724
rect 29276 23672 29328 23724
rect 29920 23715 29972 23724
rect 29920 23681 29929 23715
rect 29929 23681 29963 23715
rect 29963 23681 29972 23715
rect 29920 23672 29972 23681
rect 30288 23672 30340 23724
rect 28816 23604 28868 23656
rect 30380 23604 30432 23656
rect 31944 23740 31996 23792
rect 30748 23715 30800 23724
rect 30748 23681 30757 23715
rect 30757 23681 30791 23715
rect 30791 23681 30800 23715
rect 30748 23672 30800 23681
rect 30840 23715 30892 23724
rect 30840 23681 30849 23715
rect 30849 23681 30883 23715
rect 30883 23681 30892 23715
rect 32220 23715 32272 23724
rect 30840 23672 30892 23681
rect 32220 23681 32229 23715
rect 32229 23681 32263 23715
rect 32263 23681 32272 23715
rect 32220 23672 32272 23681
rect 33048 23715 33100 23724
rect 31944 23604 31996 23656
rect 32312 23604 32364 23656
rect 33048 23681 33057 23715
rect 33057 23681 33091 23715
rect 33091 23681 33100 23715
rect 33048 23672 33100 23681
rect 29828 23536 29880 23588
rect 31576 23536 31628 23588
rect 33600 23740 33652 23792
rect 33324 23672 33376 23724
rect 35348 23851 35400 23860
rect 35348 23817 35357 23851
rect 35357 23817 35391 23851
rect 35391 23817 35400 23851
rect 35348 23808 35400 23817
rect 40776 23851 40828 23860
rect 40776 23817 40785 23851
rect 40785 23817 40819 23851
rect 40819 23817 40828 23851
rect 40776 23808 40828 23817
rect 40868 23808 40920 23860
rect 42340 23808 42392 23860
rect 42524 23851 42576 23860
rect 42524 23817 42533 23851
rect 42533 23817 42567 23851
rect 42567 23817 42576 23851
rect 42524 23808 42576 23817
rect 44180 23783 44232 23792
rect 35348 23672 35400 23724
rect 35808 23672 35860 23724
rect 37648 23715 37700 23724
rect 37648 23681 37657 23715
rect 37657 23681 37691 23715
rect 37691 23681 37700 23715
rect 37648 23672 37700 23681
rect 16488 23468 16540 23520
rect 23664 23468 23716 23520
rect 28264 23511 28316 23520
rect 28264 23477 28273 23511
rect 28273 23477 28307 23511
rect 28307 23477 28316 23511
rect 28264 23468 28316 23477
rect 29920 23468 29972 23520
rect 30748 23468 30800 23520
rect 33232 23468 33284 23520
rect 33692 23511 33744 23520
rect 33692 23477 33701 23511
rect 33701 23477 33735 23511
rect 33735 23477 33744 23511
rect 33692 23468 33744 23477
rect 38660 23647 38712 23656
rect 38660 23613 38669 23647
rect 38669 23613 38703 23647
rect 38703 23613 38712 23647
rect 38660 23604 38712 23613
rect 44180 23749 44189 23783
rect 44189 23749 44223 23783
rect 44223 23749 44232 23783
rect 44180 23740 44232 23749
rect 44640 23740 44692 23792
rect 47584 23740 47636 23792
rect 41236 23715 41288 23724
rect 41236 23681 41245 23715
rect 41245 23681 41279 23715
rect 41279 23681 41288 23715
rect 41236 23672 41288 23681
rect 43260 23715 43312 23724
rect 39764 23647 39816 23656
rect 39764 23613 39773 23647
rect 39773 23613 39807 23647
rect 39807 23613 39816 23647
rect 39764 23604 39816 23613
rect 43260 23681 43269 23715
rect 43269 23681 43303 23715
rect 43303 23681 43312 23715
rect 43260 23672 43312 23681
rect 43628 23672 43680 23724
rect 48688 23715 48740 23724
rect 48688 23681 48697 23715
rect 48697 23681 48731 23715
rect 48731 23681 48740 23715
rect 48688 23672 48740 23681
rect 57704 23672 57756 23724
rect 42800 23604 42852 23656
rect 44272 23604 44324 23656
rect 46020 23604 46072 23656
rect 46848 23604 46900 23656
rect 46940 23536 46992 23588
rect 44548 23468 44600 23520
rect 47400 23468 47452 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 65654 23366 65706 23418
rect 65718 23366 65770 23418
rect 65782 23366 65834 23418
rect 65846 23366 65898 23418
rect 65910 23366 65962 23418
rect 8300 23307 8352 23316
rect 8300 23273 8309 23307
rect 8309 23273 8343 23307
rect 8343 23273 8352 23307
rect 8300 23264 8352 23273
rect 11152 23307 11204 23316
rect 11152 23273 11161 23307
rect 11161 23273 11195 23307
rect 11195 23273 11204 23307
rect 11152 23264 11204 23273
rect 14004 23264 14056 23316
rect 16764 23307 16816 23316
rect 16764 23273 16773 23307
rect 16773 23273 16807 23307
rect 16807 23273 16816 23307
rect 19248 23307 19300 23316
rect 16764 23264 16816 23273
rect 11428 23196 11480 23248
rect 11520 23196 11572 23248
rect 11704 23171 11756 23180
rect 11704 23137 11713 23171
rect 11713 23137 11747 23171
rect 11747 23137 11756 23171
rect 11704 23128 11756 23137
rect 17684 23196 17736 23248
rect 19248 23273 19257 23307
rect 19257 23273 19291 23307
rect 19291 23273 19300 23307
rect 19248 23264 19300 23273
rect 20260 23264 20312 23316
rect 28172 23264 28224 23316
rect 29276 23264 29328 23316
rect 35440 23264 35492 23316
rect 37832 23264 37884 23316
rect 38108 23264 38160 23316
rect 23388 23196 23440 23248
rect 30840 23196 30892 23248
rect 33324 23239 33376 23248
rect 33324 23205 33333 23239
rect 33333 23205 33367 23239
rect 33367 23205 33376 23239
rect 33324 23196 33376 23205
rect 38660 23264 38712 23316
rect 41236 23307 41288 23316
rect 41236 23273 41245 23307
rect 41245 23273 41279 23307
rect 41279 23273 41288 23307
rect 41236 23264 41288 23273
rect 43260 23264 43312 23316
rect 5356 23103 5408 23112
rect 5356 23069 5365 23103
rect 5365 23069 5399 23103
rect 5399 23069 5408 23103
rect 5356 23060 5408 23069
rect 5540 23103 5592 23112
rect 5540 23069 5547 23103
rect 5547 23069 5592 23103
rect 5540 23060 5592 23069
rect 5724 23103 5776 23112
rect 5724 23069 5733 23103
rect 5733 23069 5767 23103
rect 5767 23069 5776 23103
rect 5724 23060 5776 23069
rect 5816 23103 5868 23112
rect 5816 23069 5830 23103
rect 5830 23069 5864 23103
rect 5864 23069 5868 23103
rect 5816 23060 5868 23069
rect 14096 23128 14148 23180
rect 14464 23128 14516 23180
rect 19524 23128 19576 23180
rect 20168 23128 20220 23180
rect 22100 23128 22152 23180
rect 30380 23128 30432 23180
rect 31576 23128 31628 23180
rect 13912 23060 13964 23112
rect 15660 23103 15712 23112
rect 15660 23069 15694 23103
rect 15694 23069 15712 23103
rect 15660 23060 15712 23069
rect 17776 23060 17828 23112
rect 18328 23060 18380 23112
rect 19340 23060 19392 23112
rect 6368 22992 6420 23044
rect 12900 22992 12952 23044
rect 13820 22992 13872 23044
rect 12440 22924 12492 22976
rect 13728 22924 13780 22976
rect 14556 22967 14608 22976
rect 14556 22933 14565 22967
rect 14565 22933 14599 22967
rect 14599 22933 14608 22967
rect 14556 22924 14608 22933
rect 20812 23060 20864 23112
rect 22836 23060 22888 23112
rect 26424 23103 26476 23112
rect 26424 23069 26433 23103
rect 26433 23069 26467 23103
rect 26467 23069 26476 23103
rect 26424 23060 26476 23069
rect 26608 23103 26660 23112
rect 26608 23069 26617 23103
rect 26617 23069 26651 23103
rect 26651 23069 26660 23103
rect 26608 23060 26660 23069
rect 27712 23103 27764 23112
rect 27712 23069 27721 23103
rect 27721 23069 27755 23103
rect 27755 23069 27764 23103
rect 27712 23060 27764 23069
rect 28356 23060 28408 23112
rect 29552 23103 29604 23112
rect 29552 23069 29561 23103
rect 29561 23069 29595 23103
rect 29595 23069 29604 23103
rect 29552 23060 29604 23069
rect 29736 23103 29788 23112
rect 29736 23069 29743 23103
rect 29743 23069 29788 23103
rect 29736 23060 29788 23069
rect 29920 23103 29972 23112
rect 29920 23069 29929 23103
rect 29929 23069 29963 23103
rect 29963 23069 29972 23103
rect 29920 23060 29972 23069
rect 30104 23060 30156 23112
rect 31484 23103 31536 23112
rect 31484 23069 31493 23103
rect 31493 23069 31527 23103
rect 31527 23069 31536 23103
rect 31484 23060 31536 23069
rect 32772 23060 32824 23112
rect 37832 23128 37884 23180
rect 38568 23128 38620 23180
rect 39028 23128 39080 23180
rect 40868 23128 40920 23180
rect 42248 23196 42300 23248
rect 42800 23239 42852 23248
rect 42800 23205 42809 23239
rect 42809 23205 42843 23239
rect 42843 23205 42852 23239
rect 42800 23196 42852 23205
rect 43720 23196 43772 23248
rect 45652 23264 45704 23316
rect 46020 23196 46072 23248
rect 45284 23128 45336 23180
rect 46940 23171 46992 23180
rect 46940 23137 46949 23171
rect 46949 23137 46983 23171
rect 46983 23137 46992 23171
rect 46940 23128 46992 23137
rect 34520 23060 34572 23112
rect 35532 23060 35584 23112
rect 41880 23103 41932 23112
rect 20536 22992 20588 23044
rect 20904 22992 20956 23044
rect 20628 22967 20680 22976
rect 20628 22933 20637 22967
rect 20637 22933 20671 22967
rect 20671 22933 20680 22967
rect 20628 22924 20680 22933
rect 21916 22924 21968 22976
rect 23480 22992 23532 23044
rect 26240 22992 26292 23044
rect 29828 23035 29880 23044
rect 24676 22924 24728 22976
rect 27344 22924 27396 22976
rect 27804 22967 27856 22976
rect 27804 22933 27813 22967
rect 27813 22933 27847 22967
rect 27847 22933 27856 22967
rect 27804 22924 27856 22933
rect 29828 23001 29837 23035
rect 29837 23001 29871 23035
rect 29871 23001 29880 23035
rect 29828 22992 29880 23001
rect 31208 22992 31260 23044
rect 40776 23035 40828 23044
rect 30196 22967 30248 22976
rect 30196 22933 30205 22967
rect 30205 22933 30239 22967
rect 30239 22933 30248 22967
rect 30196 22924 30248 22933
rect 32404 22924 32456 22976
rect 35532 22924 35584 22976
rect 35716 22924 35768 22976
rect 37556 22924 37608 22976
rect 40776 23001 40785 23035
rect 40785 23001 40819 23035
rect 40819 23001 40828 23035
rect 41880 23069 41889 23103
rect 41889 23069 41923 23103
rect 41923 23069 41932 23103
rect 41880 23060 41932 23069
rect 44548 23060 44600 23112
rect 45836 23060 45888 23112
rect 47400 23103 47452 23112
rect 47400 23069 47409 23103
rect 47409 23069 47443 23103
rect 47443 23069 47452 23103
rect 47400 23060 47452 23069
rect 42616 23035 42668 23044
rect 40776 22992 40828 23001
rect 42616 23001 42625 23035
rect 42625 23001 42659 23035
rect 42659 23001 42668 23035
rect 42616 22992 42668 23001
rect 39856 22967 39908 22976
rect 39856 22933 39865 22967
rect 39865 22933 39899 22967
rect 39899 22933 39908 22967
rect 39856 22924 39908 22933
rect 39948 22924 40000 22976
rect 44180 22924 44232 22976
rect 46112 22924 46164 22976
rect 47584 22967 47636 22976
rect 47584 22933 47593 22967
rect 47593 22933 47627 22967
rect 47627 22933 47636 22967
rect 47584 22924 47636 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 5540 22763 5592 22772
rect 5540 22729 5549 22763
rect 5549 22729 5583 22763
rect 5583 22729 5592 22763
rect 5540 22720 5592 22729
rect 6368 22763 6420 22772
rect 6368 22729 6377 22763
rect 6377 22729 6411 22763
rect 6411 22729 6420 22763
rect 6368 22720 6420 22729
rect 11060 22720 11112 22772
rect 12532 22720 12584 22772
rect 5356 22627 5408 22636
rect 5356 22593 5365 22627
rect 5365 22593 5399 22627
rect 5399 22593 5408 22627
rect 5356 22584 5408 22593
rect 12440 22584 12492 22636
rect 14648 22720 14700 22772
rect 16764 22720 16816 22772
rect 17132 22763 17184 22772
rect 17132 22729 17141 22763
rect 17141 22729 17175 22763
rect 17175 22729 17184 22763
rect 17132 22720 17184 22729
rect 17224 22720 17276 22772
rect 18420 22720 18472 22772
rect 19524 22763 19576 22772
rect 19524 22729 19533 22763
rect 19533 22729 19567 22763
rect 19567 22729 19576 22763
rect 19524 22720 19576 22729
rect 23388 22720 23440 22772
rect 25872 22720 25924 22772
rect 26792 22720 26844 22772
rect 27344 22763 27396 22772
rect 13084 22695 13136 22704
rect 13084 22661 13093 22695
rect 13093 22661 13127 22695
rect 13127 22661 13136 22695
rect 13084 22652 13136 22661
rect 14556 22652 14608 22704
rect 18604 22652 18656 22704
rect 20260 22652 20312 22704
rect 12900 22584 12952 22636
rect 14188 22584 14240 22636
rect 17960 22627 18012 22636
rect 17960 22593 17969 22627
rect 17969 22593 18003 22627
rect 18003 22593 18012 22627
rect 17960 22584 18012 22593
rect 18696 22584 18748 22636
rect 20168 22584 20220 22636
rect 20536 22627 20588 22636
rect 20536 22593 20545 22627
rect 20545 22593 20579 22627
rect 20579 22593 20588 22627
rect 20536 22584 20588 22593
rect 20812 22627 20864 22636
rect 20812 22593 20821 22627
rect 20821 22593 20855 22627
rect 20855 22593 20864 22627
rect 20812 22584 20864 22593
rect 21548 22584 21600 22636
rect 5908 22448 5960 22500
rect 7932 22380 7984 22432
rect 18052 22516 18104 22568
rect 22100 22516 22152 22568
rect 22284 22516 22336 22568
rect 27344 22729 27353 22763
rect 27353 22729 27387 22763
rect 27387 22729 27396 22763
rect 27344 22720 27396 22729
rect 27436 22763 27488 22772
rect 27436 22729 27445 22763
rect 27445 22729 27479 22763
rect 27479 22729 27488 22763
rect 27436 22720 27488 22729
rect 26792 22516 26844 22568
rect 14004 22491 14056 22500
rect 14004 22457 14013 22491
rect 14013 22457 14047 22491
rect 14047 22457 14056 22491
rect 14004 22448 14056 22457
rect 17776 22448 17828 22500
rect 18880 22448 18932 22500
rect 23480 22448 23532 22500
rect 25136 22491 25188 22500
rect 25136 22457 25145 22491
rect 25145 22457 25179 22491
rect 25179 22457 25188 22491
rect 25136 22448 25188 22457
rect 30288 22720 30340 22772
rect 31944 22720 31996 22772
rect 32220 22720 32272 22772
rect 35440 22763 35492 22772
rect 27804 22652 27856 22704
rect 35440 22729 35449 22763
rect 35449 22729 35483 22763
rect 35483 22729 35492 22763
rect 35440 22720 35492 22729
rect 40776 22652 40828 22704
rect 46020 22720 46072 22772
rect 43720 22652 43772 22704
rect 44180 22695 44232 22704
rect 44180 22661 44189 22695
rect 44189 22661 44223 22695
rect 44223 22661 44232 22695
rect 44180 22652 44232 22661
rect 45468 22652 45520 22704
rect 29920 22627 29972 22636
rect 29920 22593 29929 22627
rect 29929 22593 29963 22627
rect 29963 22593 29972 22627
rect 29920 22584 29972 22593
rect 30104 22584 30156 22636
rect 31760 22584 31812 22636
rect 33416 22627 33468 22636
rect 33416 22593 33425 22627
rect 33425 22593 33459 22627
rect 33459 22593 33468 22627
rect 33416 22584 33468 22593
rect 30288 22516 30340 22568
rect 33232 22559 33284 22568
rect 31484 22491 31536 22500
rect 31484 22457 31493 22491
rect 31493 22457 31527 22491
rect 31527 22457 31536 22491
rect 31484 22448 31536 22457
rect 33232 22525 33241 22559
rect 33241 22525 33275 22559
rect 33275 22525 33284 22559
rect 33232 22516 33284 22525
rect 18512 22423 18564 22432
rect 18512 22389 18521 22423
rect 18521 22389 18555 22423
rect 18555 22389 18564 22423
rect 18512 22380 18564 22389
rect 21088 22380 21140 22432
rect 26332 22380 26384 22432
rect 32128 22380 32180 22432
rect 34704 22448 34756 22500
rect 34796 22380 34848 22432
rect 39028 22584 39080 22636
rect 39948 22584 40000 22636
rect 40040 22584 40092 22636
rect 43628 22584 43680 22636
rect 46112 22627 46164 22636
rect 46112 22593 46121 22627
rect 46121 22593 46155 22627
rect 46155 22593 46164 22627
rect 46112 22584 46164 22593
rect 39764 22516 39816 22568
rect 45376 22516 45428 22568
rect 47584 22584 47636 22636
rect 35808 22423 35860 22432
rect 35808 22389 35817 22423
rect 35817 22389 35851 22423
rect 35851 22389 35860 22423
rect 35808 22380 35860 22389
rect 41236 22423 41288 22432
rect 41236 22389 41245 22423
rect 41245 22389 41279 22423
rect 41279 22389 41288 22423
rect 41236 22380 41288 22389
rect 46020 22380 46072 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 65654 22278 65706 22330
rect 65718 22278 65770 22330
rect 65782 22278 65834 22330
rect 65846 22278 65898 22330
rect 65910 22278 65962 22330
rect 5356 22176 5408 22228
rect 10692 22176 10744 22228
rect 11060 22176 11112 22228
rect 17224 22176 17276 22228
rect 20904 22219 20956 22228
rect 20904 22185 20913 22219
rect 20913 22185 20947 22219
rect 20947 22185 20956 22219
rect 20904 22176 20956 22185
rect 21548 22219 21600 22228
rect 21548 22185 21557 22219
rect 21557 22185 21591 22219
rect 21591 22185 21600 22219
rect 21548 22176 21600 22185
rect 24308 22176 24360 22228
rect 27436 22219 27488 22228
rect 14004 22108 14056 22160
rect 15384 22108 15436 22160
rect 6644 22040 6696 22092
rect 11520 22040 11572 22092
rect 11612 22040 11664 22092
rect 13820 22040 13872 22092
rect 16488 22108 16540 22160
rect 16764 22108 16816 22160
rect 20720 22108 20772 22160
rect 27436 22185 27445 22219
rect 27445 22185 27479 22219
rect 27479 22185 27488 22219
rect 27436 22176 27488 22185
rect 33692 22176 33744 22228
rect 34704 22219 34756 22228
rect 34704 22185 34713 22219
rect 34713 22185 34747 22219
rect 34747 22185 34756 22219
rect 34704 22176 34756 22185
rect 34888 22219 34940 22228
rect 34888 22185 34897 22219
rect 34897 22185 34931 22219
rect 34931 22185 34940 22219
rect 34888 22176 34940 22185
rect 40040 22219 40092 22228
rect 40040 22185 40049 22219
rect 40049 22185 40083 22219
rect 40083 22185 40092 22219
rect 40040 22176 40092 22185
rect 41236 22176 41288 22228
rect 41880 22176 41932 22228
rect 5816 21972 5868 22024
rect 10048 22015 10100 22024
rect 10048 21981 10057 22015
rect 10057 21981 10091 22015
rect 10091 21981 10100 22015
rect 10048 21972 10100 21981
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 10692 21972 10744 22024
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 16856 21972 16908 22024
rect 8208 21904 8260 21956
rect 16948 21904 17000 21956
rect 17960 22040 18012 22092
rect 18052 22040 18104 22092
rect 20628 21972 20680 22024
rect 21088 21972 21140 22024
rect 21272 21972 21324 22024
rect 21456 21972 21508 22024
rect 22284 22040 22336 22092
rect 24400 22040 24452 22092
rect 29368 22040 29420 22092
rect 29920 22083 29972 22092
rect 29920 22049 29929 22083
rect 29929 22049 29963 22083
rect 29963 22049 29972 22083
rect 29920 22040 29972 22049
rect 30196 22040 30248 22092
rect 31484 22040 31536 22092
rect 22836 22015 22888 22024
rect 22192 21947 22244 21956
rect 22192 21913 22201 21947
rect 22201 21913 22235 21947
rect 22235 21913 22244 21947
rect 22192 21904 22244 21913
rect 22836 21981 22845 22015
rect 22845 21981 22879 22015
rect 22879 21981 22888 22015
rect 22836 21972 22888 21981
rect 23480 21972 23532 22024
rect 24492 21972 24544 22024
rect 26332 22015 26384 22024
rect 26332 21981 26366 22015
rect 26366 21981 26384 22015
rect 26332 21972 26384 21981
rect 29644 21972 29696 22024
rect 29828 22015 29880 22024
rect 29828 21981 29837 22015
rect 29837 21981 29871 22015
rect 29871 21981 29880 22015
rect 31944 22015 31996 22024
rect 29828 21972 29880 21981
rect 31944 21981 31953 22015
rect 31953 21981 31987 22015
rect 31987 21981 31996 22015
rect 31944 21972 31996 21981
rect 32220 22015 32272 22024
rect 24676 21904 24728 21956
rect 25504 21904 25556 21956
rect 9772 21836 9824 21888
rect 14188 21879 14240 21888
rect 14188 21845 14197 21879
rect 14197 21845 14231 21879
rect 14231 21845 14240 21879
rect 14188 21836 14240 21845
rect 15108 21836 15160 21888
rect 16764 21879 16816 21888
rect 16764 21845 16773 21879
rect 16773 21845 16807 21879
rect 16807 21845 16816 21879
rect 16764 21836 16816 21845
rect 18328 21836 18380 21888
rect 18604 21879 18656 21888
rect 18604 21845 18613 21879
rect 18613 21845 18647 21879
rect 18647 21845 18656 21879
rect 18604 21836 18656 21845
rect 24308 21836 24360 21888
rect 26424 21836 26476 21888
rect 31852 21904 31904 21956
rect 32220 21981 32229 22015
rect 32229 21981 32263 22015
rect 32263 21981 32272 22015
rect 32220 21972 32272 21981
rect 32404 21972 32456 22024
rect 34796 21972 34848 22024
rect 32128 21904 32180 21956
rect 35440 21904 35492 21956
rect 36728 21972 36780 22024
rect 37832 22015 37884 22024
rect 37832 21981 37841 22015
rect 37841 21981 37875 22015
rect 37875 21981 37884 22015
rect 37832 21972 37884 21981
rect 38292 21972 38344 22024
rect 39856 22015 39908 22024
rect 39856 21981 39865 22015
rect 39865 21981 39899 22015
rect 39899 21981 39908 22015
rect 39856 21972 39908 21981
rect 40500 22040 40552 22092
rect 46112 22040 46164 22092
rect 41880 21904 41932 21956
rect 37372 21879 37424 21888
rect 37372 21845 37381 21879
rect 37381 21845 37415 21879
rect 37415 21845 37424 21879
rect 37372 21836 37424 21845
rect 37740 21879 37792 21888
rect 37740 21845 37749 21879
rect 37749 21845 37783 21879
rect 37783 21845 37792 21879
rect 37740 21836 37792 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 5356 21632 5408 21684
rect 5816 21675 5868 21684
rect 5816 21641 5825 21675
rect 5825 21641 5859 21675
rect 5859 21641 5868 21675
rect 5816 21632 5868 21641
rect 5908 21632 5960 21684
rect 20260 21632 20312 21684
rect 20812 21632 20864 21684
rect 21272 21675 21324 21684
rect 21272 21641 21281 21675
rect 21281 21641 21315 21675
rect 21315 21641 21324 21675
rect 21272 21632 21324 21641
rect 21824 21632 21876 21684
rect 23664 21632 23716 21684
rect 26240 21632 26292 21684
rect 27160 21632 27212 21684
rect 7104 21539 7156 21548
rect 7104 21505 7113 21539
rect 7113 21505 7147 21539
rect 7147 21505 7156 21539
rect 7104 21496 7156 21505
rect 7932 21539 7984 21548
rect 7932 21505 7941 21539
rect 7941 21505 7975 21539
rect 7975 21505 7984 21539
rect 7932 21496 7984 21505
rect 8208 21539 8260 21548
rect 8208 21505 8217 21539
rect 8217 21505 8251 21539
rect 8251 21505 8260 21539
rect 8208 21496 8260 21505
rect 10048 21539 10100 21548
rect 10048 21505 10057 21539
rect 10057 21505 10091 21539
rect 10091 21505 10100 21539
rect 10048 21496 10100 21505
rect 10232 21539 10284 21548
rect 10232 21505 10241 21539
rect 10241 21505 10275 21539
rect 10275 21505 10284 21539
rect 10232 21496 10284 21505
rect 10784 21539 10836 21548
rect 10784 21505 10793 21539
rect 10793 21505 10827 21539
rect 10827 21505 10836 21539
rect 10784 21496 10836 21505
rect 11520 21539 11572 21548
rect 7012 21428 7064 21480
rect 8944 21471 8996 21480
rect 8944 21437 8953 21471
rect 8953 21437 8987 21471
rect 8987 21437 8996 21471
rect 8944 21428 8996 21437
rect 11060 21428 11112 21480
rect 11520 21505 11529 21539
rect 11529 21505 11563 21539
rect 11563 21505 11572 21539
rect 11520 21496 11572 21505
rect 17224 21564 17276 21616
rect 15292 21496 15344 21548
rect 16764 21496 16816 21548
rect 17868 21564 17920 21616
rect 18512 21564 18564 21616
rect 20352 21496 20404 21548
rect 21088 21564 21140 21616
rect 21180 21564 21232 21616
rect 21364 21564 21416 21616
rect 12532 21428 12584 21480
rect 5448 21360 5500 21412
rect 7564 21360 7616 21412
rect 9496 21360 9548 21412
rect 17776 21471 17828 21480
rect 17776 21437 17785 21471
rect 17785 21437 17819 21471
rect 17819 21437 17828 21471
rect 17776 21428 17828 21437
rect 20996 21496 21048 21548
rect 22928 21539 22980 21548
rect 22928 21505 22937 21539
rect 22937 21505 22971 21539
rect 22971 21505 22980 21539
rect 22928 21496 22980 21505
rect 21180 21428 21232 21480
rect 25504 21428 25556 21480
rect 25780 21471 25832 21480
rect 25780 21437 25789 21471
rect 25789 21437 25823 21471
rect 25823 21437 25832 21471
rect 25780 21428 25832 21437
rect 26056 21496 26108 21548
rect 26700 21496 26752 21548
rect 27160 21496 27212 21548
rect 27804 21496 27856 21548
rect 29644 21539 29696 21548
rect 29644 21505 29653 21539
rect 29653 21505 29687 21539
rect 29687 21505 29696 21539
rect 29644 21496 29696 21505
rect 29920 21632 29972 21684
rect 30288 21632 30340 21684
rect 30380 21632 30432 21684
rect 29828 21564 29880 21616
rect 29920 21539 29972 21548
rect 29920 21505 29929 21539
rect 29929 21505 29963 21539
rect 29963 21505 29972 21539
rect 29920 21496 29972 21505
rect 35532 21607 35584 21616
rect 35532 21573 35541 21607
rect 35541 21573 35575 21607
rect 35575 21573 35584 21607
rect 35532 21564 35584 21573
rect 45836 21564 45888 21616
rect 30748 21539 30800 21548
rect 30748 21505 30757 21539
rect 30757 21505 30791 21539
rect 30791 21505 30800 21539
rect 30748 21496 30800 21505
rect 32312 21539 32364 21548
rect 32312 21505 32321 21539
rect 32321 21505 32355 21539
rect 32355 21505 32364 21539
rect 32312 21496 32364 21505
rect 32404 21539 32456 21548
rect 32404 21505 32413 21539
rect 32413 21505 32447 21539
rect 32447 21505 32456 21539
rect 32404 21496 32456 21505
rect 35716 21496 35768 21548
rect 36728 21539 36780 21548
rect 36728 21505 36737 21539
rect 36737 21505 36771 21539
rect 36771 21505 36780 21539
rect 36728 21496 36780 21505
rect 38108 21496 38160 21548
rect 44272 21539 44324 21548
rect 44272 21505 44281 21539
rect 44281 21505 44315 21539
rect 44315 21505 44324 21539
rect 44272 21496 44324 21505
rect 46020 21539 46072 21548
rect 46020 21505 46029 21539
rect 46029 21505 46063 21539
rect 46063 21505 46072 21539
rect 46020 21496 46072 21505
rect 46848 21539 46900 21548
rect 46848 21505 46857 21539
rect 46857 21505 46891 21539
rect 46891 21505 46900 21539
rect 46848 21496 46900 21505
rect 32680 21471 32732 21480
rect 28448 21403 28500 21412
rect 7380 21335 7432 21344
rect 7380 21301 7389 21335
rect 7389 21301 7423 21335
rect 7423 21301 7432 21335
rect 7380 21292 7432 21301
rect 8392 21335 8444 21344
rect 8392 21301 8401 21335
rect 8401 21301 8435 21335
rect 8435 21301 8444 21335
rect 8392 21292 8444 21301
rect 9404 21292 9456 21344
rect 14740 21292 14792 21344
rect 16856 21335 16908 21344
rect 16856 21301 16865 21335
rect 16865 21301 16899 21335
rect 16899 21301 16908 21335
rect 16856 21292 16908 21301
rect 16948 21292 17000 21344
rect 28448 21369 28457 21403
rect 28457 21369 28491 21403
rect 28491 21369 28500 21403
rect 28448 21360 28500 21369
rect 32680 21437 32689 21471
rect 32689 21437 32723 21471
rect 32723 21437 32732 21471
rect 32680 21428 32732 21437
rect 32772 21471 32824 21480
rect 32772 21437 32781 21471
rect 32781 21437 32815 21471
rect 32815 21437 32824 21471
rect 35256 21471 35308 21480
rect 32772 21428 32824 21437
rect 35256 21437 35265 21471
rect 35265 21437 35299 21471
rect 35299 21437 35308 21471
rect 35256 21428 35308 21437
rect 35440 21471 35492 21480
rect 35440 21437 35449 21471
rect 35449 21437 35483 21471
rect 35483 21437 35492 21471
rect 35440 21428 35492 21437
rect 37372 21428 37424 21480
rect 43812 21428 43864 21480
rect 31852 21360 31904 21412
rect 31944 21360 31996 21412
rect 32864 21360 32916 21412
rect 37556 21360 37608 21412
rect 18972 21292 19024 21344
rect 20168 21292 20220 21344
rect 20904 21292 20956 21344
rect 21824 21335 21876 21344
rect 21824 21301 21833 21335
rect 21833 21301 21867 21335
rect 21867 21301 21876 21335
rect 21824 21292 21876 21301
rect 24492 21292 24544 21344
rect 24768 21292 24820 21344
rect 27804 21335 27856 21344
rect 27804 21301 27813 21335
rect 27813 21301 27847 21335
rect 27847 21301 27856 21335
rect 27804 21292 27856 21301
rect 28540 21292 28592 21344
rect 30472 21292 30524 21344
rect 34612 21292 34664 21344
rect 34888 21292 34940 21344
rect 36268 21292 36320 21344
rect 37740 21292 37792 21344
rect 39856 21292 39908 21344
rect 42340 21292 42392 21344
rect 43904 21292 43956 21344
rect 45008 21292 45060 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 65654 21190 65706 21242
rect 65718 21190 65770 21242
rect 65782 21190 65834 21242
rect 65846 21190 65898 21242
rect 65910 21190 65962 21242
rect 8944 21088 8996 21140
rect 10784 21088 10836 21140
rect 11704 21088 11756 21140
rect 7012 21020 7064 21072
rect 6644 20952 6696 21004
rect 6920 20952 6972 21004
rect 6276 20859 6328 20868
rect 6276 20825 6294 20859
rect 6294 20825 6328 20859
rect 6276 20816 6328 20825
rect 7104 20816 7156 20868
rect 7564 20995 7616 21004
rect 7564 20961 7573 20995
rect 7573 20961 7607 20995
rect 7607 20961 7616 20995
rect 7564 20952 7616 20961
rect 8300 20952 8352 21004
rect 8208 20884 8260 20936
rect 9404 20927 9456 20936
rect 9404 20893 9413 20927
rect 9413 20893 9447 20927
rect 9447 20893 9456 20927
rect 11060 20952 11112 21004
rect 14280 21088 14332 21140
rect 9404 20884 9456 20893
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 11244 20884 11296 20936
rect 9496 20859 9548 20868
rect 7012 20791 7064 20800
rect 7012 20757 7021 20791
rect 7021 20757 7055 20791
rect 7055 20757 7064 20791
rect 7012 20748 7064 20757
rect 9220 20748 9272 20800
rect 9496 20825 9505 20859
rect 9505 20825 9539 20859
rect 9539 20825 9548 20859
rect 9496 20816 9548 20825
rect 11612 20748 11664 20800
rect 12256 20952 12308 21004
rect 13912 20952 13964 21004
rect 14464 20995 14516 21004
rect 14464 20961 14473 20995
rect 14473 20961 14507 20995
rect 14507 20961 14516 20995
rect 14464 20952 14516 20961
rect 12532 20884 12584 20936
rect 14740 20927 14792 20936
rect 14740 20893 14774 20927
rect 14774 20893 14792 20927
rect 14740 20884 14792 20893
rect 15016 20884 15068 20936
rect 13544 20816 13596 20868
rect 16028 20816 16080 20868
rect 14188 20748 14240 20800
rect 15844 20791 15896 20800
rect 15844 20757 15853 20791
rect 15853 20757 15887 20791
rect 15887 20757 15896 20791
rect 15844 20748 15896 20757
rect 16948 21088 17000 21140
rect 17960 21088 18012 21140
rect 20168 21088 20220 21140
rect 21180 21088 21232 21140
rect 23572 21131 23624 21140
rect 23572 21097 23581 21131
rect 23581 21097 23615 21131
rect 23615 21097 23624 21131
rect 23572 21088 23624 21097
rect 24492 21088 24544 21140
rect 25596 21088 25648 21140
rect 28448 21131 28500 21140
rect 28448 21097 28457 21131
rect 28457 21097 28491 21131
rect 28491 21097 28500 21131
rect 28448 21088 28500 21097
rect 25044 21063 25096 21072
rect 25044 21029 25053 21063
rect 25053 21029 25087 21063
rect 25087 21029 25096 21063
rect 25044 21020 25096 21029
rect 29920 21088 29972 21140
rect 30748 21088 30800 21140
rect 32680 21088 32732 21140
rect 35716 21131 35768 21140
rect 35716 21097 35725 21131
rect 35725 21097 35759 21131
rect 35759 21097 35768 21131
rect 35716 21088 35768 21097
rect 40132 21088 40184 21140
rect 41880 21088 41932 21140
rect 18880 20952 18932 21004
rect 19432 20952 19484 21004
rect 20904 20952 20956 21004
rect 31852 21020 31904 21072
rect 16856 20884 16908 20936
rect 17868 20884 17920 20936
rect 20812 20927 20864 20936
rect 18052 20816 18104 20868
rect 20812 20893 20821 20927
rect 20821 20893 20855 20927
rect 20855 20893 20864 20927
rect 20812 20884 20864 20893
rect 22284 20884 22336 20936
rect 25780 20884 25832 20936
rect 25964 20927 26016 20936
rect 25964 20893 25973 20927
rect 25973 20893 26007 20927
rect 26007 20893 26016 20927
rect 29552 20952 29604 21004
rect 25964 20884 26016 20893
rect 28448 20884 28500 20936
rect 21364 20816 21416 20868
rect 22468 20859 22520 20868
rect 22468 20825 22502 20859
rect 22502 20825 22520 20859
rect 24768 20859 24820 20868
rect 22468 20816 22520 20825
rect 24768 20825 24777 20859
rect 24777 20825 24811 20859
rect 24811 20825 24820 20859
rect 24768 20816 24820 20825
rect 18788 20748 18840 20800
rect 18972 20748 19024 20800
rect 22928 20748 22980 20800
rect 28540 20816 28592 20868
rect 26424 20791 26476 20800
rect 26424 20757 26433 20791
rect 26433 20757 26467 20791
rect 26467 20757 26476 20791
rect 26424 20748 26476 20757
rect 29368 20748 29420 20800
rect 30104 20884 30156 20936
rect 32496 20952 32548 21004
rect 33508 20995 33560 21004
rect 33508 20961 33517 20995
rect 33517 20961 33551 20995
rect 33551 20961 33560 20995
rect 33508 20952 33560 20961
rect 35440 21020 35492 21072
rect 42432 21020 42484 21072
rect 37832 20952 37884 21004
rect 39948 20995 40000 21004
rect 39948 20961 39957 20995
rect 39957 20961 39991 20995
rect 39991 20961 40000 20995
rect 39948 20952 40000 20961
rect 42616 20952 42668 21004
rect 46112 21088 46164 21140
rect 32220 20927 32272 20936
rect 32220 20893 32229 20927
rect 32229 20893 32263 20927
rect 32263 20893 32272 20927
rect 32220 20884 32272 20893
rect 30288 20816 30340 20868
rect 32864 20884 32916 20936
rect 37280 20859 37332 20868
rect 37280 20825 37298 20859
rect 37298 20825 37332 20859
rect 37280 20816 37332 20825
rect 37740 20884 37792 20936
rect 39856 20927 39908 20936
rect 39304 20816 39356 20868
rect 39856 20893 39865 20927
rect 39865 20893 39899 20927
rect 39899 20893 39908 20927
rect 39856 20884 39908 20893
rect 40132 20927 40184 20936
rect 40132 20893 40141 20927
rect 40141 20893 40175 20927
rect 40175 20893 40184 20927
rect 40132 20884 40184 20893
rect 42340 20884 42392 20936
rect 41236 20816 41288 20868
rect 35624 20748 35676 20800
rect 38016 20791 38068 20800
rect 38016 20757 38025 20791
rect 38025 20757 38059 20791
rect 38059 20757 38068 20791
rect 38016 20748 38068 20757
rect 41604 20748 41656 20800
rect 42800 20884 42852 20936
rect 45008 20927 45060 20936
rect 45008 20893 45017 20927
rect 45017 20893 45051 20927
rect 45051 20893 45060 20927
rect 45008 20884 45060 20893
rect 45652 20927 45704 20936
rect 45652 20893 45661 20927
rect 45661 20893 45695 20927
rect 45695 20893 45704 20927
rect 45652 20884 45704 20893
rect 42708 20748 42760 20800
rect 42800 20748 42852 20800
rect 44180 20791 44232 20800
rect 44180 20757 44189 20791
rect 44189 20757 44223 20791
rect 44223 20757 44232 20791
rect 44180 20748 44232 20757
rect 45192 20791 45244 20800
rect 45192 20757 45201 20791
rect 45201 20757 45235 20791
rect 45235 20757 45244 20791
rect 45192 20748 45244 20757
rect 46112 20748 46164 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 6276 20544 6328 20596
rect 9128 20544 9180 20596
rect 11244 20544 11296 20596
rect 11612 20544 11664 20596
rect 12348 20544 12400 20596
rect 14004 20544 14056 20596
rect 14188 20476 14240 20528
rect 15200 20476 15252 20528
rect 16948 20544 17000 20596
rect 17132 20587 17184 20596
rect 17132 20553 17141 20587
rect 17141 20553 17175 20587
rect 17175 20553 17184 20587
rect 17132 20544 17184 20553
rect 18788 20544 18840 20596
rect 15844 20476 15896 20528
rect 7012 20408 7064 20460
rect 8392 20408 8444 20460
rect 7380 20383 7432 20392
rect 7380 20349 7389 20383
rect 7389 20349 7423 20383
rect 7423 20349 7432 20383
rect 7380 20340 7432 20349
rect 8208 20340 8260 20392
rect 9036 20451 9088 20460
rect 9036 20417 9045 20451
rect 9045 20417 9079 20451
rect 9079 20417 9088 20451
rect 9220 20451 9272 20460
rect 9036 20408 9088 20417
rect 9220 20417 9229 20451
rect 9229 20417 9263 20451
rect 9263 20417 9272 20451
rect 9220 20408 9272 20417
rect 10324 20451 10376 20460
rect 10324 20417 10333 20451
rect 10333 20417 10367 20451
rect 10367 20417 10376 20451
rect 10324 20408 10376 20417
rect 11980 20408 12032 20460
rect 15476 20408 15528 20460
rect 9312 20340 9364 20392
rect 12164 20340 12216 20392
rect 9220 20272 9272 20324
rect 15292 20315 15344 20324
rect 15292 20281 15301 20315
rect 15301 20281 15335 20315
rect 15335 20281 15344 20315
rect 15292 20272 15344 20281
rect 15844 20383 15896 20392
rect 15844 20349 15853 20383
rect 15853 20349 15887 20383
rect 15887 20349 15896 20383
rect 15844 20340 15896 20349
rect 18880 20408 18932 20460
rect 19432 20476 19484 20528
rect 20720 20544 20772 20596
rect 23572 20544 23624 20596
rect 25780 20544 25832 20596
rect 28264 20587 28316 20596
rect 28264 20553 28273 20587
rect 28273 20553 28307 20587
rect 28307 20553 28316 20587
rect 28264 20544 28316 20553
rect 29368 20587 29420 20596
rect 29368 20553 29377 20587
rect 29377 20553 29411 20587
rect 29411 20553 29420 20587
rect 29368 20544 29420 20553
rect 31300 20544 31352 20596
rect 32772 20544 32824 20596
rect 20996 20476 21048 20528
rect 22100 20476 22152 20528
rect 18512 20340 18564 20392
rect 19156 20340 19208 20392
rect 22192 20340 22244 20392
rect 22836 20383 22888 20392
rect 22836 20349 22845 20383
rect 22845 20349 22879 20383
rect 22879 20349 22888 20383
rect 22836 20340 22888 20349
rect 16764 20272 16816 20324
rect 18144 20272 18196 20324
rect 5540 20247 5592 20256
rect 5540 20213 5549 20247
rect 5549 20213 5583 20247
rect 5583 20213 5592 20247
rect 5540 20204 5592 20213
rect 10600 20204 10652 20256
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 14832 20247 14884 20256
rect 14832 20213 14841 20247
rect 14841 20213 14875 20247
rect 14875 20213 14884 20247
rect 14832 20204 14884 20213
rect 16120 20204 16172 20256
rect 16948 20204 17000 20256
rect 19892 20272 19944 20324
rect 20904 20272 20956 20324
rect 19248 20247 19300 20256
rect 19248 20213 19257 20247
rect 19257 20213 19291 20247
rect 19291 20213 19300 20247
rect 19248 20204 19300 20213
rect 19340 20204 19392 20256
rect 22284 20247 22336 20256
rect 22284 20213 22293 20247
rect 22293 20213 22327 20247
rect 22327 20213 22336 20247
rect 22284 20204 22336 20213
rect 23388 20204 23440 20256
rect 24768 20408 24820 20460
rect 26424 20476 26476 20528
rect 32220 20476 32272 20528
rect 33600 20476 33652 20528
rect 37280 20544 37332 20596
rect 40132 20544 40184 20596
rect 41236 20587 41288 20596
rect 41236 20553 41245 20587
rect 41245 20553 41279 20587
rect 41279 20553 41288 20587
rect 41236 20544 41288 20553
rect 37556 20476 37608 20528
rect 29644 20408 29696 20460
rect 30104 20408 30156 20460
rect 32496 20451 32548 20460
rect 32496 20417 32505 20451
rect 32505 20417 32539 20451
rect 32539 20417 32548 20451
rect 32496 20408 32548 20417
rect 33784 20451 33836 20460
rect 33784 20417 33793 20451
rect 33793 20417 33827 20451
rect 33827 20417 33836 20451
rect 33784 20408 33836 20417
rect 36268 20451 36320 20460
rect 36268 20417 36277 20451
rect 36277 20417 36311 20451
rect 36311 20417 36320 20451
rect 36268 20408 36320 20417
rect 40040 20451 40092 20460
rect 40040 20417 40049 20451
rect 40049 20417 40083 20451
rect 40083 20417 40092 20451
rect 40040 20408 40092 20417
rect 40316 20451 40368 20460
rect 25964 20340 26016 20392
rect 27344 20340 27396 20392
rect 29828 20383 29880 20392
rect 29828 20349 29837 20383
rect 29837 20349 29871 20383
rect 29871 20349 29880 20383
rect 29828 20340 29880 20349
rect 33508 20340 33560 20392
rect 39304 20340 39356 20392
rect 40316 20417 40325 20451
rect 40325 20417 40359 20451
rect 40359 20417 40368 20451
rect 40316 20408 40368 20417
rect 40408 20451 40460 20460
rect 40408 20417 40417 20451
rect 40417 20417 40451 20451
rect 40451 20417 40460 20451
rect 40408 20408 40460 20417
rect 42616 20544 42668 20596
rect 43812 20476 43864 20528
rect 44180 20476 44232 20528
rect 42432 20451 42484 20460
rect 42432 20417 42441 20451
rect 42441 20417 42475 20451
rect 42475 20417 42484 20451
rect 42432 20408 42484 20417
rect 42708 20451 42760 20460
rect 42708 20417 42717 20451
rect 42717 20417 42751 20451
rect 42751 20417 42760 20451
rect 42708 20408 42760 20417
rect 45008 20408 45060 20460
rect 45192 20408 45244 20460
rect 46112 20451 46164 20460
rect 46112 20417 46121 20451
rect 46121 20417 46155 20451
rect 46155 20417 46164 20451
rect 46112 20408 46164 20417
rect 24952 20204 25004 20256
rect 25780 20247 25832 20256
rect 25780 20213 25789 20247
rect 25789 20213 25823 20247
rect 25823 20213 25832 20247
rect 25780 20204 25832 20213
rect 27804 20204 27856 20256
rect 28448 20204 28500 20256
rect 35808 20247 35860 20256
rect 35808 20213 35817 20247
rect 35817 20213 35851 20247
rect 35851 20213 35860 20247
rect 35808 20204 35860 20213
rect 41420 20204 41472 20256
rect 41604 20272 41656 20324
rect 43352 20340 43404 20392
rect 44272 20340 44324 20392
rect 44916 20340 44968 20392
rect 43076 20204 43128 20256
rect 45192 20204 45244 20256
rect 55128 20204 55180 20256
rect 60556 20204 60608 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 65654 20102 65706 20154
rect 65718 20102 65770 20154
rect 65782 20102 65834 20154
rect 65846 20102 65898 20154
rect 65910 20102 65962 20154
rect 7932 20000 7984 20052
rect 11980 20043 12032 20052
rect 11980 20009 11989 20043
rect 11989 20009 12023 20043
rect 12023 20009 12032 20043
rect 11980 20000 12032 20009
rect 12164 20000 12216 20052
rect 22192 20000 22244 20052
rect 22468 20043 22520 20052
rect 22468 20009 22477 20043
rect 22477 20009 22511 20043
rect 22511 20009 22520 20043
rect 22468 20000 22520 20009
rect 23756 20000 23808 20052
rect 27344 20043 27396 20052
rect 27344 20009 27353 20043
rect 27353 20009 27387 20043
rect 27387 20009 27396 20043
rect 27344 20000 27396 20009
rect 31668 20000 31720 20052
rect 33784 20000 33836 20052
rect 5724 19864 5776 19916
rect 5540 19796 5592 19848
rect 7104 19796 7156 19848
rect 8300 19932 8352 19984
rect 14188 19975 14240 19984
rect 14188 19941 14197 19975
rect 14197 19941 14231 19975
rect 14231 19941 14240 19975
rect 14188 19932 14240 19941
rect 17132 19975 17184 19984
rect 8484 19864 8536 19916
rect 11152 19864 11204 19916
rect 12256 19864 12308 19916
rect 14464 19864 14516 19916
rect 17132 19941 17141 19975
rect 17141 19941 17175 19975
rect 17175 19941 17184 19975
rect 17132 19932 17184 19941
rect 18052 19975 18104 19984
rect 18052 19941 18061 19975
rect 18061 19941 18095 19975
rect 18095 19941 18104 19975
rect 18052 19932 18104 19941
rect 18788 19932 18840 19984
rect 8208 19796 8260 19848
rect 9496 19796 9548 19848
rect 4620 19728 4672 19780
rect 11520 19796 11572 19848
rect 12348 19796 12400 19848
rect 14832 19839 14884 19848
rect 14832 19805 14841 19839
rect 14841 19805 14875 19839
rect 14875 19805 14884 19839
rect 14832 19796 14884 19805
rect 18512 19839 18564 19848
rect 18512 19805 18521 19839
rect 18521 19805 18555 19839
rect 18555 19805 18564 19839
rect 18512 19796 18564 19805
rect 10784 19728 10836 19780
rect 15936 19728 15988 19780
rect 19156 19796 19208 19848
rect 19984 19864 20036 19916
rect 5448 19660 5500 19712
rect 6552 19703 6604 19712
rect 6552 19669 6561 19703
rect 6561 19669 6595 19703
rect 6595 19669 6604 19703
rect 6552 19660 6604 19669
rect 7104 19703 7156 19712
rect 7104 19669 7113 19703
rect 7113 19669 7147 19703
rect 7147 19669 7156 19703
rect 7104 19660 7156 19669
rect 9036 19660 9088 19712
rect 9312 19703 9364 19712
rect 9312 19669 9321 19703
rect 9321 19669 9355 19703
rect 9355 19669 9364 19703
rect 9312 19660 9364 19669
rect 11060 19660 11112 19712
rect 14648 19703 14700 19712
rect 14648 19669 14657 19703
rect 14657 19669 14691 19703
rect 14691 19669 14700 19703
rect 14648 19660 14700 19669
rect 15476 19660 15528 19712
rect 18880 19728 18932 19780
rect 19524 19728 19576 19780
rect 18696 19703 18748 19712
rect 18696 19669 18705 19703
rect 18705 19669 18739 19703
rect 18739 19669 18748 19703
rect 18696 19660 18748 19669
rect 19432 19703 19484 19712
rect 19432 19669 19441 19703
rect 19441 19669 19475 19703
rect 19475 19669 19484 19703
rect 19432 19660 19484 19669
rect 19800 19796 19852 19848
rect 20812 19932 20864 19984
rect 20904 19932 20956 19984
rect 26056 19975 26108 19984
rect 26056 19941 26065 19975
rect 26065 19941 26099 19975
rect 26099 19941 26108 19975
rect 26056 19932 26108 19941
rect 25780 19907 25832 19916
rect 25780 19873 25789 19907
rect 25789 19873 25823 19907
rect 25823 19873 25832 19907
rect 25780 19864 25832 19873
rect 22284 19839 22336 19848
rect 22284 19805 22293 19839
rect 22293 19805 22327 19839
rect 22327 19805 22336 19839
rect 22284 19796 22336 19805
rect 23020 19796 23072 19848
rect 26240 19796 26292 19848
rect 32496 19932 32548 19984
rect 27160 19907 27212 19916
rect 27160 19873 27169 19907
rect 27169 19873 27203 19907
rect 27203 19873 27212 19907
rect 27160 19864 27212 19873
rect 27344 19864 27396 19916
rect 29276 19864 29328 19916
rect 29828 19864 29880 19916
rect 37924 20000 37976 20052
rect 40040 20043 40092 20052
rect 40040 20009 40049 20043
rect 40049 20009 40083 20043
rect 40083 20009 40092 20043
rect 40040 20000 40092 20009
rect 41420 20043 41472 20052
rect 41420 20009 41429 20043
rect 41429 20009 41463 20043
rect 41463 20009 41472 20043
rect 41420 20000 41472 20009
rect 42708 20000 42760 20052
rect 45652 20000 45704 20052
rect 39948 19932 40000 19984
rect 35440 19907 35492 19916
rect 35440 19873 35449 19907
rect 35449 19873 35483 19907
rect 35483 19873 35492 19907
rect 35440 19864 35492 19873
rect 38016 19864 38068 19916
rect 40316 19932 40368 19984
rect 43812 19932 43864 19984
rect 45100 19932 45152 19984
rect 42800 19907 42852 19916
rect 42800 19873 42809 19907
rect 42809 19873 42843 19907
rect 42843 19873 42852 19907
rect 42800 19864 42852 19873
rect 44916 19864 44968 19916
rect 30104 19839 30156 19848
rect 30104 19805 30113 19839
rect 30113 19805 30147 19839
rect 30147 19805 30156 19839
rect 30104 19796 30156 19805
rect 19892 19728 19944 19780
rect 33324 19796 33376 19848
rect 35808 19796 35860 19848
rect 40408 19796 40460 19848
rect 43076 19839 43128 19848
rect 43076 19805 43085 19839
rect 43085 19805 43119 19839
rect 43119 19805 43128 19839
rect 43076 19796 43128 19805
rect 35532 19728 35584 19780
rect 40592 19771 40644 19780
rect 40592 19737 40601 19771
rect 40601 19737 40635 19771
rect 40635 19737 40644 19771
rect 40592 19728 40644 19737
rect 40684 19771 40736 19780
rect 40684 19737 40693 19771
rect 40693 19737 40727 19771
rect 40727 19737 40736 19771
rect 40684 19728 40736 19737
rect 41144 19728 41196 19780
rect 42432 19728 42484 19780
rect 20076 19660 20128 19712
rect 20628 19703 20680 19712
rect 20628 19669 20637 19703
rect 20637 19669 20671 19703
rect 20671 19669 20680 19703
rect 20628 19660 20680 19669
rect 31116 19703 31168 19712
rect 31116 19669 31125 19703
rect 31125 19669 31159 19703
rect 31159 19669 31168 19703
rect 31116 19660 31168 19669
rect 32496 19660 32548 19712
rect 43628 19660 43680 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 5724 19499 5776 19508
rect 5724 19465 5733 19499
rect 5733 19465 5767 19499
rect 5767 19465 5776 19499
rect 5724 19456 5776 19465
rect 15476 19499 15528 19508
rect 7104 19388 7156 19440
rect 15476 19465 15485 19499
rect 15485 19465 15519 19499
rect 15519 19465 15528 19499
rect 15476 19456 15528 19465
rect 15936 19499 15988 19508
rect 15936 19465 15945 19499
rect 15945 19465 15979 19499
rect 15979 19465 15988 19499
rect 15936 19456 15988 19465
rect 14648 19388 14700 19440
rect 4436 19320 4488 19372
rect 6552 19320 6604 19372
rect 7380 19363 7432 19372
rect 7380 19329 7389 19363
rect 7389 19329 7423 19363
rect 7423 19329 7432 19363
rect 7380 19320 7432 19329
rect 5724 19184 5776 19236
rect 8300 19320 8352 19372
rect 11060 19320 11112 19372
rect 11520 19320 11572 19372
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 18788 19363 18840 19372
rect 18788 19329 18797 19363
rect 18797 19329 18831 19363
rect 18831 19329 18840 19363
rect 18788 19320 18840 19329
rect 20628 19456 20680 19508
rect 23664 19456 23716 19508
rect 30380 19456 30432 19508
rect 31760 19456 31812 19508
rect 33600 19499 33652 19508
rect 33600 19465 33609 19499
rect 33609 19465 33643 19499
rect 33643 19465 33652 19499
rect 33600 19456 33652 19465
rect 40684 19456 40736 19508
rect 45100 19499 45152 19508
rect 45100 19465 45109 19499
rect 45109 19465 45143 19499
rect 45143 19465 45152 19499
rect 45100 19456 45152 19465
rect 19432 19388 19484 19440
rect 19984 19388 20036 19440
rect 20996 19388 21048 19440
rect 22928 19388 22980 19440
rect 9588 19252 9640 19304
rect 10600 19295 10652 19304
rect 10600 19261 10609 19295
rect 10609 19261 10643 19295
rect 10643 19261 10652 19295
rect 10600 19252 10652 19261
rect 16764 19295 16816 19304
rect 4988 19116 5040 19168
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 20076 19320 20128 19372
rect 21180 19320 21232 19372
rect 25228 19388 25280 19440
rect 33508 19388 33560 19440
rect 39304 19388 39356 19440
rect 43628 19431 43680 19440
rect 23388 19363 23440 19372
rect 23388 19329 23397 19363
rect 23397 19329 23431 19363
rect 23431 19329 23440 19363
rect 23388 19320 23440 19329
rect 24400 19363 24452 19372
rect 24400 19329 24409 19363
rect 24409 19329 24443 19363
rect 24443 19329 24452 19363
rect 24400 19320 24452 19329
rect 24676 19363 24728 19372
rect 24676 19329 24710 19363
rect 24710 19329 24728 19363
rect 24676 19320 24728 19329
rect 32036 19320 32088 19372
rect 32220 19363 32272 19372
rect 32220 19329 32229 19363
rect 32229 19329 32263 19363
rect 32263 19329 32272 19363
rect 32220 19320 32272 19329
rect 32496 19363 32548 19372
rect 32496 19329 32530 19363
rect 32530 19329 32548 19363
rect 32496 19320 32548 19329
rect 38844 19320 38896 19372
rect 39672 19363 39724 19372
rect 39672 19329 39681 19363
rect 39681 19329 39715 19363
rect 39715 19329 39724 19363
rect 39672 19320 39724 19329
rect 21088 19295 21140 19304
rect 21088 19261 21097 19295
rect 21097 19261 21131 19295
rect 21131 19261 21140 19295
rect 21088 19252 21140 19261
rect 23020 19252 23072 19304
rect 39212 19252 39264 19304
rect 39764 19295 39816 19304
rect 39764 19261 39773 19295
rect 39773 19261 39807 19295
rect 39807 19261 39816 19295
rect 39764 19252 39816 19261
rect 40132 19320 40184 19372
rect 40684 19363 40736 19372
rect 40684 19329 40693 19363
rect 40693 19329 40727 19363
rect 40727 19329 40736 19363
rect 40684 19320 40736 19329
rect 43628 19397 43637 19431
rect 43637 19397 43671 19431
rect 43671 19397 43680 19431
rect 43628 19388 43680 19397
rect 44272 19388 44324 19440
rect 43352 19363 43404 19372
rect 43352 19329 43361 19363
rect 43361 19329 43395 19363
rect 43395 19329 43404 19363
rect 43352 19320 43404 19329
rect 20812 19184 20864 19236
rect 20904 19184 20956 19236
rect 24308 19184 24360 19236
rect 18880 19159 18932 19168
rect 18880 19125 18889 19159
rect 18889 19125 18923 19159
rect 18923 19125 18932 19159
rect 18880 19116 18932 19125
rect 19432 19116 19484 19168
rect 20352 19116 20404 19168
rect 20536 19159 20588 19168
rect 20536 19125 20545 19159
rect 20545 19125 20579 19159
rect 20579 19125 20588 19159
rect 20536 19116 20588 19125
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 26240 19159 26292 19168
rect 26240 19125 26249 19159
rect 26249 19125 26283 19159
rect 26283 19125 26292 19159
rect 26240 19116 26292 19125
rect 35440 19116 35492 19168
rect 36452 19116 36504 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 65654 19014 65706 19066
rect 65718 19014 65770 19066
rect 65782 19014 65834 19066
rect 65846 19014 65898 19066
rect 65910 19014 65962 19066
rect 4988 18955 5040 18964
rect 4988 18921 4997 18955
rect 4997 18921 5031 18955
rect 5031 18921 5040 18955
rect 4988 18912 5040 18921
rect 5540 18912 5592 18964
rect 11152 18844 11204 18896
rect 12900 18844 12952 18896
rect 18880 18912 18932 18964
rect 19248 18912 19300 18964
rect 24676 18955 24728 18964
rect 24676 18921 24685 18955
rect 24685 18921 24719 18955
rect 24719 18921 24728 18955
rect 24676 18912 24728 18921
rect 27804 18912 27856 18964
rect 7104 18776 7156 18828
rect 5724 18708 5776 18760
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 16948 18751 17000 18760
rect 16948 18717 16957 18751
rect 16957 18717 16991 18751
rect 16991 18717 17000 18751
rect 16948 18708 17000 18717
rect 10968 18640 11020 18692
rect 6184 18572 6236 18624
rect 6460 18572 6512 18624
rect 7748 18615 7800 18624
rect 7748 18581 7757 18615
rect 7757 18581 7791 18615
rect 7791 18581 7800 18615
rect 7748 18572 7800 18581
rect 10324 18572 10376 18624
rect 11612 18615 11664 18624
rect 11612 18581 11621 18615
rect 11621 18581 11655 18615
rect 11655 18581 11664 18615
rect 11612 18572 11664 18581
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 16396 18640 16448 18692
rect 19340 18776 19392 18828
rect 18696 18708 18748 18760
rect 19156 18708 19208 18760
rect 20536 18751 20588 18760
rect 20536 18717 20545 18751
rect 20545 18717 20579 18751
rect 20579 18717 20588 18751
rect 20536 18708 20588 18717
rect 21272 18708 21324 18760
rect 26424 18844 26476 18896
rect 27252 18844 27304 18896
rect 25780 18819 25832 18828
rect 25780 18785 25789 18819
rect 25789 18785 25823 18819
rect 25823 18785 25832 18819
rect 25780 18776 25832 18785
rect 27068 18776 27120 18828
rect 25412 18708 25464 18760
rect 29368 18912 29420 18964
rect 29644 18912 29696 18964
rect 32588 18912 32640 18964
rect 33324 18955 33376 18964
rect 33324 18921 33333 18955
rect 33333 18921 33367 18955
rect 33367 18921 33376 18955
rect 33324 18912 33376 18921
rect 40592 18912 40644 18964
rect 44272 18955 44324 18964
rect 44272 18921 44281 18955
rect 44281 18921 44315 18955
rect 44315 18921 44324 18955
rect 44272 18912 44324 18921
rect 45008 18912 45060 18964
rect 30104 18844 30156 18896
rect 33600 18776 33652 18828
rect 33876 18819 33928 18828
rect 33876 18785 33885 18819
rect 33885 18785 33919 18819
rect 33919 18785 33928 18819
rect 39304 18819 39356 18828
rect 33876 18776 33928 18785
rect 39304 18785 39313 18819
rect 39313 18785 39347 18819
rect 39347 18785 39356 18819
rect 39304 18776 39356 18785
rect 27252 18708 27304 18760
rect 19340 18640 19392 18692
rect 13544 18572 13596 18624
rect 17132 18615 17184 18624
rect 17132 18581 17141 18615
rect 17141 18581 17175 18615
rect 17175 18581 17184 18615
rect 17132 18572 17184 18581
rect 19984 18572 20036 18624
rect 23020 18640 23072 18692
rect 26240 18640 26292 18692
rect 32220 18708 32272 18760
rect 40132 18751 40184 18760
rect 40132 18717 40141 18751
rect 40141 18717 40175 18751
rect 40175 18717 40184 18751
rect 40132 18708 40184 18717
rect 29184 18640 29236 18692
rect 31116 18640 31168 18692
rect 31760 18683 31812 18692
rect 31760 18649 31794 18683
rect 31794 18649 31812 18683
rect 31760 18640 31812 18649
rect 32496 18640 32548 18692
rect 38016 18640 38068 18692
rect 38844 18640 38896 18692
rect 25688 18615 25740 18624
rect 25688 18581 25697 18615
rect 25697 18581 25731 18615
rect 25731 18581 25740 18615
rect 25688 18572 25740 18581
rect 30196 18572 30248 18624
rect 34520 18572 34572 18624
rect 37924 18615 37976 18624
rect 37924 18581 37933 18615
rect 37933 18581 37967 18615
rect 37967 18581 37976 18615
rect 40684 18708 40736 18760
rect 41880 18708 41932 18760
rect 67824 18751 67876 18760
rect 67824 18717 67833 18751
rect 67833 18717 67867 18751
rect 67867 18717 67876 18751
rect 67824 18708 67876 18717
rect 37924 18572 37976 18581
rect 55128 18572 55180 18624
rect 55772 18572 55824 18624
rect 68008 18615 68060 18624
rect 68008 18581 68017 18615
rect 68017 18581 68051 18615
rect 68051 18581 68060 18615
rect 68008 18572 68060 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 7380 18368 7432 18420
rect 8484 18411 8536 18420
rect 8484 18377 8493 18411
rect 8493 18377 8527 18411
rect 8527 18377 8536 18411
rect 8484 18368 8536 18377
rect 15384 18368 15436 18420
rect 18972 18368 19024 18420
rect 19248 18411 19300 18420
rect 19248 18377 19257 18411
rect 19257 18377 19291 18411
rect 19291 18377 19300 18411
rect 19248 18368 19300 18377
rect 19340 18368 19392 18420
rect 5448 18300 5500 18352
rect 7748 18232 7800 18284
rect 11612 18300 11664 18352
rect 11520 18275 11572 18284
rect 11520 18241 11529 18275
rect 11529 18241 11563 18275
rect 11563 18241 11572 18275
rect 11520 18232 11572 18241
rect 16396 18232 16448 18284
rect 17132 18232 17184 18284
rect 18880 18232 18932 18284
rect 19156 18232 19208 18284
rect 20720 18368 20772 18420
rect 22744 18368 22796 18420
rect 23664 18368 23716 18420
rect 26332 18368 26384 18420
rect 29184 18411 29236 18420
rect 29184 18377 29193 18411
rect 29193 18377 29227 18411
rect 29227 18377 29236 18411
rect 29184 18368 29236 18377
rect 32036 18368 32088 18420
rect 32588 18411 32640 18420
rect 32588 18377 32597 18411
rect 32597 18377 32631 18411
rect 32631 18377 32640 18411
rect 32588 18368 32640 18377
rect 33876 18368 33928 18420
rect 37924 18411 37976 18420
rect 37924 18377 37933 18411
rect 37933 18377 37967 18411
rect 37967 18377 37976 18411
rect 37924 18368 37976 18377
rect 38016 18411 38068 18420
rect 38016 18377 38025 18411
rect 38025 18377 38059 18411
rect 38059 18377 38068 18411
rect 38016 18368 38068 18377
rect 38844 18411 38896 18420
rect 23388 18232 23440 18284
rect 24952 18275 25004 18284
rect 24952 18241 24961 18275
rect 24961 18241 24995 18275
rect 24995 18241 25004 18275
rect 24952 18232 25004 18241
rect 8116 18207 8168 18216
rect 8116 18173 8125 18207
rect 8125 18173 8159 18207
rect 8159 18173 8168 18207
rect 8116 18164 8168 18173
rect 12900 18164 12952 18216
rect 15936 18207 15988 18216
rect 15936 18173 15945 18207
rect 15945 18173 15979 18207
rect 15979 18173 15988 18207
rect 15936 18164 15988 18173
rect 12532 18096 12584 18148
rect 13544 18139 13596 18148
rect 13544 18105 13553 18139
rect 13553 18105 13587 18139
rect 13587 18105 13596 18139
rect 13544 18096 13596 18105
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 12900 18071 12952 18080
rect 12900 18037 12909 18071
rect 12909 18037 12943 18071
rect 12943 18037 12952 18071
rect 12900 18028 12952 18037
rect 15384 18028 15436 18080
rect 15752 18096 15804 18148
rect 20812 18164 20864 18216
rect 25044 18207 25096 18216
rect 20904 18096 20956 18148
rect 23112 18096 23164 18148
rect 23480 18096 23532 18148
rect 25044 18173 25053 18207
rect 25053 18173 25087 18207
rect 25087 18173 25096 18207
rect 25044 18164 25096 18173
rect 26240 18232 26292 18284
rect 27160 18232 27212 18284
rect 31668 18232 31720 18284
rect 32496 18275 32548 18284
rect 32496 18241 32505 18275
rect 32505 18241 32539 18275
rect 32539 18241 32548 18275
rect 32496 18232 32548 18241
rect 34520 18275 34572 18284
rect 26976 18207 27028 18216
rect 18972 18028 19024 18080
rect 20996 18028 21048 18080
rect 24032 18028 24084 18080
rect 26976 18173 26985 18207
rect 26985 18173 27019 18207
rect 27019 18173 27028 18207
rect 26976 18164 27028 18173
rect 32680 18207 32732 18216
rect 26332 18096 26384 18148
rect 27528 18096 27580 18148
rect 32680 18173 32689 18207
rect 32689 18173 32723 18207
rect 32723 18173 32732 18207
rect 32680 18164 32732 18173
rect 33508 18164 33560 18216
rect 34520 18241 34529 18275
rect 34529 18241 34563 18275
rect 34563 18241 34572 18275
rect 34520 18232 34572 18241
rect 34704 18164 34756 18216
rect 37832 18207 37884 18216
rect 37832 18173 37841 18207
rect 37841 18173 37875 18207
rect 37875 18173 37884 18207
rect 37832 18164 37884 18173
rect 38844 18377 38853 18411
rect 38853 18377 38887 18411
rect 38887 18377 38896 18411
rect 38844 18368 38896 18377
rect 41604 18164 41656 18216
rect 25872 18071 25924 18080
rect 25872 18037 25881 18071
rect 25881 18037 25915 18071
rect 25915 18037 25924 18071
rect 25872 18028 25924 18037
rect 39672 18096 39724 18148
rect 32588 18028 32640 18080
rect 34704 18071 34756 18080
rect 34704 18037 34713 18071
rect 34713 18037 34747 18071
rect 34747 18037 34756 18071
rect 34704 18028 34756 18037
rect 43536 18071 43588 18080
rect 43536 18037 43545 18071
rect 43545 18037 43579 18071
rect 43579 18037 43588 18071
rect 43536 18028 43588 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 65654 17926 65706 17978
rect 65718 17926 65770 17978
rect 65782 17926 65834 17978
rect 65846 17926 65898 17978
rect 65910 17926 65962 17978
rect 11796 17824 11848 17876
rect 16396 17867 16448 17876
rect 16396 17833 16405 17867
rect 16405 17833 16439 17867
rect 16439 17833 16448 17867
rect 16396 17824 16448 17833
rect 16948 17824 17000 17876
rect 20444 17824 20496 17876
rect 30288 17824 30340 17876
rect 33508 17867 33560 17876
rect 6460 17756 6512 17808
rect 5448 17731 5500 17740
rect 5448 17697 5457 17731
rect 5457 17697 5491 17731
rect 5491 17697 5500 17731
rect 5448 17688 5500 17697
rect 7380 17688 7432 17740
rect 7656 17731 7708 17740
rect 7656 17697 7665 17731
rect 7665 17697 7699 17731
rect 7699 17697 7708 17731
rect 7656 17688 7708 17697
rect 8116 17688 8168 17740
rect 10968 17688 11020 17740
rect 5724 17620 5776 17672
rect 10416 17620 10468 17672
rect 8116 17552 8168 17604
rect 12900 17620 12952 17672
rect 12532 17552 12584 17604
rect 17408 17756 17460 17808
rect 21088 17756 21140 17808
rect 23020 17799 23072 17808
rect 23020 17765 23029 17799
rect 23029 17765 23063 17799
rect 23063 17765 23072 17799
rect 23020 17756 23072 17765
rect 27252 17756 27304 17808
rect 15752 17620 15804 17672
rect 17868 17620 17920 17672
rect 20260 17688 20312 17740
rect 20628 17663 20680 17672
rect 20628 17629 20637 17663
rect 20637 17629 20671 17663
rect 20671 17629 20680 17663
rect 20628 17620 20680 17629
rect 20812 17663 20864 17672
rect 20812 17629 20821 17663
rect 20821 17629 20855 17663
rect 20855 17629 20864 17663
rect 20812 17620 20864 17629
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 23664 17663 23716 17672
rect 23664 17629 23673 17663
rect 23673 17629 23707 17663
rect 23707 17629 23716 17663
rect 23664 17620 23716 17629
rect 25872 17688 25924 17740
rect 25136 17620 25188 17672
rect 25688 17620 25740 17672
rect 6920 17484 6972 17536
rect 7012 17484 7064 17536
rect 10784 17484 10836 17536
rect 11796 17484 11848 17536
rect 12348 17484 12400 17536
rect 15108 17552 15160 17604
rect 15292 17595 15344 17604
rect 15292 17561 15326 17595
rect 15326 17561 15344 17595
rect 15292 17552 15344 17561
rect 16488 17552 16540 17604
rect 13360 17484 13412 17536
rect 14188 17527 14240 17536
rect 14188 17493 14197 17527
rect 14197 17493 14231 17527
rect 14231 17493 14240 17527
rect 14188 17484 14240 17493
rect 17316 17484 17368 17536
rect 18604 17484 18656 17536
rect 22560 17552 22612 17604
rect 26240 17552 26292 17604
rect 27160 17595 27212 17604
rect 27160 17561 27169 17595
rect 27169 17561 27203 17595
rect 27203 17561 27212 17595
rect 27160 17552 27212 17561
rect 21180 17484 21232 17536
rect 23388 17484 23440 17536
rect 33508 17833 33517 17867
rect 33517 17833 33551 17867
rect 33551 17833 33560 17867
rect 33508 17824 33560 17833
rect 37832 17824 37884 17876
rect 31668 17688 31720 17740
rect 35072 17688 35124 17740
rect 43812 17688 43864 17740
rect 30748 17552 30800 17604
rect 32036 17620 32088 17672
rect 34704 17620 34756 17672
rect 36084 17663 36136 17672
rect 36084 17629 36093 17663
rect 36093 17629 36127 17663
rect 36127 17629 36136 17663
rect 36084 17620 36136 17629
rect 38660 17620 38712 17672
rect 39304 17620 39356 17672
rect 40132 17620 40184 17672
rect 43076 17663 43128 17672
rect 43076 17629 43085 17663
rect 43085 17629 43119 17663
rect 43119 17629 43128 17663
rect 43076 17620 43128 17629
rect 54668 17620 54720 17672
rect 31760 17552 31812 17604
rect 32220 17552 32272 17604
rect 32496 17552 32548 17604
rect 33784 17552 33836 17604
rect 31024 17484 31076 17536
rect 31944 17527 31996 17536
rect 31944 17493 31953 17527
rect 31953 17493 31987 17527
rect 31987 17493 31996 17527
rect 31944 17484 31996 17493
rect 34796 17484 34848 17536
rect 36452 17552 36504 17604
rect 37464 17552 37516 17604
rect 43536 17552 43588 17604
rect 38936 17527 38988 17536
rect 38936 17493 38945 17527
rect 38945 17493 38979 17527
rect 38979 17493 38988 17527
rect 38936 17484 38988 17493
rect 39856 17527 39908 17536
rect 39856 17493 39865 17527
rect 39865 17493 39899 17527
rect 39899 17493 39908 17527
rect 39856 17484 39908 17493
rect 41604 17484 41656 17536
rect 41972 17484 42024 17536
rect 42708 17484 42760 17536
rect 43260 17527 43312 17536
rect 43260 17493 43269 17527
rect 43269 17493 43303 17527
rect 43303 17493 43312 17527
rect 43260 17484 43312 17493
rect 43720 17527 43772 17536
rect 43720 17493 43729 17527
rect 43729 17493 43763 17527
rect 43763 17493 43772 17527
rect 43720 17484 43772 17493
rect 45560 17484 45612 17536
rect 67824 17552 67876 17604
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 6460 17323 6512 17332
rect 6460 17289 6469 17323
rect 6469 17289 6503 17323
rect 6503 17289 6512 17323
rect 6460 17280 6512 17289
rect 7656 17323 7708 17332
rect 7656 17289 7665 17323
rect 7665 17289 7699 17323
rect 7699 17289 7708 17323
rect 7656 17280 7708 17289
rect 15292 17280 15344 17332
rect 19432 17280 19484 17332
rect 20812 17280 20864 17332
rect 22560 17323 22612 17332
rect 22560 17289 22569 17323
rect 22569 17289 22603 17323
rect 22603 17289 22612 17323
rect 22560 17280 22612 17289
rect 27712 17280 27764 17332
rect 5724 17144 5776 17196
rect 7564 17212 7616 17264
rect 11060 17212 11112 17264
rect 10784 17187 10836 17196
rect 10784 17153 10793 17187
rect 10793 17153 10827 17187
rect 10827 17153 10836 17187
rect 10784 17144 10836 17153
rect 12624 17212 12676 17264
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 12716 17187 12768 17196
rect 12716 17153 12725 17187
rect 12725 17153 12759 17187
rect 12759 17153 12768 17187
rect 12716 17144 12768 17153
rect 7104 17076 7156 17128
rect 7472 17076 7524 17128
rect 10416 17076 10468 17128
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 12348 17076 12400 17128
rect 16580 17212 16632 17264
rect 15384 17187 15436 17196
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 17684 17119 17736 17128
rect 17684 17085 17693 17119
rect 17693 17085 17727 17119
rect 17727 17085 17736 17119
rect 17684 17076 17736 17085
rect 10784 17008 10836 17060
rect 12624 17008 12676 17060
rect 19984 17212 20036 17264
rect 18972 17187 19024 17196
rect 17868 17008 17920 17060
rect 4712 16940 4764 16992
rect 10508 16983 10560 16992
rect 10508 16949 10517 16983
rect 10517 16949 10551 16983
rect 10551 16949 10560 16983
rect 10508 16940 10560 16949
rect 11796 16940 11848 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 18236 16940 18288 16992
rect 18972 17153 18981 17187
rect 18981 17153 19015 17187
rect 19015 17153 19024 17187
rect 18972 17144 19024 17153
rect 19156 17144 19208 17196
rect 19432 17144 19484 17196
rect 20076 17144 20128 17196
rect 20168 17187 20220 17196
rect 20168 17153 20177 17187
rect 20177 17153 20211 17187
rect 20211 17153 20220 17187
rect 20168 17144 20220 17153
rect 20628 17144 20680 17196
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 22284 17144 22336 17196
rect 24492 17212 24544 17264
rect 23112 17187 23164 17196
rect 23112 17153 23121 17187
rect 23121 17153 23155 17187
rect 23155 17153 23164 17187
rect 23112 17144 23164 17153
rect 23388 17144 23440 17196
rect 25044 17144 25096 17196
rect 26976 17187 27028 17196
rect 23756 17076 23808 17128
rect 24584 17119 24636 17128
rect 24584 17085 24593 17119
rect 24593 17085 24627 17119
rect 24627 17085 24636 17119
rect 24584 17076 24636 17085
rect 26424 17119 26476 17128
rect 26424 17085 26433 17119
rect 26433 17085 26467 17119
rect 26467 17085 26476 17119
rect 26424 17076 26476 17085
rect 26976 17153 26985 17187
rect 26985 17153 27019 17187
rect 27019 17153 27028 17187
rect 26976 17144 27028 17153
rect 27988 17280 28040 17332
rect 32588 17255 32640 17264
rect 32588 17221 32597 17255
rect 32597 17221 32631 17255
rect 32631 17221 32640 17255
rect 32588 17212 32640 17221
rect 34520 17280 34572 17332
rect 35072 17280 35124 17332
rect 37188 17280 37240 17332
rect 37464 17323 37516 17332
rect 37464 17289 37473 17323
rect 37473 17289 37507 17323
rect 37507 17289 37516 17323
rect 37464 17280 37516 17289
rect 35348 17212 35400 17264
rect 28080 17187 28132 17196
rect 28080 17153 28089 17187
rect 28089 17153 28123 17187
rect 28123 17153 28132 17187
rect 28080 17144 28132 17153
rect 31944 17144 31996 17196
rect 23480 17051 23532 17060
rect 23480 17017 23489 17051
rect 23489 17017 23523 17051
rect 23523 17017 23532 17051
rect 23480 17008 23532 17017
rect 25412 17008 25464 17060
rect 31024 17076 31076 17128
rect 32496 17076 32548 17128
rect 30748 17051 30800 17060
rect 22928 16940 22980 16992
rect 23296 16940 23348 16992
rect 24032 16983 24084 16992
rect 24032 16949 24041 16983
rect 24041 16949 24075 16983
rect 24075 16949 24084 16983
rect 30748 17017 30757 17051
rect 30757 17017 30791 17051
rect 30791 17017 30800 17051
rect 30748 17008 30800 17017
rect 24032 16940 24084 16949
rect 32404 17008 32456 17060
rect 31208 16940 31260 16992
rect 32680 16983 32732 16992
rect 32680 16949 32689 16983
rect 32689 16949 32723 16983
rect 32723 16949 32732 16983
rect 34796 17076 34848 17128
rect 37280 17187 37332 17196
rect 37280 17153 37289 17187
rect 37289 17153 37323 17187
rect 37323 17153 37332 17187
rect 37280 17144 37332 17153
rect 42616 17280 42668 17332
rect 38660 17212 38712 17264
rect 38936 17212 38988 17264
rect 39856 17144 39908 17196
rect 41604 17187 41656 17196
rect 41604 17153 41613 17187
rect 41613 17153 41647 17187
rect 41647 17153 41656 17187
rect 41604 17144 41656 17153
rect 43260 17212 43312 17264
rect 44732 17212 44784 17264
rect 43352 17144 43404 17196
rect 41788 17076 41840 17128
rect 42156 17008 42208 17060
rect 55312 17212 55364 17264
rect 46020 17051 46072 17060
rect 46020 17017 46029 17051
rect 46029 17017 46063 17051
rect 46063 17017 46072 17051
rect 46020 17008 46072 17017
rect 36452 16983 36504 16992
rect 32680 16940 32732 16949
rect 36452 16949 36461 16983
rect 36461 16949 36495 16983
rect 36495 16949 36504 16983
rect 36452 16940 36504 16949
rect 40040 16940 40092 16992
rect 41880 16940 41932 16992
rect 44916 16940 44968 16992
rect 45008 16983 45060 16992
rect 45008 16949 45017 16983
rect 45017 16949 45051 16983
rect 45051 16949 45060 16983
rect 45008 16940 45060 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 65654 16838 65706 16890
rect 65718 16838 65770 16890
rect 65782 16838 65834 16890
rect 65846 16838 65898 16890
rect 65910 16838 65962 16890
rect 4620 16736 4672 16788
rect 5724 16779 5776 16788
rect 5724 16745 5733 16779
rect 5733 16745 5767 16779
rect 5767 16745 5776 16779
rect 5724 16736 5776 16745
rect 11152 16736 11204 16788
rect 12624 16779 12676 16788
rect 12624 16745 12633 16779
rect 12633 16745 12667 16779
rect 12667 16745 12676 16779
rect 12624 16736 12676 16745
rect 16488 16736 16540 16788
rect 9680 16668 9732 16720
rect 10968 16668 11020 16720
rect 12440 16668 12492 16720
rect 4344 16643 4396 16652
rect 4344 16609 4353 16643
rect 4353 16609 4387 16643
rect 4387 16609 4396 16643
rect 4344 16600 4396 16609
rect 6920 16643 6972 16652
rect 6920 16609 6929 16643
rect 6929 16609 6963 16643
rect 6963 16609 6972 16643
rect 6920 16600 6972 16609
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 9036 16643 9088 16652
rect 9036 16609 9045 16643
rect 9045 16609 9079 16643
rect 9079 16609 9088 16643
rect 9036 16600 9088 16609
rect 7012 16575 7064 16584
rect 7012 16541 7021 16575
rect 7021 16541 7055 16575
rect 7055 16541 7064 16575
rect 7012 16532 7064 16541
rect 7656 16532 7708 16584
rect 9220 16575 9272 16584
rect 9220 16541 9229 16575
rect 9229 16541 9263 16575
rect 9263 16541 9272 16575
rect 9220 16532 9272 16541
rect 18236 16736 18288 16788
rect 18880 16736 18932 16788
rect 23388 16779 23440 16788
rect 23388 16745 23397 16779
rect 23397 16745 23431 16779
rect 23431 16745 23440 16779
rect 23388 16736 23440 16745
rect 26424 16736 26476 16788
rect 17040 16668 17092 16720
rect 17684 16668 17736 16720
rect 19156 16668 19208 16720
rect 4712 16464 4764 16516
rect 9128 16464 9180 16516
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 11428 16532 11480 16584
rect 11796 16575 11848 16584
rect 11796 16541 11805 16575
rect 11805 16541 11839 16575
rect 11839 16541 11848 16575
rect 11796 16532 11848 16541
rect 15752 16532 15804 16584
rect 18144 16532 18196 16584
rect 23112 16668 23164 16720
rect 22192 16643 22244 16652
rect 22192 16609 22201 16643
rect 22201 16609 22235 16643
rect 22235 16609 22244 16643
rect 22192 16600 22244 16609
rect 25136 16643 25188 16652
rect 25136 16609 25145 16643
rect 25145 16609 25179 16643
rect 25179 16609 25188 16643
rect 25136 16600 25188 16609
rect 32404 16736 32456 16788
rect 36452 16736 36504 16788
rect 37280 16779 37332 16788
rect 37280 16745 37289 16779
rect 37289 16745 37323 16779
rect 37323 16745 37332 16779
rect 37280 16736 37332 16745
rect 38568 16736 38620 16788
rect 42432 16779 42484 16788
rect 31760 16668 31812 16720
rect 32680 16600 32732 16652
rect 19984 16532 20036 16584
rect 21640 16532 21692 16584
rect 23572 16575 23624 16584
rect 23572 16541 23581 16575
rect 23581 16541 23615 16575
rect 23615 16541 23624 16575
rect 24860 16575 24912 16584
rect 23572 16532 23624 16541
rect 24860 16541 24869 16575
rect 24869 16541 24903 16575
rect 24903 16541 24912 16575
rect 24860 16532 24912 16541
rect 27712 16532 27764 16584
rect 29460 16532 29512 16584
rect 32312 16575 32364 16584
rect 32312 16541 32321 16575
rect 32321 16541 32355 16575
rect 32355 16541 32364 16575
rect 32312 16532 32364 16541
rect 34520 16668 34572 16720
rect 36084 16643 36136 16652
rect 36084 16609 36093 16643
rect 36093 16609 36127 16643
rect 36127 16609 36136 16643
rect 36084 16600 36136 16609
rect 38936 16668 38988 16720
rect 37832 16600 37884 16652
rect 38568 16643 38620 16652
rect 38568 16609 38577 16643
rect 38577 16609 38611 16643
rect 38611 16609 38620 16643
rect 38568 16600 38620 16609
rect 33784 16575 33836 16584
rect 33784 16541 33793 16575
rect 33793 16541 33827 16575
rect 33827 16541 33836 16575
rect 33784 16532 33836 16541
rect 40316 16600 40368 16652
rect 41512 16668 41564 16720
rect 42432 16745 42441 16779
rect 42441 16745 42475 16779
rect 42475 16745 42484 16779
rect 42432 16736 42484 16745
rect 43076 16736 43128 16788
rect 43812 16736 43864 16788
rect 40040 16575 40092 16584
rect 40040 16541 40049 16575
rect 40049 16541 40083 16575
rect 40083 16541 40092 16575
rect 40040 16532 40092 16541
rect 41052 16575 41104 16584
rect 41052 16541 41061 16575
rect 41061 16541 41095 16575
rect 41095 16541 41104 16575
rect 41052 16532 41104 16541
rect 16672 16464 16724 16516
rect 17868 16464 17920 16516
rect 19340 16464 19392 16516
rect 24584 16464 24636 16516
rect 25044 16464 25096 16516
rect 10600 16396 10652 16448
rect 11428 16396 11480 16448
rect 12164 16396 12216 16448
rect 17040 16396 17092 16448
rect 20076 16396 20128 16448
rect 22836 16396 22888 16448
rect 26148 16439 26200 16448
rect 26148 16405 26157 16439
rect 26157 16405 26191 16439
rect 26191 16405 26200 16439
rect 26148 16396 26200 16405
rect 33968 16464 34020 16516
rect 29920 16396 29972 16448
rect 32496 16439 32548 16448
rect 32496 16405 32505 16439
rect 32505 16405 32539 16439
rect 32539 16405 32548 16439
rect 32496 16396 32548 16405
rect 34152 16439 34204 16448
rect 34152 16405 34161 16439
rect 34161 16405 34195 16439
rect 34195 16405 34204 16439
rect 34152 16396 34204 16405
rect 34428 16396 34480 16448
rect 38108 16396 38160 16448
rect 38844 16439 38896 16448
rect 38844 16405 38853 16439
rect 38853 16405 38887 16439
rect 38887 16405 38896 16439
rect 38844 16396 38896 16405
rect 40132 16396 40184 16448
rect 40408 16396 40460 16448
rect 42156 16575 42208 16584
rect 42156 16541 42165 16575
rect 42165 16541 42199 16575
rect 42199 16541 42208 16575
rect 43812 16643 43864 16652
rect 43812 16609 43821 16643
rect 43821 16609 43855 16643
rect 43855 16609 43864 16643
rect 43812 16600 43864 16609
rect 45008 16600 45060 16652
rect 45192 16711 45244 16720
rect 45192 16677 45201 16711
rect 45201 16677 45235 16711
rect 45235 16677 45244 16711
rect 45192 16668 45244 16677
rect 45560 16643 45612 16652
rect 45560 16609 45569 16643
rect 45569 16609 45603 16643
rect 45603 16609 45612 16643
rect 45560 16600 45612 16609
rect 45376 16575 45428 16584
rect 42156 16532 42208 16541
rect 45376 16541 45385 16575
rect 45385 16541 45419 16575
rect 45419 16541 45428 16575
rect 45376 16532 45428 16541
rect 46020 16575 46072 16584
rect 46020 16541 46029 16575
rect 46029 16541 46063 16575
rect 46063 16541 46072 16575
rect 46020 16532 46072 16541
rect 42616 16464 42668 16516
rect 44916 16464 44968 16516
rect 43260 16396 43312 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 7472 16192 7524 16244
rect 9036 16192 9088 16244
rect 11152 16192 11204 16244
rect 15108 16192 15160 16244
rect 11520 16124 11572 16176
rect 11980 16167 12032 16176
rect 11980 16133 11989 16167
rect 11989 16133 12023 16167
rect 12023 16133 12032 16167
rect 11980 16124 12032 16133
rect 12808 16167 12860 16176
rect 12808 16133 12817 16167
rect 12817 16133 12851 16167
rect 12851 16133 12860 16167
rect 18236 16192 18288 16244
rect 20444 16192 20496 16244
rect 23572 16192 23624 16244
rect 25412 16192 25464 16244
rect 26148 16192 26200 16244
rect 27712 16235 27764 16244
rect 12808 16124 12860 16133
rect 22836 16124 22888 16176
rect 27712 16201 27721 16235
rect 27721 16201 27755 16235
rect 27755 16201 27764 16235
rect 27712 16192 27764 16201
rect 29460 16235 29512 16244
rect 29460 16201 29469 16235
rect 29469 16201 29503 16235
rect 29503 16201 29512 16235
rect 29460 16192 29512 16201
rect 29920 16235 29972 16244
rect 29920 16201 29929 16235
rect 29929 16201 29963 16235
rect 29963 16201 29972 16235
rect 29920 16192 29972 16201
rect 32312 16235 32364 16244
rect 32312 16201 32321 16235
rect 32321 16201 32355 16235
rect 32355 16201 32364 16235
rect 32312 16192 32364 16201
rect 33968 16235 34020 16244
rect 33968 16201 33977 16235
rect 33977 16201 34011 16235
rect 34011 16201 34020 16235
rect 33968 16192 34020 16201
rect 42616 16192 42668 16244
rect 4344 16056 4396 16108
rect 5172 16056 5224 16108
rect 7748 16099 7800 16108
rect 7748 16065 7757 16099
rect 7757 16065 7791 16099
rect 7791 16065 7800 16099
rect 7748 16056 7800 16065
rect 10600 16099 10652 16108
rect 10600 16065 10609 16099
rect 10609 16065 10643 16099
rect 10643 16065 10652 16099
rect 10600 16056 10652 16065
rect 16948 16056 17000 16108
rect 24768 16099 24820 16108
rect 24768 16065 24777 16099
rect 24777 16065 24811 16099
rect 24811 16065 24820 16099
rect 33508 16124 33560 16176
rect 34428 16124 34480 16176
rect 45560 16192 45612 16244
rect 24768 16056 24820 16065
rect 29828 16099 29880 16108
rect 5448 15920 5500 15972
rect 6920 16031 6972 16040
rect 6920 15997 6929 16031
rect 6929 15997 6963 16031
rect 6963 15997 6972 16031
rect 7840 16031 7892 16040
rect 6920 15988 6972 15997
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 10508 16031 10560 16040
rect 10508 15997 10517 16031
rect 10517 15997 10551 16031
rect 10551 15997 10560 16031
rect 10508 15988 10560 15997
rect 15936 16031 15988 16040
rect 15936 15997 15945 16031
rect 15945 15997 15979 16031
rect 15979 15997 15988 16031
rect 15936 15988 15988 15997
rect 18144 16031 18196 16040
rect 18144 15997 18153 16031
rect 18153 15997 18187 16031
rect 18187 15997 18196 16031
rect 18144 15988 18196 15997
rect 22652 15988 22704 16040
rect 27068 16031 27120 16040
rect 27068 15997 27077 16031
rect 27077 15997 27111 16031
rect 27111 15997 27120 16031
rect 27068 15988 27120 15997
rect 29828 16065 29837 16099
rect 29837 16065 29871 16099
rect 29871 16065 29880 16099
rect 29828 16056 29880 16065
rect 34152 16056 34204 16108
rect 34796 16099 34848 16108
rect 34796 16065 34805 16099
rect 34805 16065 34839 16099
rect 34839 16065 34848 16099
rect 34796 16056 34848 16065
rect 43720 16056 43772 16108
rect 32772 16031 32824 16040
rect 12164 15920 12216 15972
rect 24676 15920 24728 15972
rect 28080 15920 28132 15972
rect 32772 15997 32781 16031
rect 32781 15997 32815 16031
rect 32815 15997 32824 16031
rect 32772 15988 32824 15997
rect 32680 15920 32732 15972
rect 34612 15988 34664 16040
rect 42432 15988 42484 16040
rect 8576 15895 8628 15904
rect 8576 15861 8585 15895
rect 8585 15861 8619 15895
rect 8619 15861 8628 15895
rect 8576 15852 8628 15861
rect 14096 15852 14148 15904
rect 15292 15895 15344 15904
rect 15292 15861 15301 15895
rect 15301 15861 15335 15895
rect 15335 15861 15344 15895
rect 15292 15852 15344 15861
rect 28264 15895 28316 15904
rect 28264 15861 28273 15895
rect 28273 15861 28307 15895
rect 28307 15861 28316 15895
rect 28264 15852 28316 15861
rect 28908 15895 28960 15904
rect 28908 15861 28917 15895
rect 28917 15861 28951 15895
rect 28951 15861 28960 15895
rect 28908 15852 28960 15861
rect 34428 15895 34480 15904
rect 34428 15861 34437 15895
rect 34437 15861 34471 15895
rect 34471 15861 34480 15895
rect 34428 15852 34480 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 65654 15750 65706 15802
rect 65718 15750 65770 15802
rect 65782 15750 65834 15802
rect 65846 15750 65898 15802
rect 65910 15750 65962 15802
rect 5172 15691 5224 15700
rect 5172 15657 5181 15691
rect 5181 15657 5215 15691
rect 5215 15657 5224 15691
rect 5172 15648 5224 15657
rect 6460 15648 6512 15700
rect 7012 15648 7064 15700
rect 7748 15648 7800 15700
rect 6828 15580 6880 15632
rect 4620 15512 4672 15564
rect 5448 15444 5500 15496
rect 7104 15512 7156 15564
rect 15752 15648 15804 15700
rect 16856 15648 16908 15700
rect 22192 15648 22244 15700
rect 16764 15580 16816 15632
rect 24032 15648 24084 15700
rect 28080 15648 28132 15700
rect 28264 15648 28316 15700
rect 28908 15648 28960 15700
rect 38384 15648 38436 15700
rect 40040 15648 40092 15700
rect 41328 15648 41380 15700
rect 23572 15580 23624 15632
rect 17224 15555 17276 15564
rect 8300 15444 8352 15496
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 6368 15376 6420 15428
rect 9680 15419 9732 15428
rect 9680 15385 9689 15419
rect 9689 15385 9723 15419
rect 9723 15385 9732 15419
rect 17224 15521 17233 15555
rect 17233 15521 17267 15555
rect 17267 15521 17276 15555
rect 17224 15512 17276 15521
rect 26148 15512 26200 15564
rect 40316 15580 40368 15632
rect 41788 15623 41840 15632
rect 41788 15589 41797 15623
rect 41797 15589 41831 15623
rect 41831 15589 41840 15623
rect 41788 15580 41840 15589
rect 42616 15648 42668 15700
rect 45376 15580 45428 15632
rect 28172 15512 28224 15564
rect 41604 15512 41656 15564
rect 11980 15444 12032 15496
rect 15292 15444 15344 15496
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 19340 15444 19392 15496
rect 19984 15444 20036 15496
rect 22284 15487 22336 15496
rect 22284 15453 22293 15487
rect 22293 15453 22327 15487
rect 22327 15453 22336 15487
rect 22284 15444 22336 15453
rect 22468 15487 22520 15496
rect 22468 15453 22477 15487
rect 22477 15453 22511 15487
rect 22511 15453 22520 15487
rect 22468 15444 22520 15453
rect 23756 15444 23808 15496
rect 12532 15419 12584 15428
rect 9680 15376 9732 15385
rect 8208 15308 8260 15360
rect 10140 15308 10192 15360
rect 11060 15308 11112 15360
rect 11428 15351 11480 15360
rect 11428 15317 11437 15351
rect 11437 15317 11471 15351
rect 11471 15317 11480 15351
rect 11428 15308 11480 15317
rect 12532 15385 12550 15419
rect 12550 15385 12584 15419
rect 12532 15376 12584 15385
rect 13728 15308 13780 15360
rect 16580 15376 16632 15428
rect 23388 15376 23440 15428
rect 24860 15376 24912 15428
rect 16948 15308 17000 15360
rect 19340 15351 19392 15360
rect 19340 15317 19349 15351
rect 19349 15317 19383 15351
rect 19383 15317 19392 15351
rect 19340 15308 19392 15317
rect 20628 15308 20680 15360
rect 22376 15351 22428 15360
rect 22376 15317 22385 15351
rect 22385 15317 22419 15351
rect 22419 15317 22428 15351
rect 22376 15308 22428 15317
rect 22928 15351 22980 15360
rect 22928 15317 22937 15351
rect 22937 15317 22971 15351
rect 22971 15317 22980 15351
rect 22928 15308 22980 15317
rect 23664 15308 23716 15360
rect 25688 15308 25740 15360
rect 29368 15444 29420 15496
rect 29920 15487 29972 15496
rect 29920 15453 29929 15487
rect 29929 15453 29963 15487
rect 29963 15453 29972 15487
rect 29920 15444 29972 15453
rect 32864 15444 32916 15496
rect 32496 15376 32548 15428
rect 39672 15376 39724 15428
rect 43168 15444 43220 15496
rect 43260 15487 43312 15496
rect 43260 15453 43269 15487
rect 43269 15453 43303 15487
rect 43303 15453 43312 15487
rect 43260 15444 43312 15453
rect 28172 15308 28224 15360
rect 28540 15351 28592 15360
rect 28540 15317 28549 15351
rect 28549 15317 28583 15351
rect 28583 15317 28592 15351
rect 28540 15308 28592 15317
rect 29552 15351 29604 15360
rect 29552 15317 29561 15351
rect 29561 15317 29595 15351
rect 29595 15317 29604 15351
rect 29552 15308 29604 15317
rect 32772 15308 32824 15360
rect 40408 15308 40460 15360
rect 41512 15308 41564 15360
rect 43536 15308 43588 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 7012 15147 7064 15156
rect 7012 15113 7021 15147
rect 7021 15113 7055 15147
rect 7055 15113 7064 15147
rect 7012 15104 7064 15113
rect 10600 15147 10652 15156
rect 10600 15113 10609 15147
rect 10609 15113 10643 15147
rect 10643 15113 10652 15147
rect 10600 15104 10652 15113
rect 11060 15104 11112 15156
rect 12348 15104 12400 15156
rect 12532 15147 12584 15156
rect 12532 15113 12541 15147
rect 12541 15113 12575 15147
rect 12575 15113 12584 15147
rect 12532 15104 12584 15113
rect 8300 14968 8352 15020
rect 9956 14968 10008 15020
rect 20628 15104 20680 15156
rect 22284 15104 22336 15156
rect 26240 15104 26292 15156
rect 27068 15104 27120 15156
rect 27252 15147 27304 15156
rect 27252 15113 27261 15147
rect 27261 15113 27295 15147
rect 27295 15113 27304 15147
rect 27252 15104 27304 15113
rect 27344 15104 27396 15156
rect 13452 15036 13504 15088
rect 15936 15036 15988 15088
rect 7380 14900 7432 14952
rect 11428 14900 11480 14952
rect 14096 14968 14148 15020
rect 14464 14968 14516 15020
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 17224 15011 17276 15020
rect 17224 14977 17233 15011
rect 17233 14977 17267 15011
rect 17267 14977 17276 15011
rect 17224 14968 17276 14977
rect 14740 14900 14792 14952
rect 18144 14943 18196 14952
rect 18144 14909 18153 14943
rect 18153 14909 18187 14943
rect 18187 14909 18196 14943
rect 21640 15036 21692 15088
rect 22008 15079 22060 15088
rect 22008 15045 22033 15079
rect 22033 15045 22060 15079
rect 22008 15036 22060 15045
rect 22376 15036 22428 15088
rect 23664 15036 23716 15088
rect 18420 15011 18472 15020
rect 18420 14977 18454 15011
rect 18454 14977 18472 15011
rect 18420 14968 18472 14977
rect 19432 14968 19484 15020
rect 20536 14968 20588 15020
rect 21272 14968 21324 15020
rect 24216 14968 24268 15020
rect 27528 15036 27580 15088
rect 32864 15036 32916 15088
rect 34520 15104 34572 15156
rect 38844 15147 38896 15156
rect 38844 15113 38853 15147
rect 38853 15113 38887 15147
rect 38887 15113 38896 15147
rect 38844 15104 38896 15113
rect 39764 15147 39816 15156
rect 39764 15113 39773 15147
rect 39773 15113 39807 15147
rect 39807 15113 39816 15147
rect 39764 15104 39816 15113
rect 26792 14968 26844 15020
rect 28080 15011 28132 15020
rect 28080 14977 28084 15011
rect 28084 14977 28118 15011
rect 28118 14977 28132 15011
rect 28080 14968 28132 14977
rect 18144 14900 18196 14909
rect 26516 14900 26568 14952
rect 28264 15011 28316 15020
rect 28264 14977 28273 15011
rect 28273 14977 28307 15011
rect 28307 14977 28316 15011
rect 28264 14968 28316 14977
rect 6552 14764 6604 14816
rect 12440 14832 12492 14884
rect 28540 15011 28592 15020
rect 28540 14977 28549 15011
rect 28549 14977 28583 15011
rect 28583 14977 28592 15011
rect 29460 15011 29512 15020
rect 28540 14968 28592 14977
rect 29460 14977 29469 15011
rect 29469 14977 29503 15011
rect 29503 14977 29512 15011
rect 29460 14968 29512 14977
rect 30104 14968 30156 15020
rect 32312 14968 32364 15020
rect 29552 14943 29604 14952
rect 29552 14909 29561 14943
rect 29561 14909 29595 14943
rect 29595 14909 29604 14943
rect 29552 14900 29604 14909
rect 30564 14943 30616 14952
rect 30564 14909 30573 14943
rect 30573 14909 30607 14943
rect 30607 14909 30616 14943
rect 30564 14900 30616 14909
rect 31484 14900 31536 14952
rect 31852 14900 31904 14952
rect 33232 15011 33284 15020
rect 33232 14977 33241 15011
rect 33241 14977 33275 15011
rect 33275 14977 33284 15011
rect 34428 15036 34480 15088
rect 40040 15079 40092 15088
rect 40040 15045 40049 15079
rect 40049 15045 40083 15079
rect 40083 15045 40092 15079
rect 40040 15036 40092 15045
rect 40408 15104 40460 15156
rect 41052 15104 41104 15156
rect 33232 14968 33284 14977
rect 37188 14968 37240 15020
rect 37280 14943 37332 14952
rect 37280 14909 37289 14943
rect 37289 14909 37323 14943
rect 37323 14909 37332 14943
rect 37280 14900 37332 14909
rect 39212 14968 39264 15020
rect 41604 15036 41656 15088
rect 43536 15036 43588 15088
rect 40408 15011 40460 15020
rect 40408 14977 40417 15011
rect 40417 14977 40451 15011
rect 40451 14977 40460 15011
rect 40408 14968 40460 14977
rect 41328 15011 41380 15020
rect 41328 14977 41330 15011
rect 41330 14977 41364 15011
rect 41364 14977 41380 15011
rect 38752 14943 38804 14952
rect 38752 14909 38761 14943
rect 38761 14909 38795 14943
rect 38795 14909 38804 14943
rect 38752 14900 38804 14909
rect 41328 14968 41380 14977
rect 41512 15011 41564 15020
rect 41512 14977 41521 15011
rect 41521 14977 41555 15011
rect 41555 14977 41564 15011
rect 41512 14968 41564 14977
rect 43168 14968 43220 15020
rect 43352 15011 43404 15020
rect 43352 14977 43361 15011
rect 43361 14977 43395 15011
rect 43395 14977 43404 15011
rect 43352 14968 43404 14977
rect 44088 15011 44140 15020
rect 44088 14977 44122 15011
rect 44122 14977 44140 15011
rect 44088 14968 44140 14977
rect 42432 14900 42484 14952
rect 8576 14764 8628 14816
rect 12532 14764 12584 14816
rect 19340 14764 19392 14816
rect 19616 14764 19668 14816
rect 21732 14764 21784 14816
rect 24492 14764 24544 14816
rect 27344 14764 27396 14816
rect 31944 14764 31996 14816
rect 36452 14764 36504 14816
rect 41144 14832 41196 14884
rect 39120 14764 39172 14816
rect 45192 14807 45244 14816
rect 45192 14773 45201 14807
rect 45201 14773 45235 14807
rect 45235 14773 45244 14807
rect 45192 14764 45244 14773
rect 45468 14764 45520 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 65654 14662 65706 14714
rect 65718 14662 65770 14714
rect 65782 14662 65834 14714
rect 65846 14662 65898 14714
rect 65910 14662 65962 14714
rect 6368 14603 6420 14612
rect 6368 14569 6377 14603
rect 6377 14569 6411 14603
rect 6411 14569 6420 14603
rect 6368 14560 6420 14569
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 12532 14560 12584 14612
rect 13452 14603 13504 14612
rect 13452 14569 13461 14603
rect 13461 14569 13495 14603
rect 13495 14569 13504 14603
rect 13452 14560 13504 14569
rect 18420 14560 18472 14612
rect 20536 14603 20588 14612
rect 20536 14569 20545 14603
rect 20545 14569 20579 14603
rect 20579 14569 20588 14603
rect 20536 14560 20588 14569
rect 22468 14560 22520 14612
rect 24216 14560 24268 14612
rect 26792 14560 26844 14612
rect 28356 14560 28408 14612
rect 29460 14560 29512 14612
rect 32312 14603 32364 14612
rect 32312 14569 32321 14603
rect 32321 14569 32355 14603
rect 32355 14569 32364 14603
rect 32312 14560 32364 14569
rect 37280 14603 37332 14612
rect 37280 14569 37289 14603
rect 37289 14569 37323 14603
rect 37323 14569 37332 14603
rect 37280 14560 37332 14569
rect 39212 14603 39264 14612
rect 39212 14569 39221 14603
rect 39221 14569 39255 14603
rect 39255 14569 39264 14603
rect 39212 14560 39264 14569
rect 40316 14603 40368 14612
rect 40316 14569 40325 14603
rect 40325 14569 40359 14603
rect 40359 14569 40368 14603
rect 40316 14560 40368 14569
rect 40408 14560 40460 14612
rect 17224 14492 17276 14544
rect 18328 14492 18380 14544
rect 24676 14492 24728 14544
rect 15752 14467 15804 14476
rect 15752 14433 15761 14467
rect 15761 14433 15795 14467
rect 15795 14433 15804 14467
rect 15752 14424 15804 14433
rect 19432 14424 19484 14476
rect 20536 14424 20588 14476
rect 6552 14399 6604 14408
rect 6552 14365 6561 14399
rect 6561 14365 6595 14399
rect 6595 14365 6604 14399
rect 6552 14356 6604 14365
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 8208 14356 8260 14365
rect 10140 14399 10192 14408
rect 10140 14365 10149 14399
rect 10149 14365 10183 14399
rect 10183 14365 10192 14399
rect 10140 14356 10192 14365
rect 14372 14356 14424 14408
rect 16764 14356 16816 14408
rect 16120 14288 16172 14340
rect 16948 14356 17000 14408
rect 18512 14356 18564 14408
rect 19248 14356 19300 14408
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 24768 14424 24820 14476
rect 28172 14492 28224 14544
rect 35532 14492 35584 14544
rect 48688 14492 48740 14544
rect 56324 14492 56376 14544
rect 30104 14424 30156 14476
rect 31944 14467 31996 14476
rect 31944 14433 31953 14467
rect 31953 14433 31987 14467
rect 31987 14433 31996 14467
rect 31944 14424 31996 14433
rect 37188 14424 37240 14476
rect 7104 14263 7156 14272
rect 7104 14229 7113 14263
rect 7113 14229 7147 14263
rect 7147 14229 7156 14263
rect 7104 14220 7156 14229
rect 7380 14220 7432 14272
rect 15200 14220 15252 14272
rect 19156 14220 19208 14272
rect 19340 14220 19392 14272
rect 20904 14356 20956 14408
rect 19800 14288 19852 14340
rect 22100 14356 22152 14408
rect 23664 14356 23716 14408
rect 29368 14356 29420 14408
rect 30564 14356 30616 14408
rect 32772 14356 32824 14408
rect 33140 14399 33192 14408
rect 33140 14365 33149 14399
rect 33149 14365 33183 14399
rect 33183 14365 33192 14399
rect 33140 14356 33192 14365
rect 38476 14356 38528 14408
rect 21640 14288 21692 14340
rect 23296 14288 23348 14340
rect 20996 14220 21048 14272
rect 21732 14220 21784 14272
rect 26516 14288 26568 14340
rect 36176 14331 36228 14340
rect 36176 14297 36210 14331
rect 36210 14297 36228 14331
rect 36176 14288 36228 14297
rect 37280 14288 37332 14340
rect 38752 14356 38804 14408
rect 39856 14356 39908 14408
rect 40040 14399 40092 14408
rect 40040 14365 40049 14399
rect 40049 14365 40083 14399
rect 40083 14365 40092 14399
rect 40868 14399 40920 14408
rect 40040 14356 40092 14365
rect 40868 14365 40877 14399
rect 40877 14365 40911 14399
rect 40911 14365 40920 14399
rect 40868 14356 40920 14365
rect 41144 14399 41196 14408
rect 41144 14365 41153 14399
rect 41153 14365 41187 14399
rect 41187 14365 41196 14399
rect 41144 14356 41196 14365
rect 42616 14356 42668 14408
rect 45192 14356 45244 14408
rect 45468 14356 45520 14408
rect 43352 14288 43404 14340
rect 26424 14263 26476 14272
rect 26424 14229 26433 14263
rect 26433 14229 26467 14263
rect 26467 14229 26476 14263
rect 26424 14220 26476 14229
rect 27436 14263 27488 14272
rect 27436 14229 27445 14263
rect 27445 14229 27479 14263
rect 27479 14229 27488 14263
rect 27436 14220 27488 14229
rect 29736 14263 29788 14272
rect 29736 14229 29745 14263
rect 29745 14229 29779 14263
rect 29779 14229 29788 14263
rect 29736 14220 29788 14229
rect 33416 14220 33468 14272
rect 37372 14220 37424 14272
rect 38108 14263 38160 14272
rect 38108 14229 38117 14263
rect 38117 14229 38151 14263
rect 38151 14229 38160 14263
rect 38108 14220 38160 14229
rect 41696 14220 41748 14272
rect 43076 14220 43128 14272
rect 43628 14220 43680 14272
rect 44180 14220 44232 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 12072 14016 12124 14068
rect 15200 14016 15252 14068
rect 16764 14059 16816 14068
rect 16764 14025 16773 14059
rect 16773 14025 16807 14059
rect 16807 14025 16816 14059
rect 16764 14016 16816 14025
rect 17500 14016 17552 14068
rect 19340 14016 19392 14068
rect 12532 13948 12584 14000
rect 13820 13991 13872 14000
rect 13820 13957 13829 13991
rect 13829 13957 13863 13991
rect 13863 13957 13872 13991
rect 13820 13948 13872 13957
rect 4896 13880 4948 13932
rect 10784 13923 10836 13932
rect 10784 13889 10793 13923
rect 10793 13889 10827 13923
rect 10827 13889 10836 13923
rect 10784 13880 10836 13889
rect 16396 13948 16448 14000
rect 17224 13948 17276 14000
rect 14372 13880 14424 13932
rect 14924 13923 14976 13932
rect 6736 13855 6788 13864
rect 6736 13821 6745 13855
rect 6745 13821 6779 13855
rect 6779 13821 6788 13855
rect 6736 13812 6788 13821
rect 10876 13812 10928 13864
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 19156 13880 19208 13932
rect 20720 14016 20772 14068
rect 23296 14059 23348 14068
rect 23296 14025 23305 14059
rect 23305 14025 23339 14059
rect 23339 14025 23348 14059
rect 23296 14016 23348 14025
rect 23664 14059 23716 14068
rect 23664 14025 23673 14059
rect 23673 14025 23707 14059
rect 23707 14025 23716 14059
rect 23664 14016 23716 14025
rect 19892 13880 19944 13932
rect 20996 13923 21048 13932
rect 20996 13889 21005 13923
rect 21005 13889 21039 13923
rect 21039 13889 21048 13923
rect 20996 13880 21048 13889
rect 21640 13948 21692 14000
rect 26424 14016 26476 14068
rect 35992 14016 36044 14068
rect 36176 14059 36228 14068
rect 36176 14025 36185 14059
rect 36185 14025 36219 14059
rect 36219 14025 36228 14059
rect 36176 14016 36228 14025
rect 39856 14059 39908 14068
rect 39856 14025 39865 14059
rect 39865 14025 39899 14059
rect 39899 14025 39908 14059
rect 39856 14016 39908 14025
rect 35624 13948 35676 14000
rect 22008 13923 22060 13932
rect 22008 13889 22017 13923
rect 22017 13889 22051 13923
rect 22051 13889 22060 13923
rect 22008 13880 22060 13889
rect 14740 13855 14792 13864
rect 7104 13787 7156 13796
rect 7104 13753 7113 13787
rect 7113 13753 7147 13787
rect 7147 13753 7156 13787
rect 7104 13744 7156 13753
rect 7748 13744 7800 13796
rect 10600 13744 10652 13796
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 15476 13812 15528 13864
rect 12624 13744 12676 13796
rect 16488 13744 16540 13796
rect 20536 13812 20588 13864
rect 20812 13812 20864 13864
rect 23388 13880 23440 13932
rect 25320 13880 25372 13932
rect 26516 13880 26568 13932
rect 33416 13923 33468 13932
rect 33416 13889 33450 13923
rect 33450 13889 33468 13923
rect 33416 13880 33468 13889
rect 37372 13880 37424 13932
rect 25688 13855 25740 13864
rect 25688 13821 25697 13855
rect 25697 13821 25731 13855
rect 25731 13821 25740 13855
rect 25688 13812 25740 13821
rect 26332 13812 26384 13864
rect 27436 13855 27488 13864
rect 27436 13821 27445 13855
rect 27445 13821 27479 13855
rect 27479 13821 27488 13855
rect 27436 13812 27488 13821
rect 27068 13744 27120 13796
rect 32864 13812 32916 13864
rect 37280 13812 37332 13864
rect 39672 13948 39724 14000
rect 43168 14016 43220 14068
rect 45192 13948 45244 14000
rect 38476 13923 38528 13932
rect 38476 13889 38485 13923
rect 38485 13889 38519 13923
rect 38519 13889 38528 13923
rect 38476 13880 38528 13889
rect 38752 13923 38804 13932
rect 38752 13889 38786 13923
rect 38786 13889 38804 13923
rect 41696 13923 41748 13932
rect 38752 13880 38804 13889
rect 41696 13889 41705 13923
rect 41705 13889 41739 13923
rect 41739 13889 41748 13923
rect 41696 13880 41748 13889
rect 39856 13812 39908 13864
rect 40868 13812 40920 13864
rect 41604 13812 41656 13864
rect 42432 13855 42484 13864
rect 42432 13821 42441 13855
rect 42441 13821 42475 13855
rect 42475 13821 42484 13855
rect 42432 13812 42484 13821
rect 29828 13744 29880 13796
rect 32496 13744 32548 13796
rect 32588 13744 32640 13796
rect 33048 13744 33100 13796
rect 44364 13787 44416 13796
rect 44364 13753 44373 13787
rect 44373 13753 44407 13787
rect 44407 13753 44416 13787
rect 44364 13744 44416 13753
rect 45468 13744 45520 13796
rect 4988 13676 5040 13728
rect 7656 13719 7708 13728
rect 7656 13685 7665 13719
rect 7665 13685 7699 13719
rect 7699 13685 7708 13719
rect 7656 13676 7708 13685
rect 9772 13676 9824 13728
rect 11704 13676 11756 13728
rect 19340 13719 19392 13728
rect 19340 13685 19349 13719
rect 19349 13685 19383 13719
rect 19383 13685 19392 13719
rect 19340 13676 19392 13685
rect 19892 13676 19944 13728
rect 21088 13676 21140 13728
rect 21824 13719 21876 13728
rect 21824 13685 21833 13719
rect 21833 13685 21867 13719
rect 21867 13685 21876 13719
rect 21824 13676 21876 13685
rect 34520 13719 34572 13728
rect 34520 13685 34529 13719
rect 34529 13685 34563 13719
rect 34563 13685 34572 13719
rect 34520 13676 34572 13685
rect 43076 13676 43128 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 65654 13574 65706 13626
rect 65718 13574 65770 13626
rect 65782 13574 65834 13626
rect 65846 13574 65898 13626
rect 65910 13574 65962 13626
rect 7656 13472 7708 13524
rect 12072 13472 12124 13524
rect 14740 13472 14792 13524
rect 16120 13472 16172 13524
rect 16396 13472 16448 13524
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 19156 13472 19208 13524
rect 4712 13311 4764 13320
rect 4712 13277 4721 13311
rect 4721 13277 4755 13311
rect 4755 13277 4764 13311
rect 4712 13268 4764 13277
rect 4988 13311 5040 13320
rect 4988 13277 5022 13311
rect 5022 13277 5040 13311
rect 4988 13268 5040 13277
rect 6736 13268 6788 13320
rect 7748 13311 7800 13320
rect 7748 13277 7757 13311
rect 7757 13277 7791 13311
rect 7791 13277 7800 13311
rect 7748 13268 7800 13277
rect 11520 13268 11572 13320
rect 14556 13268 14608 13320
rect 16212 13336 16264 13388
rect 20904 13472 20956 13524
rect 30104 13515 30156 13524
rect 23388 13447 23440 13456
rect 23388 13413 23397 13447
rect 23397 13413 23431 13447
rect 23431 13413 23440 13447
rect 23388 13404 23440 13413
rect 26424 13404 26476 13456
rect 30104 13481 30113 13515
rect 30113 13481 30147 13515
rect 30147 13481 30156 13515
rect 30104 13472 30156 13481
rect 33140 13472 33192 13524
rect 35992 13472 36044 13524
rect 17868 13336 17920 13388
rect 27528 13379 27580 13388
rect 27528 13345 27537 13379
rect 27537 13345 27571 13379
rect 27571 13345 27580 13379
rect 27528 13336 27580 13345
rect 28080 13336 28132 13388
rect 15752 13268 15804 13320
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 21824 13311 21876 13320
rect 21824 13277 21858 13311
rect 21858 13277 21876 13311
rect 21824 13268 21876 13277
rect 27712 13268 27764 13320
rect 33232 13404 33284 13456
rect 32588 13336 32640 13388
rect 33876 13336 33928 13388
rect 8392 13200 8444 13252
rect 11428 13200 11480 13252
rect 12808 13200 12860 13252
rect 14096 13200 14148 13252
rect 6092 13175 6144 13184
rect 6092 13141 6101 13175
rect 6101 13141 6135 13175
rect 6135 13141 6144 13175
rect 6092 13132 6144 13141
rect 7840 13132 7892 13184
rect 19432 13200 19484 13252
rect 20904 13200 20956 13252
rect 24952 13200 25004 13252
rect 31944 13268 31996 13320
rect 33416 13311 33468 13320
rect 33416 13277 33425 13311
rect 33425 13277 33459 13311
rect 33459 13277 33468 13311
rect 33416 13268 33468 13277
rect 34520 13268 34572 13320
rect 38108 13472 38160 13524
rect 38384 13515 38436 13524
rect 38384 13481 38393 13515
rect 38393 13481 38427 13515
rect 38427 13481 38436 13515
rect 38384 13472 38436 13481
rect 38752 13472 38804 13524
rect 42248 13472 42300 13524
rect 43352 13515 43404 13524
rect 43352 13481 43361 13515
rect 43361 13481 43395 13515
rect 43395 13481 43404 13515
rect 43352 13472 43404 13481
rect 43536 13515 43588 13524
rect 43536 13481 43545 13515
rect 43545 13481 43579 13515
rect 43579 13481 43588 13515
rect 43536 13472 43588 13481
rect 44088 13472 44140 13524
rect 39856 13379 39908 13388
rect 39856 13345 39865 13379
rect 39865 13345 39899 13379
rect 39899 13345 39908 13379
rect 39856 13336 39908 13345
rect 39120 13311 39172 13320
rect 39120 13277 39129 13311
rect 39129 13277 39163 13311
rect 39163 13277 39172 13311
rect 39120 13268 39172 13277
rect 22468 13132 22520 13184
rect 26148 13175 26200 13184
rect 26148 13141 26157 13175
rect 26157 13141 26191 13175
rect 26191 13141 26200 13175
rect 26148 13132 26200 13141
rect 36452 13200 36504 13252
rect 36544 13243 36596 13252
rect 36544 13209 36553 13243
rect 36553 13209 36587 13243
rect 36587 13209 36596 13243
rect 36544 13200 36596 13209
rect 32496 13132 32548 13184
rect 38844 13200 38896 13252
rect 41420 13132 41472 13184
rect 43076 13311 43128 13320
rect 43076 13277 43085 13311
rect 43085 13277 43119 13311
rect 43119 13277 43128 13311
rect 43076 13268 43128 13277
rect 44180 13311 44232 13320
rect 44180 13277 44189 13311
rect 44189 13277 44223 13311
rect 44223 13277 44232 13311
rect 44180 13268 44232 13277
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 4896 12928 4948 12980
rect 6092 12928 6144 12980
rect 7656 12928 7708 12980
rect 7748 12860 7800 12912
rect 7104 12792 7156 12844
rect 6460 12724 6512 12776
rect 8300 12724 8352 12776
rect 5632 12656 5684 12708
rect 6092 12656 6144 12708
rect 8668 12724 8720 12776
rect 11428 12928 11480 12980
rect 13728 12928 13780 12980
rect 20168 12928 20220 12980
rect 22008 12971 22060 12980
rect 22008 12937 22017 12971
rect 22017 12937 22051 12971
rect 22051 12937 22060 12971
rect 22008 12928 22060 12937
rect 22468 12971 22520 12980
rect 22468 12937 22477 12971
rect 22477 12937 22511 12971
rect 22511 12937 22520 12971
rect 22468 12928 22520 12937
rect 24860 12928 24912 12980
rect 26332 12971 26384 12980
rect 26332 12937 26341 12971
rect 26341 12937 26375 12971
rect 26375 12937 26384 12971
rect 26332 12928 26384 12937
rect 27712 12971 27764 12980
rect 27712 12937 27721 12971
rect 27721 12937 27755 12971
rect 27755 12937 27764 12971
rect 27712 12928 27764 12937
rect 12716 12860 12768 12912
rect 13820 12860 13872 12912
rect 10416 12835 10468 12844
rect 10416 12801 10425 12835
rect 10425 12801 10459 12835
rect 10459 12801 10468 12835
rect 10416 12792 10468 12801
rect 10600 12835 10652 12844
rect 10600 12801 10609 12835
rect 10609 12801 10643 12835
rect 10643 12801 10652 12835
rect 10600 12792 10652 12801
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 15752 12860 15804 12912
rect 17868 12860 17920 12912
rect 18604 12860 18656 12912
rect 19156 12860 19208 12912
rect 15200 12835 15252 12844
rect 15200 12801 15209 12835
rect 15209 12801 15243 12835
rect 15243 12801 15252 12835
rect 15200 12792 15252 12801
rect 18236 12792 18288 12844
rect 18696 12792 18748 12844
rect 19340 12792 19392 12844
rect 15292 12767 15344 12776
rect 15292 12733 15301 12767
rect 15301 12733 15335 12767
rect 15335 12733 15344 12767
rect 15292 12724 15344 12733
rect 8484 12588 8536 12640
rect 8668 12588 8720 12640
rect 12624 12699 12676 12708
rect 12624 12665 12633 12699
rect 12633 12665 12667 12699
rect 12667 12665 12676 12699
rect 12624 12656 12676 12665
rect 13084 12656 13136 12708
rect 17776 12724 17828 12776
rect 19616 12835 19668 12844
rect 19616 12801 19625 12835
rect 19625 12801 19659 12835
rect 19659 12801 19668 12835
rect 25320 12860 25372 12912
rect 26148 12860 26200 12912
rect 36544 12928 36596 12980
rect 40040 12928 40092 12980
rect 43352 12928 43404 12980
rect 43720 12971 43772 12980
rect 43720 12937 43729 12971
rect 43729 12937 43763 12971
rect 43763 12937 43772 12971
rect 43720 12928 43772 12937
rect 33324 12860 33376 12912
rect 33784 12860 33836 12912
rect 35532 12860 35584 12912
rect 36360 12860 36412 12912
rect 38476 12860 38528 12912
rect 41236 12860 41288 12912
rect 44364 12860 44416 12912
rect 48964 12860 49016 12912
rect 19616 12792 19668 12801
rect 20352 12792 20404 12844
rect 20720 12835 20772 12844
rect 20720 12801 20729 12835
rect 20729 12801 20763 12835
rect 20763 12801 20772 12835
rect 20720 12792 20772 12801
rect 21916 12792 21968 12844
rect 26240 12792 26292 12844
rect 26424 12792 26476 12844
rect 26516 12792 26568 12844
rect 33416 12792 33468 12844
rect 38568 12792 38620 12844
rect 38752 12835 38804 12844
rect 38752 12801 38761 12835
rect 38761 12801 38795 12835
rect 38795 12801 38804 12835
rect 38752 12792 38804 12801
rect 40316 12835 40368 12844
rect 40316 12801 40325 12835
rect 40325 12801 40359 12835
rect 40359 12801 40368 12835
rect 40316 12792 40368 12801
rect 43628 12792 43680 12844
rect 48596 12835 48648 12844
rect 48596 12801 48605 12835
rect 48605 12801 48639 12835
rect 48639 12801 48648 12835
rect 48596 12792 48648 12801
rect 20168 12724 20220 12776
rect 22652 12767 22704 12776
rect 22652 12733 22661 12767
rect 22661 12733 22695 12767
rect 22695 12733 22704 12767
rect 22652 12724 22704 12733
rect 23112 12724 23164 12776
rect 24860 12724 24912 12776
rect 25596 12724 25648 12776
rect 27068 12767 27120 12776
rect 27068 12733 27077 12767
rect 27077 12733 27111 12767
rect 27111 12733 27120 12767
rect 27068 12724 27120 12733
rect 33600 12767 33652 12776
rect 16396 12656 16448 12708
rect 25688 12656 25740 12708
rect 27436 12656 27488 12708
rect 33600 12733 33609 12767
rect 33609 12733 33643 12767
rect 33643 12733 33652 12767
rect 33600 12724 33652 12733
rect 33692 12724 33744 12776
rect 33876 12724 33928 12776
rect 49424 12724 49476 12776
rect 28816 12656 28868 12708
rect 14924 12631 14976 12640
rect 14924 12597 14933 12631
rect 14933 12597 14967 12631
rect 14967 12597 14976 12631
rect 14924 12588 14976 12597
rect 16304 12588 16356 12640
rect 19340 12588 19392 12640
rect 19616 12588 19668 12640
rect 20444 12588 20496 12640
rect 21272 12631 21324 12640
rect 21272 12597 21281 12631
rect 21281 12597 21315 12631
rect 21315 12597 21324 12631
rect 21272 12588 21324 12597
rect 24952 12588 25004 12640
rect 33140 12631 33192 12640
rect 33140 12597 33149 12631
rect 33149 12597 33183 12631
rect 33183 12597 33192 12631
rect 33140 12588 33192 12597
rect 37740 12631 37792 12640
rect 37740 12597 37749 12631
rect 37749 12597 37783 12631
rect 37783 12597 37792 12631
rect 37740 12588 37792 12597
rect 38200 12588 38252 12640
rect 49056 12588 49108 12640
rect 50160 12588 50212 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 65654 12486 65706 12538
rect 65718 12486 65770 12538
rect 65782 12486 65834 12538
rect 65846 12486 65898 12538
rect 65910 12486 65962 12538
rect 8300 12384 8352 12436
rect 8668 12384 8720 12436
rect 10416 12384 10468 12436
rect 12716 12427 12768 12436
rect 12716 12393 12725 12427
rect 12725 12393 12759 12427
rect 12759 12393 12768 12427
rect 12716 12384 12768 12393
rect 12808 12384 12860 12436
rect 16028 12384 16080 12436
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 20168 12427 20220 12436
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 20904 12384 20956 12436
rect 21088 12384 21140 12436
rect 21916 12427 21968 12436
rect 21916 12393 21925 12427
rect 21925 12393 21959 12427
rect 21959 12393 21968 12427
rect 21916 12384 21968 12393
rect 29276 12384 29328 12436
rect 7932 12316 7984 12368
rect 15200 12316 15252 12368
rect 16396 12316 16448 12368
rect 4712 12248 4764 12300
rect 7380 12291 7432 12300
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 9312 12291 9364 12300
rect 9312 12257 9321 12291
rect 9321 12257 9355 12291
rect 9355 12257 9364 12291
rect 9312 12248 9364 12257
rect 21732 12316 21784 12368
rect 5632 12180 5684 12232
rect 5264 12112 5316 12164
rect 7104 12155 7156 12164
rect 7104 12121 7113 12155
rect 7113 12121 7147 12155
rect 7147 12121 7156 12155
rect 7104 12112 7156 12121
rect 6736 12087 6788 12096
rect 6736 12053 6745 12087
rect 6745 12053 6779 12087
rect 6779 12053 6788 12087
rect 6736 12044 6788 12053
rect 8668 12180 8720 12232
rect 10416 12180 10468 12232
rect 12256 12180 12308 12232
rect 16304 12223 16356 12232
rect 16304 12189 16308 12223
rect 16308 12189 16342 12223
rect 16342 12189 16356 12223
rect 16304 12180 16356 12189
rect 17776 12248 17828 12300
rect 36084 12291 36136 12300
rect 36084 12257 36093 12291
rect 36093 12257 36127 12291
rect 36127 12257 36136 12291
rect 36084 12248 36136 12257
rect 37740 12384 37792 12436
rect 38752 12384 38804 12436
rect 40316 12316 40368 12368
rect 47952 12316 48004 12368
rect 48872 12427 48924 12436
rect 48872 12393 48881 12427
rect 48881 12393 48915 12427
rect 48915 12393 48924 12427
rect 48872 12384 48924 12393
rect 48964 12316 49016 12368
rect 36360 12291 36412 12300
rect 36360 12257 36369 12291
rect 36369 12257 36403 12291
rect 36403 12257 36412 12291
rect 36360 12248 36412 12257
rect 16580 12223 16632 12232
rect 16580 12189 16625 12223
rect 16625 12189 16632 12223
rect 16580 12180 16632 12189
rect 16764 12223 16816 12232
rect 16764 12189 16773 12223
rect 16773 12189 16807 12223
rect 16807 12189 16816 12223
rect 19432 12223 19484 12232
rect 16764 12180 16816 12189
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 8576 12112 8628 12164
rect 15016 12112 15068 12164
rect 15292 12112 15344 12164
rect 20904 12180 20956 12232
rect 21272 12180 21324 12232
rect 23480 12180 23532 12232
rect 23756 12180 23808 12232
rect 24676 12180 24728 12232
rect 25228 12223 25280 12232
rect 25228 12189 25237 12223
rect 25237 12189 25271 12223
rect 25271 12189 25280 12223
rect 25228 12180 25280 12189
rect 25596 12223 25648 12232
rect 25596 12189 25605 12223
rect 25605 12189 25639 12223
rect 25639 12189 25648 12223
rect 25596 12180 25648 12189
rect 26148 12223 26200 12232
rect 26148 12189 26157 12223
rect 26157 12189 26191 12223
rect 26191 12189 26200 12223
rect 26148 12180 26200 12189
rect 26608 12223 26660 12232
rect 26608 12189 26617 12223
rect 26617 12189 26651 12223
rect 26651 12189 26660 12223
rect 26608 12180 26660 12189
rect 26792 12223 26844 12232
rect 26792 12189 26801 12223
rect 26801 12189 26835 12223
rect 26835 12189 26844 12223
rect 26792 12180 26844 12189
rect 31300 12180 31352 12232
rect 36912 12180 36964 12232
rect 37188 12180 37240 12232
rect 20444 12155 20496 12164
rect 7288 12044 7340 12096
rect 8760 12044 8812 12096
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 11060 12087 11112 12096
rect 11060 12053 11069 12087
rect 11069 12053 11103 12087
rect 11103 12053 11112 12087
rect 11060 12044 11112 12053
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 14832 12044 14884 12096
rect 16672 12044 16724 12096
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 19248 12087 19300 12096
rect 19248 12053 19257 12087
rect 19257 12053 19291 12087
rect 19291 12053 19300 12087
rect 19248 12044 19300 12053
rect 20444 12121 20453 12155
rect 20453 12121 20487 12155
rect 20487 12121 20496 12155
rect 20444 12112 20496 12121
rect 32036 12112 32088 12164
rect 20628 12044 20680 12096
rect 20996 12044 21048 12096
rect 24400 12044 24452 12096
rect 31668 12087 31720 12096
rect 31668 12053 31677 12087
rect 31677 12053 31711 12087
rect 31711 12053 31720 12087
rect 31668 12044 31720 12053
rect 32864 12112 32916 12164
rect 33048 12112 33100 12164
rect 37372 12180 37424 12232
rect 38200 12180 38252 12232
rect 38568 12223 38620 12232
rect 38568 12189 38577 12223
rect 38577 12189 38611 12223
rect 38611 12189 38620 12223
rect 38568 12180 38620 12189
rect 40132 12180 40184 12232
rect 43720 12180 43772 12232
rect 44272 12180 44324 12232
rect 45468 12180 45520 12232
rect 48044 12223 48096 12232
rect 48044 12189 48053 12223
rect 48053 12189 48087 12223
rect 48087 12189 48096 12223
rect 48044 12180 48096 12189
rect 33968 12044 34020 12096
rect 36912 12044 36964 12096
rect 48136 12112 48188 12164
rect 49056 12155 49108 12164
rect 49056 12121 49065 12155
rect 49065 12121 49099 12155
rect 49099 12121 49108 12155
rect 49056 12112 49108 12121
rect 38292 12044 38344 12096
rect 40684 12044 40736 12096
rect 41328 12044 41380 12096
rect 45100 12087 45152 12096
rect 45100 12053 45109 12087
rect 45109 12053 45143 12087
rect 45143 12053 45152 12087
rect 45100 12044 45152 12053
rect 45560 12044 45612 12096
rect 46848 12044 46900 12096
rect 48320 12044 48372 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 5264 11883 5316 11892
rect 5264 11849 5273 11883
rect 5273 11849 5307 11883
rect 5307 11849 5316 11883
rect 5264 11840 5316 11849
rect 8116 11840 8168 11892
rect 10416 11883 10468 11892
rect 10416 11849 10425 11883
rect 10425 11849 10459 11883
rect 10459 11849 10468 11883
rect 10416 11840 10468 11849
rect 16764 11840 16816 11892
rect 8392 11772 8444 11824
rect 6736 11704 6788 11756
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 8300 11704 8352 11756
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 11980 11772 12032 11824
rect 17960 11840 18012 11892
rect 18512 11840 18564 11892
rect 20444 11883 20496 11892
rect 20444 11849 20453 11883
rect 20453 11849 20487 11883
rect 20487 11849 20496 11883
rect 20444 11840 20496 11849
rect 25320 11840 25372 11892
rect 26884 11840 26936 11892
rect 11244 11704 11296 11756
rect 17868 11772 17920 11824
rect 8116 11679 8168 11688
rect 8116 11645 8125 11679
rect 8125 11645 8159 11679
rect 8159 11645 8168 11679
rect 8116 11636 8168 11645
rect 10692 11679 10744 11688
rect 10692 11645 10701 11679
rect 10701 11645 10735 11679
rect 10735 11645 10744 11679
rect 10692 11636 10744 11645
rect 11060 11636 11112 11688
rect 11520 11636 11572 11688
rect 12624 11568 12676 11620
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 19248 11704 19300 11756
rect 20812 11704 20864 11756
rect 20996 11747 21048 11756
rect 20996 11713 21005 11747
rect 21005 11713 21039 11747
rect 21039 11713 21048 11747
rect 20996 11704 21048 11713
rect 25228 11772 25280 11824
rect 32128 11772 32180 11824
rect 37280 11840 37332 11892
rect 37740 11840 37792 11892
rect 38476 11840 38528 11892
rect 41604 11840 41656 11892
rect 42156 11840 42208 11892
rect 45560 11840 45612 11892
rect 48044 11840 48096 11892
rect 49240 11840 49292 11892
rect 49700 11840 49752 11892
rect 38292 11815 38344 11824
rect 24400 11704 24452 11756
rect 24952 11704 25004 11756
rect 26240 11747 26292 11756
rect 26240 11713 26249 11747
rect 26249 11713 26283 11747
rect 26283 11713 26292 11747
rect 26976 11747 27028 11756
rect 26240 11704 26292 11713
rect 26976 11713 26985 11747
rect 26985 11713 27019 11747
rect 27019 11713 27028 11747
rect 26976 11704 27028 11713
rect 27436 11704 27488 11756
rect 28908 11747 28960 11756
rect 28908 11713 28917 11747
rect 28917 11713 28951 11747
rect 28951 11713 28960 11747
rect 28908 11704 28960 11713
rect 15660 11679 15712 11688
rect 15660 11645 15669 11679
rect 15669 11645 15703 11679
rect 15703 11645 15712 11679
rect 15660 11636 15712 11645
rect 16304 11636 16356 11688
rect 23296 11679 23348 11688
rect 14924 11568 14976 11620
rect 7288 11543 7340 11552
rect 7288 11509 7297 11543
rect 7297 11509 7331 11543
rect 7331 11509 7340 11543
rect 7288 11500 7340 11509
rect 8116 11500 8168 11552
rect 9496 11500 9548 11552
rect 14740 11500 14792 11552
rect 15292 11500 15344 11552
rect 16672 11500 16724 11552
rect 23296 11645 23305 11679
rect 23305 11645 23339 11679
rect 23339 11645 23348 11679
rect 23296 11636 23348 11645
rect 25044 11636 25096 11688
rect 28816 11679 28868 11688
rect 28816 11645 28825 11679
rect 28825 11645 28859 11679
rect 28859 11645 28868 11679
rect 28816 11636 28868 11645
rect 19800 11500 19852 11552
rect 19984 11543 20036 11552
rect 19984 11509 19993 11543
rect 19993 11509 20027 11543
rect 20027 11509 20036 11543
rect 19984 11500 20036 11509
rect 20720 11543 20772 11552
rect 20720 11509 20729 11543
rect 20729 11509 20763 11543
rect 20763 11509 20772 11543
rect 20720 11500 20772 11509
rect 26608 11568 26660 11620
rect 29000 11568 29052 11620
rect 30656 11747 30708 11756
rect 30656 11713 30665 11747
rect 30665 11713 30699 11747
rect 30699 11713 30708 11747
rect 30656 11704 30708 11713
rect 30932 11747 30984 11756
rect 30932 11713 30941 11747
rect 30941 11713 30975 11747
rect 30975 11713 30984 11747
rect 30932 11704 30984 11713
rect 31116 11747 31168 11756
rect 31116 11713 31125 11747
rect 31125 11713 31159 11747
rect 31159 11713 31168 11747
rect 31116 11704 31168 11713
rect 31392 11747 31444 11756
rect 31392 11713 31401 11747
rect 31401 11713 31435 11747
rect 31435 11713 31444 11747
rect 31392 11704 31444 11713
rect 33140 11704 33192 11756
rect 33784 11704 33836 11756
rect 38292 11781 38301 11815
rect 38301 11781 38335 11815
rect 38335 11781 38344 11815
rect 38292 11772 38344 11781
rect 48136 11772 48188 11824
rect 33048 11636 33100 11688
rect 33140 11568 33192 11620
rect 31392 11500 31444 11552
rect 33600 11500 33652 11552
rect 34704 11500 34756 11552
rect 36084 11500 36136 11552
rect 36912 11636 36964 11688
rect 41420 11704 41472 11756
rect 41880 11704 41932 11756
rect 45468 11704 45520 11756
rect 47952 11704 48004 11756
rect 48504 11747 48556 11756
rect 48504 11713 48513 11747
rect 48513 11713 48547 11747
rect 48547 11713 48556 11747
rect 48504 11704 48556 11713
rect 49148 11704 49200 11756
rect 49240 11747 49292 11756
rect 49240 11713 49249 11747
rect 49249 11713 49283 11747
rect 49283 11713 49292 11747
rect 49240 11704 49292 11713
rect 49424 11747 49476 11756
rect 49424 11713 49433 11747
rect 49433 11713 49467 11747
rect 49467 11713 49476 11747
rect 49884 11747 49936 11756
rect 49424 11704 49476 11713
rect 49884 11713 49893 11747
rect 49893 11713 49927 11747
rect 49927 11713 49936 11747
rect 49884 11704 49936 11713
rect 67364 11747 67416 11756
rect 43904 11679 43956 11688
rect 43904 11645 43913 11679
rect 43913 11645 43947 11679
rect 43947 11645 43956 11679
rect 43904 11636 43956 11645
rect 46756 11568 46808 11620
rect 48596 11568 48648 11620
rect 37832 11500 37884 11552
rect 42708 11500 42760 11552
rect 46940 11500 46992 11552
rect 48872 11500 48924 11552
rect 67364 11713 67373 11747
rect 67373 11713 67407 11747
rect 67407 11713 67416 11747
rect 67364 11704 67416 11713
rect 67548 11543 67600 11552
rect 67548 11509 67557 11543
rect 67557 11509 67591 11543
rect 67591 11509 67600 11543
rect 67548 11500 67600 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 65654 11398 65706 11450
rect 65718 11398 65770 11450
rect 65782 11398 65834 11450
rect 65846 11398 65898 11450
rect 65910 11398 65962 11450
rect 7288 11296 7340 11348
rect 8392 11296 8444 11348
rect 11244 11339 11296 11348
rect 11244 11305 11253 11339
rect 11253 11305 11287 11339
rect 11287 11305 11296 11339
rect 11244 11296 11296 11305
rect 12256 11339 12308 11348
rect 12256 11305 12265 11339
rect 12265 11305 12299 11339
rect 12299 11305 12308 11339
rect 12256 11296 12308 11305
rect 14832 11296 14884 11348
rect 4712 11160 4764 11212
rect 6736 11160 6788 11212
rect 7932 11160 7984 11212
rect 5172 11024 5224 11076
rect 8484 11160 8536 11212
rect 13452 11228 13504 11280
rect 16764 11228 16816 11280
rect 18604 11228 18656 11280
rect 19432 11296 19484 11348
rect 19800 11296 19852 11348
rect 21180 11296 21232 11348
rect 13084 11160 13136 11212
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 14740 11160 14792 11169
rect 16856 11160 16908 11212
rect 21088 11228 21140 11280
rect 8392 11092 8444 11144
rect 12624 11135 12676 11144
rect 12624 11101 12633 11135
rect 12633 11101 12667 11135
rect 12667 11101 12676 11135
rect 12624 11092 12676 11101
rect 8576 11024 8628 11076
rect 9496 10999 9548 11008
rect 9496 10965 9505 10999
rect 9505 10965 9539 10999
rect 9539 10965 9548 10999
rect 9496 10956 9548 10965
rect 9588 10956 9640 11008
rect 16948 11024 17000 11076
rect 17132 11067 17184 11076
rect 17132 11033 17141 11067
rect 17141 11033 17175 11067
rect 17175 11033 17184 11067
rect 17132 11024 17184 11033
rect 20076 11160 20128 11212
rect 20536 11160 20588 11212
rect 19984 11092 20036 11144
rect 23296 11296 23348 11348
rect 28908 11296 28960 11348
rect 29000 11296 29052 11348
rect 30196 11296 30248 11348
rect 31300 11339 31352 11348
rect 31300 11305 31309 11339
rect 31309 11305 31343 11339
rect 31343 11305 31352 11339
rect 31300 11296 31352 11305
rect 33784 11339 33836 11348
rect 33784 11305 33793 11339
rect 33793 11305 33827 11339
rect 33827 11305 33836 11339
rect 33784 11296 33836 11305
rect 36084 11296 36136 11348
rect 38568 11296 38620 11348
rect 43812 11296 43864 11348
rect 44180 11296 44232 11348
rect 46756 11339 46808 11348
rect 46756 11305 46765 11339
rect 46765 11305 46799 11339
rect 46799 11305 46808 11339
rect 46756 11296 46808 11305
rect 48136 11339 48188 11348
rect 48136 11305 48145 11339
rect 48145 11305 48179 11339
rect 48179 11305 48188 11339
rect 48136 11296 48188 11305
rect 49884 11296 49936 11348
rect 67364 11339 67416 11348
rect 21916 11228 21968 11280
rect 23572 11228 23624 11280
rect 26792 11228 26844 11280
rect 28264 11271 28316 11280
rect 28264 11237 28273 11271
rect 28273 11237 28307 11271
rect 28307 11237 28316 11271
rect 28264 11228 28316 11237
rect 29460 11228 29512 11280
rect 33140 11228 33192 11280
rect 22100 11160 22152 11212
rect 22652 11160 22704 11212
rect 24860 11135 24912 11144
rect 21180 11024 21232 11076
rect 24860 11101 24869 11135
rect 24869 11101 24903 11135
rect 24903 11101 24912 11135
rect 24860 11092 24912 11101
rect 25228 11160 25280 11212
rect 26332 11160 26384 11212
rect 28080 11160 28132 11212
rect 29092 11160 29144 11212
rect 24492 11024 24544 11076
rect 26240 11135 26292 11144
rect 26240 11101 26249 11135
rect 26249 11101 26283 11135
rect 26283 11101 26292 11135
rect 26240 11092 26292 11101
rect 30472 11092 30524 11144
rect 31208 11092 31260 11144
rect 29184 11024 29236 11076
rect 30748 11024 30800 11076
rect 36912 11160 36964 11212
rect 31668 11092 31720 11144
rect 33048 11092 33100 11144
rect 33600 11135 33652 11144
rect 33600 11101 33609 11135
rect 33609 11101 33643 11135
rect 33643 11101 33652 11135
rect 33600 11092 33652 11101
rect 37280 11135 37332 11144
rect 37280 11101 37289 11135
rect 37289 11101 37323 11135
rect 37323 11101 37332 11135
rect 37280 11092 37332 11101
rect 38200 11203 38252 11212
rect 38200 11169 38209 11203
rect 38209 11169 38243 11203
rect 38243 11169 38252 11203
rect 38200 11160 38252 11169
rect 38936 11160 38988 11212
rect 41604 11203 41656 11212
rect 41604 11169 41613 11203
rect 41613 11169 41647 11203
rect 41647 11169 41656 11203
rect 41604 11160 41656 11169
rect 43904 11160 43956 11212
rect 48044 11228 48096 11280
rect 48964 11228 49016 11280
rect 67364 11305 67373 11339
rect 67373 11305 67407 11339
rect 67407 11305 67416 11339
rect 67364 11296 67416 11305
rect 50620 11228 50672 11280
rect 38384 11092 38436 11144
rect 16764 10956 16816 11008
rect 19984 10956 20036 11008
rect 21364 10999 21416 11008
rect 21364 10965 21373 10999
rect 21373 10965 21407 10999
rect 21407 10965 21416 10999
rect 21364 10956 21416 10965
rect 33692 11024 33744 11076
rect 36176 11067 36228 11076
rect 36176 11033 36185 11067
rect 36185 11033 36219 11067
rect 36219 11033 36228 11067
rect 36176 11024 36228 11033
rect 39856 11092 39908 11144
rect 42156 11135 42208 11144
rect 42156 11101 42165 11135
rect 42165 11101 42199 11135
rect 42199 11101 42208 11135
rect 42156 11092 42208 11101
rect 42708 11092 42760 11144
rect 44272 11135 44324 11144
rect 44272 11101 44281 11135
rect 44281 11101 44315 11135
rect 44315 11101 44324 11135
rect 44272 11092 44324 11101
rect 47400 11135 47452 11144
rect 47400 11101 47409 11135
rect 47409 11101 47443 11135
rect 47443 11101 47452 11135
rect 47400 11092 47452 11101
rect 48320 11160 48372 11212
rect 40776 11024 40828 11076
rect 47032 11024 47084 11076
rect 48504 11092 48556 11144
rect 48964 11092 49016 11144
rect 49148 11092 49200 11144
rect 49976 11092 50028 11144
rect 50160 11067 50212 11076
rect 50160 11033 50169 11067
rect 50169 11033 50203 11067
rect 50203 11033 50212 11067
rect 50160 11024 50212 11033
rect 49424 10956 49476 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 5172 10795 5224 10804
rect 5172 10761 5181 10795
rect 5181 10761 5215 10795
rect 5215 10761 5224 10795
rect 5172 10752 5224 10761
rect 6736 10795 6788 10804
rect 6736 10761 6745 10795
rect 6745 10761 6779 10795
rect 6779 10761 6788 10795
rect 6736 10752 6788 10761
rect 9588 10752 9640 10804
rect 13728 10795 13780 10804
rect 8300 10684 8352 10736
rect 12900 10684 12952 10736
rect 13728 10761 13737 10795
rect 13737 10761 13771 10795
rect 13771 10761 13780 10795
rect 13728 10752 13780 10761
rect 16764 10795 16816 10804
rect 16764 10761 16773 10795
rect 16773 10761 16807 10795
rect 16807 10761 16816 10795
rect 16764 10752 16816 10761
rect 20352 10795 20404 10804
rect 20352 10761 20361 10795
rect 20361 10761 20395 10795
rect 20395 10761 20404 10795
rect 20352 10752 20404 10761
rect 21916 10795 21968 10804
rect 21916 10761 21925 10795
rect 21925 10761 21959 10795
rect 21959 10761 21968 10795
rect 21916 10752 21968 10761
rect 22008 10752 22060 10804
rect 22928 10752 22980 10804
rect 30656 10752 30708 10804
rect 31944 10752 31996 10804
rect 33508 10795 33560 10804
rect 33508 10761 33517 10795
rect 33517 10761 33551 10795
rect 33551 10761 33560 10795
rect 33508 10752 33560 10761
rect 33600 10752 33652 10804
rect 38936 10752 38988 10804
rect 40776 10795 40828 10804
rect 40776 10761 40785 10795
rect 40785 10761 40819 10795
rect 40819 10761 40828 10795
rect 40776 10752 40828 10761
rect 42708 10752 42760 10804
rect 6460 10616 6512 10668
rect 8116 10659 8168 10668
rect 8116 10625 8125 10659
rect 8125 10625 8159 10659
rect 8159 10625 8168 10659
rect 8116 10616 8168 10625
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 12164 10659 12216 10668
rect 12164 10625 12198 10659
rect 12198 10625 12216 10659
rect 23480 10684 23532 10736
rect 30840 10684 30892 10736
rect 12164 10616 12216 10625
rect 15660 10616 15712 10668
rect 20812 10659 20864 10668
rect 20812 10625 20821 10659
rect 20821 10625 20855 10659
rect 20855 10625 20864 10659
rect 20812 10616 20864 10625
rect 26424 10616 26476 10668
rect 26976 10616 27028 10668
rect 30748 10616 30800 10668
rect 34704 10684 34756 10736
rect 31484 10616 31536 10668
rect 32312 10659 32364 10668
rect 32312 10625 32321 10659
rect 32321 10625 32355 10659
rect 32355 10625 32364 10659
rect 32312 10616 32364 10625
rect 32588 10659 32640 10668
rect 32588 10625 32597 10659
rect 32597 10625 32631 10659
rect 32631 10625 32640 10659
rect 38200 10684 38252 10736
rect 38384 10684 38436 10736
rect 32588 10616 32640 10625
rect 37832 10659 37884 10668
rect 37832 10625 37841 10659
rect 37841 10625 37875 10659
rect 37875 10625 37884 10659
rect 37832 10616 37884 10625
rect 40500 10616 40552 10668
rect 41420 10616 41472 10668
rect 46940 10752 46992 10804
rect 47032 10795 47084 10804
rect 47032 10761 47041 10795
rect 47041 10761 47075 10795
rect 47075 10761 47084 10795
rect 47032 10752 47084 10761
rect 47400 10752 47452 10804
rect 49424 10752 49476 10804
rect 45100 10684 45152 10736
rect 50068 10684 50120 10736
rect 46848 10659 46900 10668
rect 46848 10625 46857 10659
rect 46857 10625 46891 10659
rect 46891 10625 46900 10659
rect 46848 10616 46900 10625
rect 48596 10659 48648 10668
rect 11520 10548 11572 10600
rect 16580 10548 16632 10600
rect 20536 10591 20588 10600
rect 20536 10557 20545 10591
rect 20545 10557 20579 10591
rect 20579 10557 20588 10591
rect 20536 10548 20588 10557
rect 8392 10523 8444 10532
rect 8392 10489 8401 10523
rect 8401 10489 8435 10523
rect 8435 10489 8444 10523
rect 8392 10480 8444 10489
rect 6828 10412 6880 10464
rect 7656 10455 7708 10464
rect 7656 10421 7665 10455
rect 7665 10421 7699 10455
rect 7699 10421 7708 10455
rect 7656 10412 7708 10421
rect 11796 10412 11848 10464
rect 20260 10480 20312 10532
rect 21364 10548 21416 10600
rect 25964 10591 26016 10600
rect 25964 10557 25973 10591
rect 25973 10557 26007 10591
rect 26007 10557 26016 10591
rect 25964 10548 26016 10557
rect 26148 10548 26200 10600
rect 29184 10591 29236 10600
rect 29184 10557 29193 10591
rect 29193 10557 29227 10591
rect 29227 10557 29236 10591
rect 29184 10548 29236 10557
rect 20996 10480 21048 10532
rect 20628 10412 20680 10464
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 33692 10548 33744 10600
rect 43628 10548 43680 10600
rect 46756 10548 46808 10600
rect 48596 10625 48605 10659
rect 48605 10625 48639 10659
rect 48639 10625 48648 10659
rect 48596 10616 48648 10625
rect 50160 10659 50212 10668
rect 49792 10548 49844 10600
rect 50160 10625 50169 10659
rect 50169 10625 50203 10659
rect 50203 10625 50212 10659
rect 50160 10616 50212 10625
rect 50620 10659 50672 10668
rect 50620 10625 50629 10659
rect 50629 10625 50663 10659
rect 50663 10625 50672 10659
rect 50620 10616 50672 10625
rect 50804 10659 50856 10668
rect 50804 10625 50813 10659
rect 50813 10625 50847 10659
rect 50847 10625 50856 10659
rect 50804 10616 50856 10625
rect 40592 10480 40644 10532
rect 43536 10480 43588 10532
rect 49424 10480 49476 10532
rect 49608 10480 49660 10532
rect 50712 10548 50764 10600
rect 29552 10412 29604 10464
rect 30380 10412 30432 10464
rect 30840 10412 30892 10464
rect 31852 10412 31904 10464
rect 39028 10412 39080 10464
rect 42616 10455 42668 10464
rect 42616 10421 42625 10455
rect 42625 10421 42659 10455
rect 42659 10421 42668 10455
rect 42616 10412 42668 10421
rect 48412 10455 48464 10464
rect 48412 10421 48421 10455
rect 48421 10421 48455 10455
rect 48455 10421 48464 10455
rect 48412 10412 48464 10421
rect 50896 10412 50948 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 65654 10310 65706 10362
rect 65718 10310 65770 10362
rect 65782 10310 65834 10362
rect 65846 10310 65898 10362
rect 65910 10310 65962 10362
rect 7656 10208 7708 10260
rect 9128 10140 9180 10192
rect 12164 10208 12216 10260
rect 17132 10208 17184 10260
rect 20536 10208 20588 10260
rect 21548 10208 21600 10260
rect 25964 10251 26016 10260
rect 25964 10217 25973 10251
rect 25973 10217 26007 10251
rect 26007 10217 26016 10251
rect 25964 10208 26016 10217
rect 26240 10208 26292 10260
rect 29184 10208 29236 10260
rect 30932 10208 30984 10260
rect 31208 10251 31260 10260
rect 31208 10217 31217 10251
rect 31217 10217 31251 10251
rect 31251 10217 31260 10251
rect 31208 10208 31260 10217
rect 33508 10208 33560 10260
rect 40500 10251 40552 10260
rect 40500 10217 40509 10251
rect 40509 10217 40543 10251
rect 40543 10217 40552 10251
rect 40500 10208 40552 10217
rect 46848 10208 46900 10260
rect 48504 10208 48556 10260
rect 48596 10208 48648 10260
rect 49792 10208 49844 10260
rect 50252 10208 50304 10260
rect 16120 10183 16172 10192
rect 6552 10115 6604 10124
rect 6552 10081 6561 10115
rect 6561 10081 6595 10115
rect 6595 10081 6604 10115
rect 6552 10072 6604 10081
rect 8116 10072 8168 10124
rect 8944 10115 8996 10124
rect 8944 10081 8953 10115
rect 8953 10081 8987 10115
rect 8987 10081 8996 10115
rect 8944 10072 8996 10081
rect 9496 10072 9548 10124
rect 16120 10149 16129 10183
rect 16129 10149 16163 10183
rect 16163 10149 16172 10183
rect 16120 10140 16172 10149
rect 16580 10140 16632 10192
rect 13084 10115 13136 10124
rect 8208 10004 8260 10056
rect 9036 10047 9088 10056
rect 9036 10013 9045 10047
rect 9045 10013 9079 10047
rect 9079 10013 9088 10047
rect 9036 10004 9088 10013
rect 9128 10004 9180 10056
rect 8300 9936 8352 9988
rect 13084 10081 13093 10115
rect 13093 10081 13127 10115
rect 13127 10081 13136 10115
rect 13084 10072 13136 10081
rect 15660 10072 15712 10124
rect 16948 10072 17000 10124
rect 18052 10072 18104 10124
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 18696 10140 18748 10192
rect 21548 10072 21600 10124
rect 21180 10004 21232 10056
rect 24124 10072 24176 10124
rect 24584 10047 24636 10056
rect 19892 9936 19944 9988
rect 24584 10013 24593 10047
rect 24593 10013 24627 10047
rect 24627 10013 24636 10047
rect 24584 10004 24636 10013
rect 29552 10140 29604 10192
rect 34428 10140 34480 10192
rect 29184 10072 29236 10124
rect 32128 10115 32180 10124
rect 26424 10004 26476 10056
rect 30380 10047 30432 10056
rect 30380 10013 30389 10047
rect 30389 10013 30423 10047
rect 30423 10013 30432 10047
rect 30380 10004 30432 10013
rect 30656 10047 30708 10056
rect 30656 10013 30665 10047
rect 30665 10013 30699 10047
rect 30699 10013 30708 10047
rect 30656 10004 30708 10013
rect 31116 10004 31168 10056
rect 32128 10081 32137 10115
rect 32137 10081 32171 10115
rect 32171 10081 32180 10115
rect 32128 10072 32180 10081
rect 32588 10072 32640 10124
rect 41236 10140 41288 10192
rect 49148 10140 49200 10192
rect 49516 10183 49568 10192
rect 49516 10149 49525 10183
rect 49525 10149 49559 10183
rect 49559 10149 49568 10183
rect 49516 10140 49568 10149
rect 41420 10072 41472 10124
rect 43536 10072 43588 10124
rect 38108 10004 38160 10056
rect 38752 10004 38804 10056
rect 40040 10047 40092 10056
rect 40040 10013 40049 10047
rect 40049 10013 40083 10047
rect 40083 10013 40092 10047
rect 40040 10004 40092 10013
rect 14556 9868 14608 9920
rect 20076 9911 20128 9920
rect 20076 9877 20085 9911
rect 20085 9877 20119 9911
rect 20119 9877 20128 9911
rect 20076 9868 20128 9877
rect 21364 9868 21416 9920
rect 26332 9936 26384 9988
rect 28172 9979 28224 9988
rect 28172 9945 28181 9979
rect 28181 9945 28215 9979
rect 28215 9945 28224 9979
rect 28172 9936 28224 9945
rect 31392 9936 31444 9988
rect 40316 9936 40368 9988
rect 24768 9868 24820 9920
rect 28632 9868 28684 9920
rect 33508 9868 33560 9920
rect 33968 9911 34020 9920
rect 33968 9877 33977 9911
rect 33977 9877 34011 9911
rect 34011 9877 34020 9911
rect 33968 9868 34020 9877
rect 36452 9868 36504 9920
rect 39948 9911 40000 9920
rect 39948 9877 39957 9911
rect 39957 9877 39991 9911
rect 39991 9877 40000 9911
rect 39948 9868 40000 9877
rect 45468 10004 45520 10056
rect 46756 10072 46808 10124
rect 49332 10115 49384 10124
rect 49332 10081 49341 10115
rect 49341 10081 49375 10115
rect 49375 10081 49384 10115
rect 49332 10072 49384 10081
rect 49792 10072 49844 10124
rect 49976 10072 50028 10124
rect 50436 10115 50488 10124
rect 50436 10081 50446 10115
rect 50446 10081 50480 10115
rect 50480 10081 50488 10115
rect 50436 10072 50488 10081
rect 47032 10004 47084 10056
rect 48228 10004 48280 10056
rect 49240 10004 49292 10056
rect 42984 9979 43036 9988
rect 42984 9945 42993 9979
rect 42993 9945 43027 9979
rect 43027 9945 43036 9979
rect 42984 9936 43036 9945
rect 48596 9936 48648 9988
rect 49976 9936 50028 9988
rect 43628 9868 43680 9920
rect 45008 9868 45060 9920
rect 47584 9911 47636 9920
rect 47584 9877 47593 9911
rect 47593 9877 47627 9911
rect 47627 9877 47636 9911
rect 47584 9868 47636 9877
rect 49148 9868 49200 9920
rect 51264 9911 51316 9920
rect 51264 9877 51273 9911
rect 51273 9877 51307 9911
rect 51307 9877 51316 9911
rect 51264 9868 51316 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 8392 9664 8444 9716
rect 8944 9664 8996 9716
rect 16120 9707 16172 9716
rect 16120 9673 16129 9707
rect 16129 9673 16163 9707
rect 16163 9673 16172 9707
rect 16120 9664 16172 9673
rect 20628 9664 20680 9716
rect 25964 9707 26016 9716
rect 25964 9673 25973 9707
rect 25973 9673 26007 9707
rect 26007 9673 26016 9707
rect 25964 9664 26016 9673
rect 32312 9664 32364 9716
rect 33968 9664 34020 9716
rect 38108 9707 38160 9716
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 9036 9596 9088 9648
rect 15384 9596 15436 9648
rect 16672 9639 16724 9648
rect 9312 9571 9364 9580
rect 6552 9503 6604 9512
rect 6552 9469 6561 9503
rect 6561 9469 6595 9503
rect 6595 9469 6604 9503
rect 6552 9460 6604 9469
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 12716 9528 12768 9580
rect 13452 9571 13504 9580
rect 13452 9537 13461 9571
rect 13461 9537 13495 9571
rect 13495 9537 13504 9571
rect 13452 9528 13504 9537
rect 15660 9571 15712 9580
rect 15660 9537 15669 9571
rect 15669 9537 15703 9571
rect 15703 9537 15712 9571
rect 15660 9528 15712 9537
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 16672 9605 16681 9639
rect 16681 9605 16715 9639
rect 16715 9605 16724 9639
rect 16672 9596 16724 9605
rect 17684 9596 17736 9648
rect 10692 9460 10744 9512
rect 10968 9460 11020 9512
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 8300 9392 8352 9444
rect 9128 9392 9180 9444
rect 13636 9435 13688 9444
rect 13636 9401 13645 9435
rect 13645 9401 13679 9435
rect 13679 9401 13688 9435
rect 13636 9392 13688 9401
rect 14740 9392 14792 9444
rect 20076 9528 20128 9580
rect 20628 9528 20680 9580
rect 20904 9528 20956 9580
rect 21916 9528 21968 9580
rect 24584 9596 24636 9648
rect 21180 9460 21232 9512
rect 20536 9392 20588 9444
rect 25780 9528 25832 9580
rect 32128 9639 32180 9648
rect 32128 9605 32137 9639
rect 32137 9605 32171 9639
rect 32171 9605 32180 9639
rect 32128 9596 32180 9605
rect 38108 9673 38117 9707
rect 38117 9673 38151 9707
rect 38151 9673 38160 9707
rect 38108 9664 38160 9673
rect 40040 9664 40092 9716
rect 39948 9596 40000 9648
rect 40316 9596 40368 9648
rect 28264 9528 28316 9580
rect 29828 9528 29880 9580
rect 33324 9528 33376 9580
rect 35348 9528 35400 9580
rect 42984 9664 43036 9716
rect 44180 9596 44232 9648
rect 49240 9664 49292 9716
rect 49976 9664 50028 9716
rect 50620 9664 50672 9716
rect 24492 9503 24544 9512
rect 24492 9469 24501 9503
rect 24501 9469 24535 9503
rect 24535 9469 24544 9503
rect 24492 9460 24544 9469
rect 26240 9460 26292 9512
rect 27988 9503 28040 9512
rect 13728 9324 13780 9376
rect 24124 9367 24176 9376
rect 24124 9333 24133 9367
rect 24133 9333 24167 9367
rect 24167 9333 24176 9367
rect 24124 9324 24176 9333
rect 26424 9324 26476 9376
rect 27988 9469 27997 9503
rect 27997 9469 28031 9503
rect 28031 9469 28040 9503
rect 27988 9460 28040 9469
rect 29644 9460 29696 9512
rect 30932 9503 30984 9512
rect 30932 9469 30941 9503
rect 30941 9469 30975 9503
rect 30975 9469 30984 9503
rect 30932 9460 30984 9469
rect 32588 9460 32640 9512
rect 45008 9528 45060 9580
rect 48596 9528 48648 9580
rect 49424 9596 49476 9648
rect 49884 9596 49936 9648
rect 49148 9571 49200 9580
rect 49148 9537 49157 9571
rect 49157 9537 49191 9571
rect 49191 9537 49200 9571
rect 49148 9528 49200 9537
rect 49700 9528 49752 9580
rect 50252 9596 50304 9648
rect 51264 9596 51316 9648
rect 35716 9503 35768 9512
rect 27068 9435 27120 9444
rect 27068 9401 27077 9435
rect 27077 9401 27111 9435
rect 27111 9401 27120 9435
rect 27068 9392 27120 9401
rect 34428 9392 34480 9444
rect 35716 9469 35725 9503
rect 35725 9469 35759 9503
rect 35759 9469 35768 9503
rect 35716 9460 35768 9469
rect 40224 9503 40276 9512
rect 40224 9469 40233 9503
rect 40233 9469 40267 9503
rect 40267 9469 40276 9503
rect 40224 9460 40276 9469
rect 43628 9503 43680 9512
rect 43628 9469 43637 9503
rect 43637 9469 43671 9503
rect 43671 9469 43680 9503
rect 43628 9460 43680 9469
rect 46756 9460 46808 9512
rect 47584 9503 47636 9512
rect 47584 9469 47593 9503
rect 47593 9469 47627 9503
rect 47627 9469 47636 9503
rect 47584 9460 47636 9469
rect 49884 9460 49936 9512
rect 50804 9460 50856 9512
rect 50988 9503 51040 9512
rect 50988 9469 50997 9503
rect 50997 9469 51031 9503
rect 51031 9469 51040 9503
rect 50988 9460 51040 9469
rect 48412 9392 48464 9444
rect 29092 9324 29144 9376
rect 30380 9367 30432 9376
rect 30380 9333 30389 9367
rect 30389 9333 30423 9367
rect 30423 9333 30432 9367
rect 30380 9324 30432 9333
rect 36728 9367 36780 9376
rect 36728 9333 36737 9367
rect 36737 9333 36771 9367
rect 36771 9333 36780 9367
rect 36728 9324 36780 9333
rect 39212 9324 39264 9376
rect 40960 9324 41012 9376
rect 47768 9367 47820 9376
rect 47768 9333 47777 9367
rect 47777 9333 47811 9367
rect 47811 9333 47820 9367
rect 47768 9324 47820 9333
rect 48780 9324 48832 9376
rect 50252 9392 50304 9444
rect 50528 9392 50580 9444
rect 50712 9324 50764 9376
rect 50988 9324 51040 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 65654 9222 65706 9274
rect 65718 9222 65770 9274
rect 65782 9222 65834 9274
rect 65846 9222 65898 9274
rect 65910 9222 65962 9274
rect 15936 9120 15988 9172
rect 19340 9120 19392 9172
rect 21548 9163 21600 9172
rect 21548 9129 21557 9163
rect 21557 9129 21591 9163
rect 21591 9129 21600 9163
rect 21548 9120 21600 9129
rect 21916 9163 21968 9172
rect 21916 9129 21925 9163
rect 21925 9129 21959 9163
rect 21959 9129 21968 9163
rect 21916 9120 21968 9129
rect 28080 9120 28132 9172
rect 29644 9163 29696 9172
rect 8116 9052 8168 9104
rect 14096 9052 14148 9104
rect 16120 9052 16172 9104
rect 27068 9052 27120 9104
rect 9772 9027 9824 9036
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 9680 8916 9732 8968
rect 15384 8984 15436 9036
rect 16488 8984 16540 9036
rect 21824 8984 21876 9036
rect 25320 9027 25372 9036
rect 25320 8993 25329 9027
rect 25329 8993 25363 9027
rect 25363 8993 25372 9027
rect 25320 8984 25372 8993
rect 26240 8984 26292 9036
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 14924 8916 14976 8968
rect 9956 8891 10008 8900
rect 9956 8857 9965 8891
rect 9965 8857 9999 8891
rect 9999 8857 10008 8891
rect 9956 8848 10008 8857
rect 15476 8848 15528 8900
rect 16488 8848 16540 8900
rect 12256 8780 12308 8832
rect 15660 8780 15712 8832
rect 18236 8916 18288 8968
rect 20168 8916 20220 8968
rect 20628 8959 20680 8968
rect 20628 8925 20637 8959
rect 20637 8925 20671 8959
rect 20671 8925 20680 8959
rect 20628 8916 20680 8925
rect 25412 8916 25464 8968
rect 28448 8916 28500 8968
rect 29000 8959 29052 8968
rect 29000 8925 29009 8959
rect 29009 8925 29043 8959
rect 29043 8925 29052 8959
rect 29000 8916 29052 8925
rect 29644 9129 29653 9163
rect 29653 9129 29687 9163
rect 29687 9129 29696 9163
rect 29644 9120 29696 9129
rect 29736 9120 29788 9172
rect 32128 9120 32180 9172
rect 34612 9120 34664 9172
rect 36728 9120 36780 9172
rect 46940 9120 46992 9172
rect 48872 9163 48924 9172
rect 48872 9129 48881 9163
rect 48881 9129 48915 9163
rect 48915 9129 48924 9163
rect 48872 9120 48924 9129
rect 49332 9163 49384 9172
rect 49332 9129 49341 9163
rect 49341 9129 49375 9163
rect 49375 9129 49384 9163
rect 49332 9120 49384 9129
rect 50068 9120 50120 9172
rect 50896 9120 50948 9172
rect 35808 9052 35860 9104
rect 33048 8916 33100 8968
rect 33140 8916 33192 8968
rect 40316 8984 40368 9036
rect 49424 9052 49476 9104
rect 49700 9052 49752 9104
rect 50804 9052 50856 9104
rect 48964 9027 49016 9036
rect 48964 8993 48973 9027
rect 48973 8993 49007 9027
rect 49007 8993 49016 9027
rect 48964 8984 49016 8993
rect 44180 8959 44232 8968
rect 44180 8925 44189 8959
rect 44189 8925 44223 8959
rect 44223 8925 44232 8959
rect 44180 8916 44232 8925
rect 47952 8959 48004 8968
rect 47952 8925 47961 8959
rect 47961 8925 47995 8959
rect 47995 8925 48004 8959
rect 47952 8916 48004 8925
rect 48780 8959 48832 8968
rect 18236 8780 18288 8832
rect 20812 8823 20864 8832
rect 20812 8789 20821 8823
rect 20821 8789 20855 8823
rect 20855 8789 20864 8823
rect 20812 8780 20864 8789
rect 23480 8848 23532 8900
rect 27988 8848 28040 8900
rect 22100 8780 22152 8832
rect 30564 8848 30616 8900
rect 32312 8848 32364 8900
rect 32680 8891 32732 8900
rect 32680 8857 32689 8891
rect 32689 8857 32723 8891
rect 32723 8857 32732 8891
rect 32680 8848 32732 8857
rect 36452 8848 36504 8900
rect 36912 8891 36964 8900
rect 36912 8857 36921 8891
rect 36921 8857 36955 8891
rect 36955 8857 36964 8891
rect 36912 8848 36964 8857
rect 40500 8848 40552 8900
rect 40960 8848 41012 8900
rect 47768 8848 47820 8900
rect 48780 8925 48789 8959
rect 48789 8925 48823 8959
rect 48823 8925 48832 8959
rect 48780 8916 48832 8925
rect 49608 8916 49660 8968
rect 50528 8959 50580 8968
rect 50528 8925 50537 8959
rect 50537 8925 50571 8959
rect 50571 8925 50580 8959
rect 50528 8916 50580 8925
rect 50896 8916 50948 8968
rect 49516 8848 49568 8900
rect 50988 8848 51040 8900
rect 35440 8823 35492 8832
rect 35440 8789 35449 8823
rect 35449 8789 35483 8823
rect 35483 8789 35492 8823
rect 35440 8780 35492 8789
rect 41696 8823 41748 8832
rect 41696 8789 41705 8823
rect 41705 8789 41739 8823
rect 41739 8789 41748 8823
rect 41696 8780 41748 8789
rect 44272 8823 44324 8832
rect 44272 8789 44281 8823
rect 44281 8789 44315 8823
rect 44315 8789 44324 8823
rect 44272 8780 44324 8789
rect 48504 8780 48556 8832
rect 50712 8780 50764 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 6644 8576 6696 8628
rect 6828 8619 6880 8628
rect 6828 8585 6837 8619
rect 6837 8585 6871 8619
rect 6871 8585 6880 8619
rect 6828 8576 6880 8585
rect 9036 8576 9088 8628
rect 9772 8551 9824 8560
rect 9772 8517 9781 8551
rect 9781 8517 9815 8551
rect 9815 8517 9824 8551
rect 9772 8508 9824 8517
rect 7380 8372 7432 8424
rect 7932 8372 7984 8424
rect 9588 8372 9640 8424
rect 14096 8576 14148 8628
rect 21824 8619 21876 8628
rect 11980 8508 12032 8560
rect 12348 8483 12400 8492
rect 12348 8449 12357 8483
rect 12357 8449 12391 8483
rect 12391 8449 12400 8483
rect 12348 8440 12400 8449
rect 16120 8551 16172 8560
rect 16120 8517 16129 8551
rect 16129 8517 16163 8551
rect 16163 8517 16172 8551
rect 16120 8508 16172 8517
rect 14740 8440 14792 8492
rect 15384 8483 15436 8492
rect 15384 8449 15393 8483
rect 15393 8449 15427 8483
rect 15427 8449 15436 8483
rect 15384 8440 15436 8449
rect 16580 8440 16632 8492
rect 17868 8508 17920 8560
rect 20628 8508 20680 8560
rect 16948 8483 17000 8492
rect 16948 8449 16982 8483
rect 16982 8449 17000 8483
rect 16948 8440 17000 8449
rect 20168 8440 20220 8492
rect 21824 8585 21833 8619
rect 21833 8585 21867 8619
rect 21867 8585 21876 8619
rect 21824 8576 21876 8585
rect 25780 8619 25832 8628
rect 25780 8585 25789 8619
rect 25789 8585 25823 8619
rect 25823 8585 25832 8619
rect 25780 8576 25832 8585
rect 26332 8619 26384 8628
rect 26332 8585 26341 8619
rect 26341 8585 26375 8619
rect 26375 8585 26384 8619
rect 26332 8576 26384 8585
rect 27988 8576 28040 8628
rect 29000 8576 29052 8628
rect 29828 8576 29880 8628
rect 31208 8619 31260 8628
rect 31208 8585 31217 8619
rect 31217 8585 31251 8619
rect 31251 8585 31260 8619
rect 31208 8576 31260 8585
rect 31944 8576 31996 8628
rect 33048 8576 33100 8628
rect 36912 8576 36964 8628
rect 40224 8576 40276 8628
rect 40500 8576 40552 8628
rect 22100 8483 22152 8492
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 12716 8415 12768 8424
rect 12716 8381 12725 8415
rect 12725 8381 12759 8415
rect 12759 8381 12768 8415
rect 12716 8372 12768 8381
rect 15660 8372 15712 8424
rect 20444 8415 20496 8424
rect 20444 8381 20453 8415
rect 20453 8381 20487 8415
rect 20487 8381 20496 8415
rect 20444 8372 20496 8381
rect 20628 8372 20680 8424
rect 9680 8304 9732 8356
rect 10784 8304 10836 8356
rect 13728 8304 13780 8356
rect 18052 8347 18104 8356
rect 18052 8313 18061 8347
rect 18061 8313 18095 8347
rect 18095 8313 18104 8347
rect 18052 8304 18104 8313
rect 19248 8304 19300 8356
rect 22100 8449 22109 8483
rect 22109 8449 22143 8483
rect 22143 8449 22152 8483
rect 22100 8440 22152 8449
rect 22652 8483 22704 8492
rect 22652 8449 22661 8483
rect 22661 8449 22695 8483
rect 22695 8449 22704 8483
rect 22652 8440 22704 8449
rect 23296 8483 23348 8492
rect 23296 8449 23305 8483
rect 23305 8449 23339 8483
rect 23339 8449 23348 8483
rect 23296 8440 23348 8449
rect 23480 8483 23532 8492
rect 23480 8449 23489 8483
rect 23489 8449 23523 8483
rect 23523 8449 23532 8483
rect 23480 8440 23532 8449
rect 25320 8483 25372 8492
rect 25320 8449 25329 8483
rect 25329 8449 25363 8483
rect 25363 8449 25372 8483
rect 25320 8440 25372 8449
rect 32680 8508 32732 8560
rect 26332 8440 26384 8492
rect 28264 8440 28316 8492
rect 24952 8372 25004 8424
rect 25780 8372 25832 8424
rect 27252 8372 27304 8424
rect 29092 8440 29144 8492
rect 29644 8483 29696 8492
rect 29644 8449 29653 8483
rect 29653 8449 29687 8483
rect 29687 8449 29696 8483
rect 29644 8440 29696 8449
rect 32312 8483 32364 8492
rect 30932 8415 30984 8424
rect 24400 8304 24452 8356
rect 5356 8236 5408 8288
rect 21916 8236 21968 8288
rect 23020 8236 23072 8288
rect 25412 8279 25464 8288
rect 25412 8245 25421 8279
rect 25421 8245 25455 8279
rect 25455 8245 25464 8279
rect 25412 8236 25464 8245
rect 26424 8304 26476 8356
rect 28172 8304 28224 8356
rect 30932 8381 30941 8415
rect 30941 8381 30975 8415
rect 30975 8381 30984 8415
rect 30932 8372 30984 8381
rect 31300 8372 31352 8424
rect 32312 8449 32351 8483
rect 32351 8449 32364 8483
rect 32312 8440 32364 8449
rect 32496 8483 32548 8492
rect 32496 8449 32505 8483
rect 32505 8449 32539 8483
rect 32539 8449 32548 8483
rect 35440 8508 35492 8560
rect 32496 8440 32548 8449
rect 30656 8304 30708 8356
rect 33600 8372 33652 8424
rect 40040 8440 40092 8492
rect 41696 8508 41748 8560
rect 29552 8236 29604 8288
rect 32956 8279 33008 8288
rect 32956 8245 32965 8279
rect 32965 8245 32999 8279
rect 32999 8245 33008 8279
rect 32956 8236 33008 8245
rect 34244 8279 34296 8288
rect 34244 8245 34253 8279
rect 34253 8245 34287 8279
rect 34287 8245 34296 8279
rect 34244 8236 34296 8245
rect 34704 8236 34756 8288
rect 40224 8347 40276 8356
rect 40224 8313 40233 8347
rect 40233 8313 40267 8347
rect 40267 8313 40276 8347
rect 40224 8304 40276 8313
rect 35716 8236 35768 8288
rect 39580 8279 39632 8288
rect 39580 8245 39589 8279
rect 39589 8245 39623 8279
rect 39623 8245 39632 8279
rect 39580 8236 39632 8245
rect 40960 8372 41012 8424
rect 43260 8440 43312 8492
rect 43720 8576 43772 8628
rect 50160 8619 50212 8628
rect 44272 8508 44324 8560
rect 50160 8585 50169 8619
rect 50169 8585 50203 8619
rect 50203 8585 50212 8619
rect 50160 8576 50212 8585
rect 48872 8508 48924 8560
rect 49332 8508 49384 8560
rect 50896 8576 50948 8628
rect 50804 8508 50856 8560
rect 48320 8440 48372 8492
rect 48964 8440 49016 8492
rect 49424 8483 49476 8492
rect 49424 8449 49433 8483
rect 49433 8449 49467 8483
rect 49467 8449 49476 8483
rect 49424 8440 49476 8449
rect 49700 8440 49752 8492
rect 41788 8372 41840 8424
rect 41144 8347 41196 8356
rect 41144 8313 41153 8347
rect 41153 8313 41187 8347
rect 41187 8313 41196 8347
rect 41144 8304 41196 8313
rect 41236 8347 41288 8356
rect 41236 8313 41245 8347
rect 41245 8313 41279 8347
rect 41279 8313 41288 8347
rect 48596 8372 48648 8424
rect 41236 8304 41288 8313
rect 49608 8304 49660 8356
rect 48596 8279 48648 8288
rect 48596 8245 48605 8279
rect 48605 8245 48639 8279
rect 48639 8245 48648 8279
rect 48596 8236 48648 8245
rect 49332 8236 49384 8288
rect 49976 8236 50028 8288
rect 50620 8236 50672 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 65654 8134 65706 8186
rect 65718 8134 65770 8186
rect 65782 8134 65834 8186
rect 65846 8134 65898 8186
rect 65910 8134 65962 8186
rect 6644 8032 6696 8084
rect 8300 8032 8352 8084
rect 9588 8075 9640 8084
rect 9588 8041 9597 8075
rect 9597 8041 9631 8075
rect 9631 8041 9640 8075
rect 9588 8032 9640 8041
rect 9956 8032 10008 8084
rect 4712 7896 4764 7948
rect 5356 7871 5408 7880
rect 5356 7837 5390 7871
rect 5390 7837 5408 7871
rect 5356 7828 5408 7837
rect 9220 7828 9272 7880
rect 10968 8007 11020 8016
rect 10968 7973 10977 8007
rect 10977 7973 11011 8007
rect 11011 7973 11020 8007
rect 10968 7964 11020 7973
rect 13268 7964 13320 8016
rect 14832 8032 14884 8084
rect 13728 7896 13780 7948
rect 14648 7896 14700 7948
rect 11428 7828 11480 7880
rect 12624 7828 12676 7880
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 14924 7828 14976 7837
rect 10876 7760 10928 7812
rect 14740 7803 14792 7812
rect 14740 7769 14749 7803
rect 14749 7769 14783 7803
rect 14783 7769 14792 7803
rect 14740 7760 14792 7769
rect 16948 8032 17000 8084
rect 20168 8032 20220 8084
rect 20812 8032 20864 8084
rect 21824 8032 21876 8084
rect 22652 8032 22704 8084
rect 24676 8032 24728 8084
rect 25320 8075 25372 8084
rect 25320 8041 25329 8075
rect 25329 8041 25363 8075
rect 25363 8041 25372 8075
rect 25320 8032 25372 8041
rect 25780 8075 25832 8084
rect 25780 8041 25789 8075
rect 25789 8041 25823 8075
rect 25823 8041 25832 8075
rect 25780 8032 25832 8041
rect 28264 8032 28316 8084
rect 28632 8032 28684 8084
rect 29644 8075 29696 8084
rect 29644 8041 29653 8075
rect 29653 8041 29687 8075
rect 29687 8041 29696 8075
rect 29644 8032 29696 8041
rect 30564 8075 30616 8084
rect 30564 8041 30573 8075
rect 30573 8041 30607 8075
rect 30607 8041 30616 8075
rect 30564 8032 30616 8041
rect 20904 7964 20956 8016
rect 26240 7964 26292 8016
rect 26332 7964 26384 8016
rect 34244 8032 34296 8084
rect 34796 8032 34848 8084
rect 35348 8032 35400 8084
rect 35716 8075 35768 8084
rect 35716 8041 35725 8075
rect 35725 8041 35759 8075
rect 35759 8041 35768 8075
rect 35716 8032 35768 8041
rect 40224 8032 40276 8084
rect 31300 7964 31352 8016
rect 40960 8032 41012 8084
rect 41696 8075 41748 8084
rect 41696 8041 41705 8075
rect 41705 8041 41739 8075
rect 41739 8041 41748 8075
rect 41696 8032 41748 8041
rect 50160 8032 50212 8084
rect 17868 7896 17920 7948
rect 19156 7896 19208 7948
rect 19248 7871 19300 7880
rect 18236 7803 18288 7812
rect 18236 7769 18245 7803
rect 18245 7769 18279 7803
rect 18279 7769 18288 7803
rect 18236 7760 18288 7769
rect 19248 7837 19257 7871
rect 19257 7837 19291 7871
rect 19291 7837 19300 7871
rect 19248 7828 19300 7837
rect 22468 7896 22520 7948
rect 27344 7939 27396 7948
rect 27344 7905 27353 7939
rect 27353 7905 27387 7939
rect 27387 7905 27396 7939
rect 27344 7896 27396 7905
rect 32588 7939 32640 7948
rect 32588 7905 32597 7939
rect 32597 7905 32631 7939
rect 32631 7905 32640 7939
rect 32588 7896 32640 7905
rect 21916 7871 21968 7880
rect 21916 7837 21925 7871
rect 21925 7837 21959 7871
rect 21959 7837 21968 7871
rect 21916 7828 21968 7837
rect 22192 7828 22244 7880
rect 23388 7871 23440 7880
rect 19432 7760 19484 7812
rect 20168 7803 20220 7812
rect 20168 7769 20202 7803
rect 20202 7769 20220 7803
rect 20168 7760 20220 7769
rect 20444 7760 20496 7812
rect 22100 7803 22152 7812
rect 22100 7769 22109 7803
rect 22109 7769 22143 7803
rect 22143 7769 22152 7803
rect 22100 7760 22152 7769
rect 7840 7735 7892 7744
rect 7840 7701 7849 7735
rect 7849 7701 7883 7735
rect 7883 7701 7892 7735
rect 7840 7692 7892 7701
rect 15936 7735 15988 7744
rect 15936 7701 15945 7735
rect 15945 7701 15979 7735
rect 15979 7701 15988 7735
rect 15936 7692 15988 7701
rect 18052 7692 18104 7744
rect 21824 7692 21876 7744
rect 23388 7837 23397 7871
rect 23397 7837 23431 7871
rect 23431 7837 23440 7871
rect 23388 7828 23440 7837
rect 23480 7871 23532 7880
rect 23480 7837 23489 7871
rect 23489 7837 23523 7871
rect 23523 7837 23532 7871
rect 24400 7871 24452 7880
rect 23480 7828 23532 7837
rect 24400 7837 24409 7871
rect 24409 7837 24443 7871
rect 24443 7837 24452 7871
rect 24400 7828 24452 7837
rect 27436 7871 27488 7880
rect 27436 7837 27445 7871
rect 27445 7837 27479 7871
rect 27479 7837 27488 7871
rect 27436 7828 27488 7837
rect 30380 7871 30432 7880
rect 25780 7760 25832 7812
rect 28356 7803 28408 7812
rect 28356 7769 28365 7803
rect 28365 7769 28399 7803
rect 28399 7769 28408 7803
rect 28356 7760 28408 7769
rect 30380 7837 30389 7871
rect 30389 7837 30423 7871
rect 30423 7837 30432 7871
rect 30380 7828 30432 7837
rect 32956 7828 33008 7880
rect 33600 7871 33652 7880
rect 33600 7837 33609 7871
rect 33609 7837 33643 7871
rect 33643 7837 33652 7871
rect 33600 7828 33652 7837
rect 35440 7896 35492 7948
rect 26424 7692 26476 7744
rect 34796 7760 34848 7812
rect 35532 7828 35584 7880
rect 39212 7828 39264 7880
rect 40868 7964 40920 8016
rect 46940 7964 46992 8016
rect 54668 7964 54720 8016
rect 41144 7896 41196 7948
rect 41604 7871 41656 7880
rect 40040 7760 40092 7812
rect 32404 7692 32456 7744
rect 34428 7692 34480 7744
rect 40408 7760 40460 7812
rect 41604 7837 41613 7871
rect 41613 7837 41647 7871
rect 41647 7837 41656 7871
rect 41604 7828 41656 7837
rect 43260 7828 43312 7880
rect 49700 7896 49752 7948
rect 43076 7760 43128 7812
rect 45008 7828 45060 7880
rect 45560 7828 45612 7880
rect 48320 7871 48372 7880
rect 48320 7837 48329 7871
rect 48329 7837 48363 7871
rect 48363 7837 48372 7871
rect 48320 7828 48372 7837
rect 48596 7828 48648 7880
rect 49332 7828 49384 7880
rect 50712 7828 50764 7880
rect 49976 7760 50028 7812
rect 41236 7692 41288 7744
rect 43996 7692 44048 7744
rect 44088 7735 44140 7744
rect 44088 7701 44097 7735
rect 44097 7701 44131 7735
rect 44131 7701 44140 7735
rect 45100 7735 45152 7744
rect 44088 7692 44140 7701
rect 45100 7701 45109 7735
rect 45109 7701 45143 7735
rect 45143 7701 45152 7735
rect 45100 7692 45152 7701
rect 48596 7692 48648 7744
rect 49700 7692 49752 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 9220 7531 9272 7540
rect 7840 7420 7892 7472
rect 9220 7497 9229 7531
rect 9229 7497 9263 7531
rect 9263 7497 9272 7531
rect 9220 7488 9272 7497
rect 9312 7488 9364 7540
rect 10876 7488 10928 7540
rect 20352 7488 20404 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 21824 7488 21876 7540
rect 28264 7531 28316 7540
rect 11980 7463 12032 7472
rect 11980 7429 11989 7463
rect 11989 7429 12023 7463
rect 12023 7429 12032 7463
rect 11980 7420 12032 7429
rect 14740 7420 14792 7472
rect 18236 7420 18288 7472
rect 22192 7420 22244 7472
rect 22284 7463 22336 7472
rect 22284 7429 22293 7463
rect 22293 7429 22327 7463
rect 22327 7429 22336 7463
rect 23020 7463 23072 7472
rect 22284 7420 22336 7429
rect 23020 7429 23029 7463
rect 23029 7429 23063 7463
rect 23063 7429 23072 7463
rect 23020 7420 23072 7429
rect 28264 7497 28273 7531
rect 28273 7497 28307 7531
rect 28307 7497 28316 7531
rect 28264 7488 28316 7497
rect 28356 7488 28408 7540
rect 28816 7531 28868 7540
rect 28816 7497 28825 7531
rect 28825 7497 28859 7531
rect 28859 7497 28868 7531
rect 28816 7488 28868 7497
rect 31208 7488 31260 7540
rect 35532 7531 35584 7540
rect 35532 7497 35541 7531
rect 35541 7497 35575 7531
rect 35575 7497 35584 7531
rect 35532 7488 35584 7497
rect 41144 7488 41196 7540
rect 41604 7488 41656 7540
rect 41788 7531 41840 7540
rect 41788 7497 41797 7531
rect 41797 7497 41831 7531
rect 41831 7497 41840 7531
rect 41788 7488 41840 7497
rect 44088 7488 44140 7540
rect 52736 7488 52788 7540
rect 29184 7420 29236 7472
rect 29552 7420 29604 7472
rect 7196 7352 7248 7404
rect 7932 7352 7984 7404
rect 15476 7395 15528 7404
rect 5356 7284 5408 7336
rect 9312 7284 9364 7336
rect 15476 7361 15485 7395
rect 15485 7361 15519 7395
rect 15519 7361 15528 7395
rect 15476 7352 15528 7361
rect 19156 7352 19208 7404
rect 19340 7352 19392 7404
rect 19800 7352 19852 7404
rect 20996 7352 21048 7404
rect 24676 7352 24728 7404
rect 25228 7395 25280 7404
rect 25228 7361 25237 7395
rect 25237 7361 25271 7395
rect 25271 7361 25280 7395
rect 25228 7352 25280 7361
rect 27712 7395 27764 7404
rect 27712 7361 27721 7395
rect 27721 7361 27755 7395
rect 27755 7361 27764 7395
rect 27712 7352 27764 7361
rect 30656 7352 30708 7404
rect 32404 7395 32456 7404
rect 32404 7361 32413 7395
rect 32413 7361 32447 7395
rect 32447 7361 32456 7395
rect 32404 7352 32456 7361
rect 34428 7395 34480 7404
rect 34428 7361 34437 7395
rect 34437 7361 34471 7395
rect 34471 7361 34480 7395
rect 34428 7352 34480 7361
rect 34704 7395 34756 7404
rect 34704 7361 34713 7395
rect 34713 7361 34747 7395
rect 34747 7361 34756 7395
rect 34704 7352 34756 7361
rect 35348 7395 35400 7404
rect 35348 7361 35357 7395
rect 35357 7361 35391 7395
rect 35391 7361 35400 7395
rect 35348 7352 35400 7361
rect 39580 7420 39632 7472
rect 40316 7420 40368 7472
rect 43996 7463 44048 7472
rect 38016 7395 38068 7404
rect 38016 7361 38025 7395
rect 38025 7361 38059 7395
rect 38059 7361 38068 7395
rect 38016 7352 38068 7361
rect 40868 7352 40920 7404
rect 10508 7216 10560 7268
rect 12624 7216 12676 7268
rect 6368 7191 6420 7200
rect 6368 7157 6377 7191
rect 6377 7157 6411 7191
rect 6411 7157 6420 7191
rect 6368 7148 6420 7157
rect 11980 7148 12032 7200
rect 14464 7284 14516 7336
rect 14648 7284 14700 7336
rect 15384 7327 15436 7336
rect 15384 7293 15393 7327
rect 15393 7293 15427 7327
rect 15427 7293 15436 7327
rect 16672 7327 16724 7336
rect 15384 7284 15436 7293
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 20260 7284 20312 7336
rect 22100 7284 22152 7336
rect 22468 7284 22520 7336
rect 24768 7327 24820 7336
rect 24768 7293 24777 7327
rect 24777 7293 24811 7327
rect 24811 7293 24820 7327
rect 24768 7284 24820 7293
rect 28632 7284 28684 7336
rect 32128 7327 32180 7336
rect 32128 7293 32137 7327
rect 32137 7293 32171 7327
rect 32171 7293 32180 7327
rect 32128 7284 32180 7293
rect 35440 7284 35492 7336
rect 40224 7327 40276 7336
rect 40224 7293 40233 7327
rect 40233 7293 40267 7327
rect 40267 7293 40276 7327
rect 40224 7284 40276 7293
rect 14096 7216 14148 7268
rect 16764 7216 16816 7268
rect 26240 7259 26292 7268
rect 26240 7225 26249 7259
rect 26249 7225 26283 7259
rect 26283 7225 26292 7259
rect 41052 7352 41104 7404
rect 41236 7352 41288 7404
rect 41788 7395 41840 7404
rect 41788 7361 41797 7395
rect 41797 7361 41831 7395
rect 41831 7361 41840 7395
rect 41788 7352 41840 7361
rect 43996 7429 44005 7463
rect 44005 7429 44039 7463
rect 44039 7429 44048 7463
rect 43996 7420 44048 7429
rect 43076 7395 43128 7404
rect 43076 7361 43085 7395
rect 43085 7361 43119 7395
rect 43119 7361 43128 7395
rect 43076 7352 43128 7361
rect 43260 7395 43312 7404
rect 43260 7361 43269 7395
rect 43269 7361 43303 7395
rect 43303 7361 43312 7395
rect 43260 7352 43312 7361
rect 45100 7352 45152 7404
rect 48504 7395 48556 7404
rect 48504 7361 48513 7395
rect 48513 7361 48547 7395
rect 48547 7361 48556 7395
rect 48504 7352 48556 7361
rect 49792 7352 49844 7404
rect 49976 7395 50028 7404
rect 49976 7361 49985 7395
rect 49985 7361 50019 7395
rect 50019 7361 50028 7395
rect 49976 7352 50028 7361
rect 43720 7327 43772 7336
rect 43720 7293 43729 7327
rect 43729 7293 43763 7327
rect 43763 7293 43772 7327
rect 43720 7284 43772 7293
rect 26240 7216 26292 7225
rect 41236 7216 41288 7268
rect 13912 7191 13964 7200
rect 13912 7157 13921 7191
rect 13921 7157 13955 7191
rect 13955 7157 13964 7191
rect 13912 7148 13964 7157
rect 33324 7148 33376 7200
rect 37464 7191 37516 7200
rect 37464 7157 37473 7191
rect 37473 7157 37507 7191
rect 37507 7157 37516 7191
rect 37464 7148 37516 7157
rect 40132 7148 40184 7200
rect 43996 7148 44048 7200
rect 44456 7148 44508 7200
rect 47860 7191 47912 7200
rect 47860 7157 47869 7191
rect 47869 7157 47903 7191
rect 47903 7157 47912 7191
rect 47860 7148 47912 7157
rect 48320 7191 48372 7200
rect 48320 7157 48329 7191
rect 48329 7157 48363 7191
rect 48363 7157 48372 7191
rect 48320 7148 48372 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 65654 7046 65706 7098
rect 65718 7046 65770 7098
rect 65782 7046 65834 7098
rect 65846 7046 65898 7098
rect 65910 7046 65962 7098
rect 7196 6987 7248 6996
rect 7196 6953 7205 6987
rect 7205 6953 7239 6987
rect 7239 6953 7248 6987
rect 7196 6944 7248 6953
rect 22192 6944 22244 6996
rect 16672 6876 16724 6928
rect 23848 6944 23900 6996
rect 26424 6944 26476 6996
rect 27160 6944 27212 6996
rect 27252 6944 27304 6996
rect 27436 6944 27488 6996
rect 34796 6987 34848 6996
rect 34796 6953 34805 6987
rect 34805 6953 34839 6987
rect 34839 6953 34848 6987
rect 34796 6944 34848 6953
rect 37464 6944 37516 6996
rect 4712 6808 4764 6860
rect 5356 6851 5408 6860
rect 5356 6817 5365 6851
rect 5365 6817 5399 6851
rect 5399 6817 5408 6851
rect 5356 6808 5408 6817
rect 7932 6808 7984 6860
rect 10416 6808 10468 6860
rect 13084 6808 13136 6860
rect 16580 6808 16632 6860
rect 17592 6808 17644 6860
rect 20628 6851 20680 6860
rect 6368 6740 6420 6792
rect 8392 6740 8444 6792
rect 10968 6740 11020 6792
rect 12348 6740 12400 6792
rect 13912 6740 13964 6792
rect 16396 6740 16448 6792
rect 9312 6672 9364 6724
rect 14004 6672 14056 6724
rect 14464 6672 14516 6724
rect 15200 6672 15252 6724
rect 16764 6740 16816 6792
rect 18052 6740 18104 6792
rect 20628 6817 20637 6851
rect 20637 6817 20671 6851
rect 20671 6817 20680 6851
rect 20628 6808 20680 6817
rect 20260 6783 20312 6792
rect 20260 6749 20269 6783
rect 20269 6749 20303 6783
rect 20303 6749 20312 6783
rect 20260 6740 20312 6749
rect 21180 6740 21232 6792
rect 22192 6783 22244 6792
rect 22192 6749 22201 6783
rect 22201 6749 22235 6783
rect 22235 6749 22244 6783
rect 22192 6740 22244 6749
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 10048 6647 10100 6656
rect 7656 6604 7708 6613
rect 10048 6613 10057 6647
rect 10057 6613 10091 6647
rect 10091 6613 10100 6647
rect 10048 6604 10100 6613
rect 10324 6604 10376 6656
rect 12072 6604 12124 6656
rect 12808 6647 12860 6656
rect 12808 6613 12817 6647
rect 12817 6613 12851 6647
rect 12851 6613 12860 6647
rect 12808 6604 12860 6613
rect 13636 6604 13688 6656
rect 15476 6604 15528 6656
rect 19340 6672 19392 6724
rect 23204 6740 23256 6792
rect 24032 6740 24084 6792
rect 23572 6715 23624 6724
rect 19432 6647 19484 6656
rect 19432 6613 19441 6647
rect 19441 6613 19475 6647
rect 19475 6613 19484 6647
rect 19432 6604 19484 6613
rect 23020 6647 23072 6656
rect 23020 6613 23029 6647
rect 23029 6613 23063 6647
rect 23063 6613 23072 6647
rect 23020 6604 23072 6613
rect 23572 6681 23581 6715
rect 23581 6681 23615 6715
rect 23615 6681 23624 6715
rect 23572 6672 23624 6681
rect 23388 6604 23440 6656
rect 23940 6604 23992 6656
rect 27344 6808 27396 6860
rect 29644 6876 29696 6928
rect 32128 6876 32180 6928
rect 32772 6876 32824 6928
rect 39948 6876 40000 6928
rect 40040 6876 40092 6928
rect 40224 6944 40276 6996
rect 40500 6944 40552 6996
rect 45192 6944 45244 6996
rect 45560 6876 45612 6928
rect 28632 6808 28684 6860
rect 35624 6808 35676 6860
rect 41144 6808 41196 6860
rect 45008 6808 45060 6860
rect 25228 6783 25280 6792
rect 25228 6749 25237 6783
rect 25237 6749 25271 6783
rect 25271 6749 25280 6783
rect 25228 6740 25280 6749
rect 26424 6783 26476 6792
rect 26424 6749 26433 6783
rect 26433 6749 26467 6783
rect 26467 6749 26476 6783
rect 26424 6740 26476 6749
rect 29276 6740 29328 6792
rect 29644 6740 29696 6792
rect 34796 6740 34848 6792
rect 35348 6740 35400 6792
rect 40500 6740 40552 6792
rect 41880 6740 41932 6792
rect 43996 6783 44048 6792
rect 43996 6749 44005 6783
rect 44005 6749 44039 6783
rect 44039 6749 44048 6783
rect 43996 6740 44048 6749
rect 44272 6740 44324 6792
rect 27160 6672 27212 6724
rect 28724 6672 28776 6724
rect 30656 6672 30708 6724
rect 24952 6604 25004 6656
rect 25228 6604 25280 6656
rect 26056 6647 26108 6656
rect 26056 6613 26065 6647
rect 26065 6613 26099 6647
rect 26099 6613 26108 6647
rect 26056 6604 26108 6613
rect 27252 6647 27304 6656
rect 27252 6613 27261 6647
rect 27261 6613 27295 6647
rect 27295 6613 27304 6647
rect 27252 6604 27304 6613
rect 30288 6604 30340 6656
rect 31116 6604 31168 6656
rect 40684 6672 40736 6724
rect 45192 6783 45244 6792
rect 45192 6749 45201 6783
rect 45201 6749 45235 6783
rect 45235 6749 45244 6783
rect 45192 6740 45244 6749
rect 47492 6672 47544 6724
rect 48412 6808 48464 6860
rect 48596 6808 48648 6860
rect 49976 6876 50028 6928
rect 48320 6740 48372 6792
rect 49424 6740 49476 6792
rect 43352 6647 43404 6656
rect 43352 6613 43361 6647
rect 43361 6613 43395 6647
rect 43395 6613 43404 6647
rect 43352 6604 43404 6613
rect 44180 6604 44232 6656
rect 45744 6647 45796 6656
rect 45744 6613 45753 6647
rect 45753 6613 45787 6647
rect 45787 6613 45796 6647
rect 45744 6604 45796 6613
rect 48504 6604 48556 6656
rect 49700 6672 49752 6724
rect 49976 6604 50028 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 8300 6400 8352 6452
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 10508 6400 10560 6452
rect 10968 6443 11020 6452
rect 10968 6409 10977 6443
rect 10977 6409 11011 6443
rect 11011 6409 11020 6443
rect 10968 6400 11020 6409
rect 12348 6400 12400 6452
rect 14740 6443 14792 6452
rect 14740 6409 14749 6443
rect 14749 6409 14783 6443
rect 14783 6409 14792 6443
rect 14740 6400 14792 6409
rect 17408 6400 17460 6452
rect 17592 6400 17644 6452
rect 18052 6443 18104 6452
rect 18052 6409 18061 6443
rect 18061 6409 18095 6443
rect 18095 6409 18104 6443
rect 18052 6400 18104 6409
rect 19432 6400 19484 6452
rect 7656 6332 7708 6384
rect 11428 6332 11480 6384
rect 11520 6332 11572 6384
rect 10048 6264 10100 6316
rect 6460 6196 6512 6248
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 11612 6264 11664 6316
rect 14004 6332 14056 6384
rect 13636 6307 13688 6316
rect 13636 6273 13670 6307
rect 13670 6273 13688 6307
rect 13636 6264 13688 6273
rect 15200 6307 15252 6316
rect 15200 6273 15209 6307
rect 15209 6273 15243 6307
rect 15243 6273 15252 6307
rect 15200 6264 15252 6273
rect 19800 6332 19852 6384
rect 20996 6375 21048 6384
rect 20996 6341 21005 6375
rect 21005 6341 21039 6375
rect 21039 6341 21048 6375
rect 20996 6332 21048 6341
rect 17960 6264 18012 6316
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 19156 6264 19208 6316
rect 23020 6332 23072 6384
rect 27344 6332 27396 6384
rect 23572 6264 23624 6316
rect 25228 6264 25280 6316
rect 27988 6400 28040 6452
rect 29644 6443 29696 6452
rect 29644 6409 29653 6443
rect 29653 6409 29687 6443
rect 29687 6409 29696 6443
rect 29644 6400 29696 6409
rect 32128 6400 32180 6452
rect 34796 6443 34848 6452
rect 34796 6409 34805 6443
rect 34805 6409 34839 6443
rect 34839 6409 34848 6443
rect 34796 6400 34848 6409
rect 41880 6443 41932 6452
rect 41880 6409 41889 6443
rect 41889 6409 41923 6443
rect 41923 6409 41932 6443
rect 41880 6400 41932 6409
rect 43352 6400 43404 6452
rect 44272 6400 44324 6452
rect 27528 6332 27580 6384
rect 28448 6332 28500 6384
rect 33324 6375 33376 6384
rect 27712 6264 27764 6316
rect 28724 6264 28776 6316
rect 29276 6307 29328 6316
rect 29276 6273 29285 6307
rect 29285 6273 29319 6307
rect 29319 6273 29328 6307
rect 33324 6341 33333 6375
rect 33333 6341 33367 6375
rect 33367 6341 33376 6375
rect 33324 6332 33376 6341
rect 33876 6332 33928 6384
rect 44180 6375 44232 6384
rect 44180 6341 44189 6375
rect 44189 6341 44223 6375
rect 44223 6341 44232 6375
rect 44180 6332 44232 6341
rect 45744 6332 45796 6384
rect 50068 6332 50120 6384
rect 29276 6264 29328 6273
rect 30288 6264 30340 6316
rect 31760 6264 31812 6316
rect 32588 6264 32640 6316
rect 38660 6264 38712 6316
rect 40960 6307 41012 6316
rect 40960 6273 40987 6307
rect 40987 6273 41012 6307
rect 41236 6307 41288 6316
rect 40960 6264 41012 6273
rect 41236 6273 41245 6307
rect 41245 6273 41279 6307
rect 41279 6273 41288 6307
rect 41236 6264 41288 6273
rect 48320 6307 48372 6316
rect 48320 6273 48329 6307
rect 48329 6273 48363 6307
rect 48363 6273 48372 6307
rect 48320 6264 48372 6273
rect 48964 6264 49016 6316
rect 49884 6307 49936 6316
rect 49884 6273 49893 6307
rect 49893 6273 49927 6307
rect 49927 6273 49936 6307
rect 49884 6264 49936 6273
rect 11060 6196 11112 6248
rect 11520 6239 11572 6248
rect 11520 6205 11529 6239
rect 11529 6205 11563 6239
rect 11563 6205 11572 6239
rect 11520 6196 11572 6205
rect 16764 6196 16816 6248
rect 17408 6239 17460 6248
rect 17408 6205 17417 6239
rect 17417 6205 17451 6239
rect 17451 6205 17460 6239
rect 17408 6196 17460 6205
rect 22192 6196 22244 6248
rect 23204 6196 23256 6248
rect 6920 6103 6972 6112
rect 6920 6069 6929 6103
rect 6929 6069 6963 6103
rect 6963 6069 6972 6103
rect 6920 6060 6972 6069
rect 9496 6060 9548 6112
rect 12164 6060 12216 6112
rect 16580 6060 16632 6112
rect 19340 6060 19392 6112
rect 27344 6196 27396 6248
rect 26424 6128 26476 6180
rect 27620 6196 27672 6248
rect 28816 6196 28868 6248
rect 26240 6060 26292 6112
rect 27620 6060 27672 6112
rect 27988 6103 28040 6112
rect 27988 6069 27997 6103
rect 27997 6069 28031 6103
rect 28031 6069 28040 6103
rect 27988 6060 28040 6069
rect 40040 6239 40092 6248
rect 40040 6205 40049 6239
rect 40049 6205 40083 6239
rect 40083 6205 40092 6239
rect 40040 6196 40092 6205
rect 40224 6239 40276 6248
rect 40224 6205 40233 6239
rect 40233 6205 40267 6239
rect 40267 6205 40276 6239
rect 40224 6196 40276 6205
rect 40316 6196 40368 6248
rect 43720 6196 43772 6248
rect 47124 6196 47176 6248
rect 48596 6239 48648 6248
rect 48596 6205 48605 6239
rect 48605 6205 48639 6239
rect 48639 6205 48648 6239
rect 51448 6307 51500 6316
rect 51448 6273 51457 6307
rect 51457 6273 51491 6307
rect 51491 6273 51500 6307
rect 51448 6264 51500 6273
rect 48596 6196 48648 6205
rect 54024 6196 54076 6248
rect 30380 6060 30432 6112
rect 37372 6103 37424 6112
rect 37372 6069 37381 6103
rect 37381 6069 37415 6103
rect 37415 6069 37424 6103
rect 37372 6060 37424 6069
rect 41788 6060 41840 6112
rect 46940 6060 46992 6112
rect 50068 6060 50120 6112
rect 50988 6128 51040 6180
rect 50896 6060 50948 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 65654 5958 65706 6010
rect 65718 5958 65770 6010
rect 65782 5958 65834 6010
rect 65846 5958 65898 6010
rect 65910 5958 65962 6010
rect 7656 5856 7708 5908
rect 8300 5788 8352 5840
rect 5356 5720 5408 5772
rect 11520 5856 11572 5908
rect 11612 5856 11664 5908
rect 11428 5831 11480 5840
rect 11428 5797 11437 5831
rect 11437 5797 11471 5831
rect 11471 5797 11480 5831
rect 11428 5788 11480 5797
rect 11060 5720 11112 5772
rect 18604 5720 18656 5772
rect 9128 5652 9180 5704
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 10324 5695 10376 5704
rect 10324 5661 10358 5695
rect 10358 5661 10376 5695
rect 10324 5652 10376 5661
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 12440 5652 12492 5704
rect 13268 5652 13320 5704
rect 14096 5695 14148 5704
rect 14096 5661 14105 5695
rect 14105 5661 14139 5695
rect 14139 5661 14148 5695
rect 14096 5652 14148 5661
rect 6368 5584 6420 5636
rect 12808 5584 12860 5636
rect 15384 5652 15436 5704
rect 17592 5652 17644 5704
rect 18144 5652 18196 5704
rect 18696 5695 18748 5704
rect 18696 5661 18705 5695
rect 18705 5661 18739 5695
rect 18739 5661 18748 5695
rect 18696 5652 18748 5661
rect 15292 5584 15344 5636
rect 15936 5584 15988 5636
rect 26240 5856 26292 5908
rect 27712 5856 27764 5908
rect 28724 5899 28776 5908
rect 28724 5865 28733 5899
rect 28733 5865 28767 5899
rect 28767 5865 28776 5899
rect 28724 5856 28776 5865
rect 31116 5856 31168 5908
rect 32772 5899 32824 5908
rect 32772 5865 32781 5899
rect 32781 5865 32815 5899
rect 32815 5865 32824 5899
rect 32772 5856 32824 5865
rect 33876 5899 33928 5908
rect 33876 5865 33885 5899
rect 33885 5865 33919 5899
rect 33919 5865 33928 5899
rect 33876 5856 33928 5865
rect 20536 5788 20588 5840
rect 20628 5788 20680 5840
rect 19800 5763 19852 5772
rect 19800 5729 19809 5763
rect 19809 5729 19843 5763
rect 19843 5729 19852 5763
rect 19800 5720 19852 5729
rect 19984 5763 20036 5772
rect 19984 5729 19993 5763
rect 19993 5729 20027 5763
rect 20027 5729 20036 5763
rect 19984 5720 20036 5729
rect 20444 5652 20496 5704
rect 24952 5788 25004 5840
rect 23112 5763 23164 5772
rect 23112 5729 23121 5763
rect 23121 5729 23155 5763
rect 23155 5729 23164 5763
rect 23112 5720 23164 5729
rect 24124 5652 24176 5704
rect 26056 5652 26108 5704
rect 9404 5516 9456 5568
rect 12900 5559 12952 5568
rect 12900 5525 12909 5559
rect 12909 5525 12943 5559
rect 12943 5525 12952 5559
rect 12900 5516 12952 5525
rect 14004 5516 14056 5568
rect 14096 5516 14148 5568
rect 14556 5516 14608 5568
rect 20628 5584 20680 5636
rect 23940 5584 23992 5636
rect 30380 5788 30432 5840
rect 26424 5695 26476 5704
rect 26424 5661 26433 5695
rect 26433 5661 26467 5695
rect 26467 5661 26476 5695
rect 26424 5652 26476 5661
rect 27528 5652 27580 5704
rect 19432 5516 19484 5568
rect 22560 5559 22612 5568
rect 22560 5525 22569 5559
rect 22569 5525 22603 5559
rect 22603 5525 22612 5559
rect 22560 5516 22612 5525
rect 31760 5720 31812 5772
rect 33784 5695 33836 5704
rect 33784 5661 33793 5695
rect 33793 5661 33827 5695
rect 33827 5661 33836 5695
rect 37464 5856 37516 5908
rect 46296 5856 46348 5908
rect 48964 5856 49016 5908
rect 51448 5856 51500 5908
rect 35808 5720 35860 5772
rect 38384 5763 38436 5772
rect 38384 5729 38393 5763
rect 38393 5729 38427 5763
rect 38427 5729 38436 5763
rect 38384 5720 38436 5729
rect 40132 5720 40184 5772
rect 41144 5763 41196 5772
rect 41144 5729 41153 5763
rect 41153 5729 41187 5763
rect 41187 5729 41196 5763
rect 41144 5720 41196 5729
rect 48596 5763 48648 5772
rect 48596 5729 48605 5763
rect 48605 5729 48639 5763
rect 48639 5729 48648 5763
rect 48596 5720 48648 5729
rect 50068 5720 50120 5772
rect 33784 5652 33836 5661
rect 37372 5652 37424 5704
rect 39304 5695 39356 5704
rect 39304 5661 39313 5695
rect 39313 5661 39347 5695
rect 39347 5661 39356 5695
rect 39304 5652 39356 5661
rect 40408 5695 40460 5704
rect 40408 5661 40417 5695
rect 40417 5661 40451 5695
rect 40451 5661 40460 5695
rect 40408 5652 40460 5661
rect 46480 5652 46532 5704
rect 48412 5652 48464 5704
rect 50896 5695 50948 5704
rect 32680 5584 32732 5636
rect 35900 5584 35952 5636
rect 39856 5584 39908 5636
rect 50896 5661 50905 5695
rect 50905 5661 50939 5695
rect 50939 5661 50948 5695
rect 50896 5652 50948 5661
rect 50988 5652 51040 5704
rect 30656 5516 30708 5568
rect 37280 5559 37332 5568
rect 37280 5525 37289 5559
rect 37289 5525 37323 5559
rect 37323 5525 37332 5559
rect 37280 5516 37332 5525
rect 37372 5516 37424 5568
rect 38108 5559 38160 5568
rect 38108 5525 38117 5559
rect 38117 5525 38151 5559
rect 38151 5525 38160 5559
rect 38108 5516 38160 5525
rect 38844 5516 38896 5568
rect 39764 5516 39816 5568
rect 46572 5516 46624 5568
rect 48412 5516 48464 5568
rect 55220 5584 55272 5636
rect 61384 5584 61436 5636
rect 49884 5516 49936 5568
rect 50160 5559 50212 5568
rect 50160 5525 50169 5559
rect 50169 5525 50203 5559
rect 50203 5525 50212 5559
rect 50160 5516 50212 5525
rect 51356 5516 51408 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 6368 5355 6420 5364
rect 6368 5321 6377 5355
rect 6377 5321 6411 5355
rect 6411 5321 6420 5355
rect 6368 5312 6420 5321
rect 10508 5355 10560 5364
rect 10508 5321 10517 5355
rect 10517 5321 10551 5355
rect 10551 5321 10560 5355
rect 10508 5312 10560 5321
rect 20444 5355 20496 5364
rect 6920 5176 6972 5228
rect 9128 5219 9180 5228
rect 9128 5185 9137 5219
rect 9137 5185 9171 5219
rect 9171 5185 9180 5219
rect 9128 5176 9180 5185
rect 9404 5219 9456 5228
rect 9404 5185 9438 5219
rect 9438 5185 9456 5219
rect 9404 5176 9456 5185
rect 9864 5176 9916 5228
rect 13176 5176 13228 5228
rect 14924 5176 14976 5228
rect 17960 5244 18012 5296
rect 20444 5321 20453 5355
rect 20453 5321 20487 5355
rect 20487 5321 20496 5355
rect 20444 5312 20496 5321
rect 20536 5312 20588 5364
rect 28632 5312 28684 5364
rect 31116 5355 31168 5364
rect 31116 5321 31125 5355
rect 31125 5321 31159 5355
rect 31159 5321 31168 5355
rect 31116 5312 31168 5321
rect 32680 5312 32732 5364
rect 35900 5312 35952 5364
rect 37280 5312 37332 5364
rect 19432 5244 19484 5296
rect 26332 5244 26384 5296
rect 40040 5312 40092 5364
rect 41328 5312 41380 5364
rect 48136 5312 48188 5364
rect 42432 5244 42484 5296
rect 49516 5244 49568 5296
rect 15752 5219 15804 5228
rect 15752 5185 15761 5219
rect 15761 5185 15795 5219
rect 15795 5185 15804 5219
rect 15752 5176 15804 5185
rect 22560 5176 22612 5228
rect 12072 5108 12124 5160
rect 13360 5108 13412 5160
rect 15936 5108 15988 5160
rect 17868 5108 17920 5160
rect 10416 5040 10468 5092
rect 12440 5040 12492 5092
rect 15016 5040 15068 5092
rect 12348 4972 12400 5024
rect 12624 5015 12676 5024
rect 12624 4981 12633 5015
rect 12633 4981 12667 5015
rect 12667 4981 12676 5015
rect 12624 4972 12676 4981
rect 13820 4972 13872 5024
rect 16028 5040 16080 5092
rect 15844 5015 15896 5024
rect 15844 4981 15853 5015
rect 15853 4981 15887 5015
rect 15887 4981 15896 5015
rect 15844 4972 15896 4981
rect 17776 4972 17828 5024
rect 18420 4972 18472 5024
rect 18604 4972 18656 5024
rect 23112 5108 23164 5160
rect 25412 5176 25464 5228
rect 25780 5176 25832 5228
rect 27528 5219 27580 5228
rect 27528 5185 27537 5219
rect 27537 5185 27571 5219
rect 27571 5185 27580 5219
rect 27528 5176 27580 5185
rect 27804 5219 27856 5228
rect 27804 5185 27838 5219
rect 27838 5185 27856 5219
rect 27804 5176 27856 5185
rect 33784 5176 33836 5228
rect 38108 5176 38160 5228
rect 38660 5219 38712 5228
rect 38660 5185 38669 5219
rect 38669 5185 38703 5219
rect 38703 5185 38712 5219
rect 38660 5176 38712 5185
rect 38844 5176 38896 5228
rect 39948 5219 40000 5228
rect 39948 5185 39957 5219
rect 39957 5185 39991 5219
rect 39991 5185 40000 5219
rect 39948 5176 40000 5185
rect 42800 5176 42852 5228
rect 38384 5108 38436 5160
rect 22744 4972 22796 5024
rect 23756 4972 23808 5024
rect 24584 4972 24636 5024
rect 30656 5015 30708 5024
rect 30656 4981 30665 5015
rect 30665 4981 30699 5015
rect 30699 4981 30708 5015
rect 30656 4972 30708 4981
rect 37188 4972 37240 5024
rect 41328 5151 41380 5160
rect 41328 5117 41337 5151
rect 41337 5117 41371 5151
rect 41371 5117 41380 5151
rect 41328 5108 41380 5117
rect 43352 5108 43404 5160
rect 49884 5176 49936 5228
rect 50068 5219 50120 5228
rect 50068 5185 50077 5219
rect 50077 5185 50111 5219
rect 50111 5185 50120 5219
rect 50068 5176 50120 5185
rect 50620 5176 50672 5228
rect 46296 5108 46348 5160
rect 40132 5040 40184 5092
rect 40316 5083 40368 5092
rect 40316 5049 40325 5083
rect 40325 5049 40359 5083
rect 40359 5049 40368 5083
rect 40316 5040 40368 5049
rect 46848 5040 46900 5092
rect 47308 5040 47360 5092
rect 48688 5040 48740 5092
rect 41788 4972 41840 5024
rect 45652 4972 45704 5024
rect 45928 4972 45980 5024
rect 46756 4972 46808 5024
rect 49056 5015 49108 5024
rect 49056 4981 49065 5015
rect 49065 4981 49099 5015
rect 49099 4981 49108 5015
rect 49056 4972 49108 4981
rect 51724 4972 51776 5024
rect 53288 4972 53340 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 65654 4870 65706 4922
rect 65718 4870 65770 4922
rect 65782 4870 65834 4922
rect 65846 4870 65898 4922
rect 65910 4870 65962 4922
rect 12716 4768 12768 4820
rect 14372 4768 14424 4820
rect 15660 4768 15712 4820
rect 9864 4743 9916 4752
rect 9864 4709 9873 4743
rect 9873 4709 9907 4743
rect 9907 4709 9916 4743
rect 9864 4700 9916 4709
rect 10416 4743 10468 4752
rect 10416 4709 10425 4743
rect 10425 4709 10459 4743
rect 10459 4709 10468 4743
rect 10416 4700 10468 4709
rect 14188 4700 14240 4752
rect 15752 4700 15804 4752
rect 13268 4632 13320 4684
rect 15660 4632 15712 4684
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 12716 4607 12768 4616
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 13452 4564 13504 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 18972 4700 19024 4752
rect 20260 4768 20312 4820
rect 24124 4768 24176 4820
rect 27804 4768 27856 4820
rect 40224 4768 40276 4820
rect 40960 4768 41012 4820
rect 48136 4768 48188 4820
rect 54024 4811 54076 4820
rect 54024 4777 54033 4811
rect 54033 4777 54067 4811
rect 54067 4777 54076 4811
rect 54024 4768 54076 4777
rect 54576 4811 54628 4820
rect 54576 4777 54585 4811
rect 54585 4777 54619 4811
rect 54619 4777 54628 4811
rect 54576 4768 54628 4777
rect 55312 4811 55364 4820
rect 55312 4777 55321 4811
rect 55321 4777 55355 4811
rect 55355 4777 55364 4811
rect 55312 4768 55364 4777
rect 22008 4700 22060 4752
rect 38108 4700 38160 4752
rect 41236 4700 41288 4752
rect 47216 4700 47268 4752
rect 49976 4700 50028 4752
rect 16028 4632 16080 4684
rect 16672 4632 16724 4684
rect 17868 4632 17920 4684
rect 22468 4675 22520 4684
rect 22468 4641 22477 4675
rect 22477 4641 22511 4675
rect 22511 4641 22520 4675
rect 22468 4632 22520 4641
rect 38936 4632 38988 4684
rect 41144 4632 41196 4684
rect 41328 4632 41380 4684
rect 44824 4632 44876 4684
rect 46204 4632 46256 4684
rect 47676 4632 47728 4684
rect 51172 4632 51224 4684
rect 16212 4607 16264 4616
rect 11612 4496 11664 4548
rect 16212 4573 16221 4607
rect 16221 4573 16255 4607
rect 16255 4573 16264 4607
rect 16212 4564 16264 4573
rect 16856 4607 16908 4616
rect 14832 4496 14884 4548
rect 15108 4539 15160 4548
rect 15108 4505 15117 4539
rect 15117 4505 15151 4539
rect 15151 4505 15160 4539
rect 15108 4496 15160 4505
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 19340 4564 19392 4616
rect 21088 4564 21140 4616
rect 22744 4607 22796 4616
rect 22744 4573 22778 4607
rect 22778 4573 22796 4607
rect 22744 4564 22796 4573
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 27988 4564 28040 4616
rect 29920 4564 29972 4616
rect 31116 4607 31168 4616
rect 31116 4573 31125 4607
rect 31125 4573 31159 4607
rect 31159 4573 31168 4607
rect 31116 4564 31168 4573
rect 31852 4564 31904 4616
rect 35808 4607 35860 4616
rect 35808 4573 35817 4607
rect 35817 4573 35851 4607
rect 35851 4573 35860 4607
rect 35808 4564 35860 4573
rect 37188 4564 37240 4616
rect 38752 4564 38804 4616
rect 16948 4496 17000 4548
rect 19248 4496 19300 4548
rect 36084 4539 36136 4548
rect 36084 4505 36093 4539
rect 36093 4505 36127 4539
rect 36127 4505 36136 4539
rect 36084 4496 36136 4505
rect 12256 4471 12308 4480
rect 12256 4437 12265 4471
rect 12265 4437 12299 4471
rect 12299 4437 12308 4471
rect 12256 4428 12308 4437
rect 15476 4428 15528 4480
rect 20996 4428 21048 4480
rect 24952 4428 25004 4480
rect 32956 4428 33008 4480
rect 42800 4564 42852 4616
rect 42984 4607 43036 4616
rect 42984 4573 42993 4607
rect 42993 4573 43027 4607
rect 43027 4573 43036 4607
rect 42984 4564 43036 4573
rect 43352 4564 43404 4616
rect 44272 4607 44324 4616
rect 44272 4573 44281 4607
rect 44281 4573 44315 4607
rect 44315 4573 44324 4607
rect 44272 4564 44324 4573
rect 45100 4564 45152 4616
rect 45376 4564 45428 4616
rect 46940 4607 46992 4616
rect 46940 4573 46949 4607
rect 46949 4573 46983 4607
rect 46983 4573 46992 4607
rect 46940 4564 46992 4573
rect 48044 4564 48096 4616
rect 48320 4564 48372 4616
rect 50896 4564 50948 4616
rect 40868 4539 40920 4548
rect 40868 4505 40877 4539
rect 40877 4505 40911 4539
rect 40911 4505 40920 4539
rect 40868 4496 40920 4505
rect 42524 4496 42576 4548
rect 42616 4496 42668 4548
rect 39856 4471 39908 4480
rect 39856 4437 39865 4471
rect 39865 4437 39899 4471
rect 39899 4437 39908 4471
rect 39856 4428 39908 4437
rect 42340 4428 42392 4480
rect 42800 4471 42852 4480
rect 42800 4437 42809 4471
rect 42809 4437 42843 4471
rect 42843 4437 42852 4471
rect 42800 4428 42852 4437
rect 43536 4471 43588 4480
rect 43536 4437 43545 4471
rect 43545 4437 43579 4471
rect 43579 4437 43588 4471
rect 43536 4428 43588 4437
rect 44180 4471 44232 4480
rect 44180 4437 44189 4471
rect 44189 4437 44223 4471
rect 44223 4437 44232 4471
rect 44180 4428 44232 4437
rect 45008 4471 45060 4480
rect 45008 4437 45017 4471
rect 45017 4437 45051 4471
rect 45051 4437 45060 4471
rect 45008 4428 45060 4437
rect 47032 4428 47084 4480
rect 48412 4471 48464 4480
rect 48412 4437 48421 4471
rect 48421 4437 48455 4471
rect 48455 4437 48464 4471
rect 48412 4428 48464 4437
rect 50712 4496 50764 4548
rect 51632 4471 51684 4480
rect 51632 4437 51641 4471
rect 51641 4437 51675 4471
rect 51675 4437 51684 4471
rect 51632 4428 51684 4437
rect 52092 4471 52144 4480
rect 52092 4437 52101 4471
rect 52101 4437 52135 4471
rect 52135 4437 52144 4471
rect 52092 4428 52144 4437
rect 55956 4471 56008 4480
rect 55956 4437 55965 4471
rect 55965 4437 55999 4471
rect 55999 4437 56008 4471
rect 55956 4428 56008 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 12072 4224 12124 4276
rect 8668 4131 8720 4140
rect 8668 4097 8677 4131
rect 8677 4097 8711 4131
rect 8711 4097 8720 4131
rect 8668 4088 8720 4097
rect 14280 4224 14332 4276
rect 15844 4267 15896 4276
rect 15844 4233 15853 4267
rect 15853 4233 15887 4267
rect 15887 4233 15896 4267
rect 15844 4224 15896 4233
rect 16856 4224 16908 4276
rect 20260 4224 20312 4276
rect 26332 4224 26384 4276
rect 33048 4267 33100 4276
rect 33048 4233 33057 4267
rect 33057 4233 33091 4267
rect 33091 4233 33100 4267
rect 33048 4224 33100 4233
rect 36084 4224 36136 4276
rect 42616 4224 42668 4276
rect 46388 4267 46440 4276
rect 46388 4233 46397 4267
rect 46397 4233 46431 4267
rect 46431 4233 46440 4267
rect 46388 4224 46440 4233
rect 48412 4224 48464 4276
rect 49516 4267 49568 4276
rect 49516 4233 49525 4267
rect 49525 4233 49559 4267
rect 49559 4233 49568 4267
rect 49516 4224 49568 4233
rect 50896 4224 50948 4276
rect 54024 4224 54076 4276
rect 67180 4224 67232 4276
rect 13728 4156 13780 4208
rect 14648 4199 14700 4208
rect 14648 4165 14657 4199
rect 14657 4165 14691 4199
rect 14691 4165 14700 4199
rect 14648 4156 14700 4165
rect 15384 4156 15436 4208
rect 12808 4088 12860 4140
rect 13544 4088 13596 4140
rect 15292 4088 15344 4140
rect 15476 4131 15528 4140
rect 15476 4097 15485 4131
rect 15485 4097 15519 4131
rect 15519 4097 15528 4131
rect 15476 4088 15528 4097
rect 15752 4131 15804 4140
rect 15752 4097 15761 4131
rect 15761 4097 15795 4131
rect 15795 4097 15804 4131
rect 15752 4088 15804 4097
rect 16212 4156 16264 4208
rect 16488 4088 16540 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 25044 4156 25096 4208
rect 12808 3952 12860 4004
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 16856 4020 16908 4072
rect 17960 4131 18012 4140
rect 17960 4097 17969 4131
rect 17969 4097 18003 4131
rect 18003 4097 18012 4131
rect 17960 4088 18012 4097
rect 18236 4088 18288 4140
rect 18604 4131 18656 4140
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 18604 4088 18656 4097
rect 19984 4088 20036 4140
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 23756 4131 23808 4140
rect 23756 4097 23765 4131
rect 23765 4097 23799 4131
rect 23799 4097 23808 4131
rect 23756 4088 23808 4097
rect 24952 4131 25004 4140
rect 24952 4097 24986 4131
rect 24986 4097 25004 4131
rect 24952 4088 25004 4097
rect 38844 4156 38896 4208
rect 42248 4156 42300 4208
rect 44180 4156 44232 4208
rect 45008 4156 45060 4208
rect 13452 3952 13504 4004
rect 14372 3952 14424 4004
rect 14924 3952 14976 4004
rect 16948 3952 17000 4004
rect 19892 4020 19944 4072
rect 31760 4088 31812 4140
rect 19156 3995 19208 4004
rect 19156 3961 19165 3995
rect 19165 3961 19199 3995
rect 19199 3961 19208 3995
rect 19156 3952 19208 3961
rect 14556 3884 14608 3936
rect 14740 3927 14792 3936
rect 14740 3893 14749 3927
rect 14749 3893 14783 3927
rect 14783 3893 14792 3927
rect 14740 3884 14792 3893
rect 14832 3884 14884 3936
rect 15568 3884 15620 3936
rect 15752 3884 15804 3936
rect 16764 3884 16816 3936
rect 20536 3884 20588 3936
rect 21732 3884 21784 3936
rect 23020 3884 23072 3936
rect 23940 3927 23992 3936
rect 23940 3893 23949 3927
rect 23949 3893 23983 3927
rect 23983 3893 23992 3927
rect 23940 3884 23992 3893
rect 24400 3884 24452 3936
rect 32128 4020 32180 4072
rect 32956 4020 33008 4072
rect 37372 4088 37424 4140
rect 37464 4131 37516 4140
rect 37464 4097 37473 4131
rect 37473 4097 37507 4131
rect 37507 4097 37516 4131
rect 37464 4088 37516 4097
rect 39856 4088 39908 4140
rect 40592 4088 40644 4140
rect 42432 4131 42484 4140
rect 42432 4097 42441 4131
rect 42441 4097 42475 4131
rect 42475 4097 42484 4131
rect 42432 4088 42484 4097
rect 45836 4088 45888 4140
rect 46572 4131 46624 4140
rect 37924 4020 37976 4072
rect 41788 4063 41840 4072
rect 41788 4029 41797 4063
rect 41797 4029 41831 4063
rect 41831 4029 41840 4063
rect 41788 4020 41840 4029
rect 45192 4063 45244 4072
rect 45192 4029 45201 4063
rect 45201 4029 45235 4063
rect 45235 4029 45244 4063
rect 45192 4020 45244 4029
rect 46296 4020 46348 4072
rect 46572 4097 46581 4131
rect 46581 4097 46615 4131
rect 46615 4097 46624 4131
rect 46572 4088 46624 4097
rect 48228 4088 48280 4140
rect 48596 4088 48648 4140
rect 49056 4088 49108 4140
rect 49332 4088 49384 4140
rect 49700 4020 49752 4072
rect 54668 4131 54720 4140
rect 54668 4097 54677 4131
rect 54677 4097 54711 4131
rect 54711 4097 54720 4131
rect 54668 4088 54720 4097
rect 55220 4131 55272 4140
rect 55220 4097 55229 4131
rect 55229 4097 55263 4131
rect 55263 4097 55272 4131
rect 55772 4131 55824 4140
rect 55220 4088 55272 4097
rect 55772 4097 55781 4131
rect 55781 4097 55815 4131
rect 55815 4097 55824 4131
rect 55772 4088 55824 4097
rect 56324 4131 56376 4140
rect 56324 4097 56333 4131
rect 56333 4097 56367 4131
rect 56367 4097 56376 4131
rect 56324 4088 56376 4097
rect 67364 4131 67416 4140
rect 67364 4097 67373 4131
rect 67373 4097 67407 4131
rect 67407 4097 67416 4131
rect 67364 4088 67416 4097
rect 50620 4063 50672 4072
rect 50620 4029 50629 4063
rect 50629 4029 50663 4063
rect 50663 4029 50672 4063
rect 50620 4020 50672 4029
rect 26424 3952 26476 4004
rect 39028 3952 39080 4004
rect 39856 3995 39908 4004
rect 39856 3961 39865 3995
rect 39865 3961 39899 3995
rect 39899 3961 39908 3995
rect 39856 3952 39908 3961
rect 40408 3952 40460 4004
rect 42432 3952 42484 4004
rect 27712 3884 27764 3936
rect 29000 3927 29052 3936
rect 29000 3893 29009 3927
rect 29009 3893 29043 3927
rect 29043 3893 29052 3927
rect 29000 3884 29052 3893
rect 29552 3927 29604 3936
rect 29552 3893 29561 3927
rect 29561 3893 29595 3927
rect 29595 3893 29604 3927
rect 29552 3884 29604 3893
rect 29644 3884 29696 3936
rect 31484 3884 31536 3936
rect 32220 3884 32272 3936
rect 37372 3927 37424 3936
rect 37372 3893 37381 3927
rect 37381 3893 37415 3927
rect 37415 3893 37424 3927
rect 37372 3884 37424 3893
rect 37648 3884 37700 3936
rect 38476 3884 38528 3936
rect 40592 3884 40644 3936
rect 41788 3884 41840 3936
rect 43444 3927 43496 3936
rect 43444 3893 43453 3927
rect 43453 3893 43487 3927
rect 43487 3893 43496 3927
rect 43444 3884 43496 3893
rect 46112 3952 46164 4004
rect 46940 3952 46992 4004
rect 50068 3952 50120 4004
rect 50160 3952 50212 4004
rect 50804 3952 50856 4004
rect 45560 3884 45612 3936
rect 46664 3884 46716 3936
rect 46848 3884 46900 3936
rect 47124 3884 47176 3936
rect 48228 3927 48280 3936
rect 48228 3893 48237 3927
rect 48237 3893 48271 3927
rect 48271 3893 48280 3927
rect 48228 3884 48280 3893
rect 49332 3884 49384 3936
rect 50252 3927 50304 3936
rect 50252 3893 50261 3927
rect 50261 3893 50295 3927
rect 50295 3893 50304 3927
rect 50252 3884 50304 3893
rect 50344 3884 50396 3936
rect 51264 3884 51316 3936
rect 51908 3884 51960 3936
rect 67548 3927 67600 3936
rect 67548 3893 67557 3927
rect 67557 3893 67591 3927
rect 67591 3893 67600 3927
rect 67548 3884 67600 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 65654 3782 65706 3834
rect 65718 3782 65770 3834
rect 65782 3782 65834 3834
rect 65846 3782 65898 3834
rect 65910 3782 65962 3834
rect 11612 3723 11664 3732
rect 11612 3689 11621 3723
rect 11621 3689 11655 3723
rect 11655 3689 11664 3723
rect 11612 3680 11664 3689
rect 12164 3680 12216 3732
rect 12808 3680 12860 3732
rect 13452 3680 13504 3732
rect 14188 3723 14240 3732
rect 14188 3689 14197 3723
rect 14197 3689 14231 3723
rect 14231 3689 14240 3723
rect 14188 3680 14240 3689
rect 14280 3680 14332 3732
rect 14924 3680 14976 3732
rect 15292 3680 15344 3732
rect 15752 3680 15804 3732
rect 16488 3723 16540 3732
rect 16488 3689 16497 3723
rect 16497 3689 16531 3723
rect 16531 3689 16540 3723
rect 16488 3680 16540 3689
rect 17500 3680 17552 3732
rect 20260 3723 20312 3732
rect 20260 3689 20269 3723
rect 20269 3689 20303 3723
rect 20303 3689 20312 3723
rect 20260 3680 20312 3689
rect 25780 3723 25832 3732
rect 25780 3689 25789 3723
rect 25789 3689 25823 3723
rect 25823 3689 25832 3723
rect 25780 3680 25832 3689
rect 31576 3680 31628 3732
rect 32588 3680 32640 3732
rect 33048 3680 33100 3732
rect 39580 3680 39632 3732
rect 42984 3680 43036 3732
rect 43812 3680 43864 3732
rect 20628 3612 20680 3664
rect 8116 3476 8168 3528
rect 11612 3544 11664 3596
rect 14004 3544 14056 3596
rect 14280 3544 14332 3596
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 8392 3451 8444 3460
rect 8392 3417 8401 3451
rect 8401 3417 8435 3451
rect 8435 3417 8444 3451
rect 8392 3408 8444 3417
rect 11888 3476 11940 3528
rect 12072 3519 12124 3528
rect 12072 3485 12081 3519
rect 12081 3485 12115 3519
rect 12115 3485 12124 3519
rect 12072 3476 12124 3485
rect 12900 3476 12952 3528
rect 13360 3476 13412 3528
rect 13636 3476 13688 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 15384 3476 15436 3528
rect 16488 3544 16540 3596
rect 19340 3544 19392 3596
rect 20536 3587 20588 3596
rect 20536 3553 20545 3587
rect 20545 3553 20579 3587
rect 20579 3553 20588 3587
rect 20536 3544 20588 3553
rect 24400 3587 24452 3596
rect 24400 3553 24409 3587
rect 24409 3553 24443 3587
rect 24443 3553 24452 3587
rect 24400 3544 24452 3553
rect 26424 3544 26476 3596
rect 29092 3544 29144 3596
rect 32312 3544 32364 3596
rect 35808 3544 35860 3596
rect 42616 3612 42668 3664
rect 45100 3680 45152 3732
rect 47768 3680 47820 3732
rect 48596 3723 48648 3732
rect 48596 3689 48605 3723
rect 48605 3689 48639 3723
rect 48639 3689 48648 3723
rect 48596 3680 48648 3689
rect 20076 3476 20128 3528
rect 21088 3476 21140 3528
rect 22008 3476 22060 3528
rect 22468 3476 22520 3528
rect 23572 3476 23624 3528
rect 9956 3340 10008 3392
rect 10692 3408 10744 3460
rect 11336 3408 11388 3460
rect 12256 3340 12308 3392
rect 12624 3340 12676 3392
rect 16120 3340 16172 3392
rect 16488 3451 16540 3460
rect 16488 3417 16497 3451
rect 16497 3417 16531 3451
rect 16531 3417 16540 3451
rect 16488 3408 16540 3417
rect 23940 3476 23992 3528
rect 26056 3476 26108 3528
rect 27436 3476 27488 3528
rect 28264 3476 28316 3528
rect 28816 3476 28868 3528
rect 29460 3476 29512 3528
rect 33232 3476 33284 3528
rect 37372 3476 37424 3528
rect 38568 3476 38620 3528
rect 39028 3476 39080 3528
rect 39856 3519 39908 3528
rect 39856 3485 39865 3519
rect 39865 3485 39899 3519
rect 39899 3485 39908 3519
rect 39856 3476 39908 3485
rect 41972 3544 42024 3596
rect 42432 3544 42484 3596
rect 42524 3544 42576 3596
rect 43444 3544 43496 3596
rect 42800 3476 42852 3528
rect 24400 3408 24452 3460
rect 31024 3451 31076 3460
rect 31024 3417 31033 3451
rect 31033 3417 31067 3451
rect 31067 3417 31076 3451
rect 31024 3408 31076 3417
rect 31484 3408 31536 3460
rect 18236 3340 18288 3392
rect 39028 3383 39080 3392
rect 39028 3349 39037 3383
rect 39037 3349 39071 3383
rect 39071 3349 39080 3383
rect 39028 3340 39080 3349
rect 40592 3408 40644 3460
rect 44548 3544 44600 3596
rect 46020 3612 46072 3664
rect 45560 3544 45612 3596
rect 46388 3544 46440 3596
rect 47124 3587 47176 3596
rect 47124 3553 47133 3587
rect 47133 3553 47167 3587
rect 47167 3553 47176 3587
rect 47124 3544 47176 3553
rect 47952 3544 48004 3596
rect 50344 3680 50396 3732
rect 48780 3612 48832 3664
rect 51816 3680 51868 3732
rect 67364 3723 67416 3732
rect 67364 3689 67373 3723
rect 67373 3689 67407 3723
rect 67407 3689 67416 3723
rect 67364 3680 67416 3689
rect 57244 3612 57296 3664
rect 48872 3544 48924 3596
rect 47032 3519 47084 3528
rect 47032 3485 47041 3519
rect 47041 3485 47075 3519
rect 47075 3485 47084 3519
rect 47032 3476 47084 3485
rect 47400 3476 47452 3528
rect 49056 3544 49108 3596
rect 49240 3544 49292 3596
rect 49792 3476 49844 3528
rect 50804 3476 50856 3528
rect 51724 3587 51776 3596
rect 51724 3553 51733 3587
rect 51733 3553 51767 3587
rect 51767 3553 51776 3587
rect 51724 3544 51776 3553
rect 54484 3544 54536 3596
rect 55864 3544 55916 3596
rect 57612 3544 57664 3596
rect 41144 3340 41196 3392
rect 46388 3408 46440 3460
rect 48044 3408 48096 3460
rect 41604 3383 41656 3392
rect 41604 3349 41613 3383
rect 41613 3349 41647 3383
rect 41647 3349 41656 3383
rect 42340 3383 42392 3392
rect 41604 3340 41656 3349
rect 42340 3349 42349 3383
rect 42349 3349 42383 3383
rect 42383 3349 42392 3383
rect 42340 3340 42392 3349
rect 42524 3340 42576 3392
rect 42708 3340 42760 3392
rect 43444 3340 43496 3392
rect 45284 3340 45336 3392
rect 48780 3340 48832 3392
rect 51264 3408 51316 3460
rect 52092 3476 52144 3528
rect 52368 3476 52420 3528
rect 54576 3476 54628 3528
rect 55404 3476 55456 3528
rect 56416 3476 56468 3528
rect 67180 3519 67232 3528
rect 67180 3485 67189 3519
rect 67189 3485 67223 3519
rect 67223 3485 67232 3519
rect 67180 3476 67232 3485
rect 53472 3451 53524 3460
rect 53472 3417 53481 3451
rect 53481 3417 53515 3451
rect 53515 3417 53524 3451
rect 53472 3408 53524 3417
rect 53932 3340 53984 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 10232 3136 10284 3188
rect 8484 3111 8536 3120
rect 8484 3077 8493 3111
rect 8493 3077 8527 3111
rect 8527 3077 8536 3111
rect 8484 3068 8536 3077
rect 12716 3179 12768 3188
rect 12716 3145 12725 3179
rect 12725 3145 12759 3179
rect 12759 3145 12768 3179
rect 12716 3136 12768 3145
rect 15108 3136 15160 3188
rect 15568 3136 15620 3188
rect 16488 3136 16540 3188
rect 19984 3179 20036 3188
rect 19984 3145 19993 3179
rect 19993 3145 20027 3179
rect 20027 3145 20036 3179
rect 19984 3136 20036 3145
rect 21088 3179 21140 3188
rect 21088 3145 21097 3179
rect 21097 3145 21131 3179
rect 21131 3145 21140 3179
rect 21088 3136 21140 3145
rect 29552 3136 29604 3188
rect 10140 3043 10192 3052
rect 10140 3009 10149 3043
rect 10149 3009 10183 3043
rect 10183 3009 10192 3043
rect 10140 3000 10192 3009
rect 10232 3000 10284 3052
rect 13360 3000 13412 3052
rect 10968 2932 11020 2984
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 12256 2932 12308 2984
rect 13912 3000 13964 3052
rect 14096 2975 14148 2984
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 15200 3068 15252 3120
rect 19064 3068 19116 3120
rect 29644 3068 29696 3120
rect 31024 3136 31076 3188
rect 32128 3179 32180 3188
rect 32128 3145 32137 3179
rect 32137 3145 32171 3179
rect 32171 3145 32180 3179
rect 32128 3136 32180 3145
rect 32588 3179 32640 3188
rect 32588 3145 32597 3179
rect 32597 3145 32631 3179
rect 32631 3145 32640 3179
rect 32588 3136 32640 3145
rect 38844 3136 38896 3188
rect 39856 3136 39908 3188
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 14740 3000 14792 3052
rect 19800 3043 19852 3052
rect 19800 3009 19809 3043
rect 19809 3009 19843 3043
rect 19843 3009 19852 3043
rect 19800 3000 19852 3009
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 29092 3043 29144 3052
rect 29092 3009 29101 3043
rect 29101 3009 29135 3043
rect 29135 3009 29144 3043
rect 29092 3000 29144 3009
rect 32220 3000 32272 3052
rect 39028 3068 39080 3120
rect 39764 3111 39816 3120
rect 39764 3077 39773 3111
rect 39773 3077 39807 3111
rect 39807 3077 39816 3111
rect 39764 3068 39816 3077
rect 43720 3136 43772 3188
rect 45192 3136 45244 3188
rect 41144 3068 41196 3120
rect 42064 3068 42116 3120
rect 42708 3068 42760 3120
rect 43536 3068 43588 3120
rect 15384 2975 15436 2984
rect 15384 2941 15393 2975
rect 15393 2941 15427 2975
rect 15427 2941 15436 2975
rect 15384 2932 15436 2941
rect 15476 2932 15528 2984
rect 20904 2932 20956 2984
rect 23848 2932 23900 2984
rect 25780 2932 25832 2984
rect 29368 2932 29420 2984
rect 32772 2975 32824 2984
rect 32772 2941 32781 2975
rect 32781 2941 32815 2975
rect 32815 2941 32824 2975
rect 32772 2932 32824 2941
rect 32956 2932 33008 2984
rect 10876 2796 10928 2848
rect 14464 2864 14516 2916
rect 15200 2864 15252 2916
rect 17316 2864 17368 2916
rect 19432 2864 19484 2916
rect 19800 2864 19852 2916
rect 21272 2864 21324 2916
rect 13084 2796 13136 2848
rect 14096 2796 14148 2848
rect 14188 2839 14240 2848
rect 14188 2805 14197 2839
rect 14197 2805 14231 2839
rect 14231 2805 14240 2839
rect 14188 2796 14240 2805
rect 15292 2796 15344 2848
rect 15568 2839 15620 2848
rect 15568 2805 15577 2839
rect 15577 2805 15611 2839
rect 15611 2805 15620 2839
rect 15568 2796 15620 2805
rect 20352 2796 20404 2848
rect 21456 2796 21508 2848
rect 23296 2796 23348 2848
rect 24952 2864 25004 2916
rect 28540 2864 28592 2916
rect 38200 2864 38252 2916
rect 41512 3043 41564 3052
rect 41512 3009 41521 3043
rect 41521 3009 41555 3043
rect 41555 3009 41564 3043
rect 41512 3000 41564 3009
rect 41880 3000 41932 3052
rect 48596 3136 48648 3188
rect 49700 3179 49752 3188
rect 48412 3068 48464 3120
rect 49240 3068 49292 3120
rect 49700 3145 49709 3179
rect 49709 3145 49743 3179
rect 49743 3145 49752 3179
rect 49700 3136 49752 3145
rect 38568 2932 38620 2984
rect 25504 2796 25556 2848
rect 26332 2796 26384 2848
rect 26884 2796 26936 2848
rect 30472 2796 30524 2848
rect 33784 2839 33836 2848
rect 33784 2805 33793 2839
rect 33793 2805 33827 2839
rect 33827 2805 33836 2839
rect 33784 2796 33836 2805
rect 34336 2796 34388 2848
rect 34796 2796 34848 2848
rect 35440 2796 35492 2848
rect 36268 2796 36320 2848
rect 36820 2796 36872 2848
rect 38660 2864 38712 2916
rect 41972 2932 42024 2984
rect 42340 2932 42392 2984
rect 44272 2932 44324 2984
rect 48228 2932 48280 2984
rect 49332 3000 49384 3052
rect 49608 3068 49660 3120
rect 50712 3136 50764 3188
rect 50068 3068 50120 3120
rect 51816 3043 51868 3052
rect 51816 3009 51825 3043
rect 51825 3009 51859 3043
rect 51859 3009 51868 3043
rect 51816 3000 51868 3009
rect 52736 3043 52788 3052
rect 52736 3009 52745 3043
rect 52745 3009 52779 3043
rect 52779 3009 52788 3043
rect 52736 3000 52788 3009
rect 54668 3068 54720 3120
rect 54760 3068 54812 3120
rect 56784 3068 56836 3120
rect 55128 3000 55180 3052
rect 55312 3000 55364 3052
rect 41052 2864 41104 2916
rect 43168 2864 43220 2916
rect 42248 2796 42300 2848
rect 42524 2796 42576 2848
rect 42800 2796 42852 2848
rect 43536 2839 43588 2848
rect 43536 2805 43545 2839
rect 43545 2805 43579 2839
rect 43579 2805 43588 2839
rect 43536 2796 43588 2805
rect 45284 2864 45336 2916
rect 47584 2907 47636 2916
rect 47584 2873 47593 2907
rect 47593 2873 47627 2907
rect 47627 2873 47636 2907
rect 47584 2864 47636 2873
rect 51724 2932 51776 2984
rect 56968 2932 57020 2984
rect 46020 2796 46072 2848
rect 49516 2839 49568 2848
rect 49516 2805 49525 2839
rect 49525 2805 49559 2839
rect 49559 2805 49568 2839
rect 49516 2796 49568 2805
rect 50620 2864 50672 2916
rect 51172 2864 51224 2916
rect 52828 2864 52880 2916
rect 54208 2864 54260 2916
rect 55128 2864 55180 2916
rect 57520 2864 57572 2916
rect 51080 2839 51132 2848
rect 51080 2805 51089 2839
rect 51089 2805 51123 2839
rect 51123 2805 51132 2839
rect 51080 2796 51132 2805
rect 51448 2796 51500 2848
rect 52276 2796 52328 2848
rect 53380 2796 53432 2848
rect 55588 2796 55640 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 65654 2694 65706 2746
rect 65718 2694 65770 2746
rect 65782 2694 65834 2746
rect 65846 2694 65898 2746
rect 65910 2694 65962 2746
rect 10968 2592 11020 2644
rect 11336 2524 11388 2576
rect 12348 2524 12400 2576
rect 12532 2524 12584 2576
rect 12440 2456 12492 2508
rect 12716 2499 12768 2508
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 10968 2431 11020 2440
rect 10968 2397 10977 2431
rect 10977 2397 11011 2431
rect 11011 2397 11020 2431
rect 10968 2388 11020 2397
rect 12716 2465 12725 2499
rect 12725 2465 12759 2499
rect 12759 2465 12768 2499
rect 12716 2456 12768 2465
rect 14648 2592 14700 2644
rect 16028 2635 16080 2644
rect 16028 2601 16037 2635
rect 16037 2601 16071 2635
rect 16071 2601 16080 2635
rect 16028 2592 16080 2601
rect 16764 2635 16816 2644
rect 16764 2601 16773 2635
rect 16773 2601 16807 2635
rect 16807 2601 16816 2635
rect 16764 2592 16816 2601
rect 19800 2592 19852 2644
rect 20260 2592 20312 2644
rect 32772 2592 32824 2644
rect 15108 2567 15160 2576
rect 15108 2533 15117 2567
rect 15117 2533 15151 2567
rect 15151 2533 15160 2567
rect 15108 2524 15160 2533
rect 17500 2567 17552 2576
rect 17500 2533 17509 2567
rect 17509 2533 17543 2567
rect 17543 2533 17552 2567
rect 17500 2524 17552 2533
rect 21180 2524 21232 2576
rect 24124 2524 24176 2576
rect 27160 2524 27212 2576
rect 30196 2524 30248 2576
rect 32404 2524 32456 2576
rect 33508 2524 33560 2576
rect 15292 2456 15344 2508
rect 22192 2456 22244 2508
rect 24676 2456 24728 2508
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 11704 2320 11756 2372
rect 11980 2320 12032 2372
rect 14740 2252 14792 2304
rect 15384 2320 15436 2372
rect 15844 2252 15896 2304
rect 16396 2320 16448 2372
rect 22744 2388 22796 2440
rect 25228 2388 25280 2440
rect 27988 2456 28040 2508
rect 30748 2456 30800 2508
rect 32680 2456 32732 2508
rect 21640 2320 21692 2372
rect 31300 2388 31352 2440
rect 32956 2388 33008 2440
rect 34060 2388 34112 2440
rect 34612 2388 34664 2440
rect 35164 2388 35216 2440
rect 35716 2388 35768 2440
rect 26608 2320 26660 2372
rect 30656 2320 30708 2372
rect 56784 2635 56836 2644
rect 56784 2601 56793 2635
rect 56793 2601 56827 2635
rect 56827 2601 56836 2635
rect 56784 2592 56836 2601
rect 40408 2524 40460 2576
rect 41604 2524 41656 2576
rect 44272 2524 44324 2576
rect 37096 2456 37148 2508
rect 39948 2456 40000 2508
rect 35992 2388 36044 2440
rect 36544 2388 36596 2440
rect 37372 2388 37424 2440
rect 40224 2431 40276 2440
rect 40224 2397 40233 2431
rect 40233 2397 40267 2431
rect 40267 2397 40276 2431
rect 40224 2388 40276 2397
rect 40960 2431 41012 2440
rect 40960 2397 40969 2431
rect 40969 2397 41003 2431
rect 41003 2397 41012 2431
rect 40960 2388 41012 2397
rect 42800 2456 42852 2508
rect 42892 2456 42944 2508
rect 46296 2524 46348 2576
rect 46664 2524 46716 2576
rect 52552 2524 52604 2576
rect 56692 2524 56744 2576
rect 47492 2456 47544 2508
rect 49884 2456 49936 2508
rect 51080 2456 51132 2508
rect 42156 2388 42208 2440
rect 42524 2388 42576 2440
rect 43904 2431 43956 2440
rect 43904 2397 43913 2431
rect 43913 2397 43947 2431
rect 43947 2397 43956 2431
rect 43904 2388 43956 2397
rect 21548 2252 21600 2304
rect 39856 2252 39908 2304
rect 40132 2252 40184 2304
rect 40868 2252 40920 2304
rect 42800 2320 42852 2372
rect 48596 2388 48648 2440
rect 46664 2363 46716 2372
rect 42708 2252 42760 2304
rect 45008 2252 45060 2304
rect 46664 2329 46673 2363
rect 46673 2329 46707 2363
rect 46707 2329 46716 2363
rect 46664 2320 46716 2329
rect 47860 2320 47912 2372
rect 48228 2320 48280 2372
rect 48964 2388 49016 2440
rect 49608 2388 49660 2440
rect 51264 2431 51316 2440
rect 51264 2397 51273 2431
rect 51273 2397 51307 2431
rect 51307 2397 51316 2431
rect 51264 2388 51316 2397
rect 51632 2388 51684 2440
rect 54024 2456 54076 2508
rect 53288 2388 53340 2440
rect 55772 2456 55824 2508
rect 57428 2456 57480 2508
rect 56324 2388 56376 2440
rect 51356 2320 51408 2372
rect 53656 2320 53708 2372
rect 46572 2252 46624 2304
rect 50896 2252 50948 2304
rect 51172 2252 51224 2304
rect 52000 2252 52052 2304
rect 53104 2252 53156 2304
rect 55496 2320 55548 2372
rect 55956 2320 56008 2372
rect 56140 2252 56192 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 8208 2048 8260 2100
rect 12716 2048 12768 2100
rect 17684 2048 17736 2100
rect 21640 2048 21692 2100
rect 40224 2048 40276 2100
rect 44364 2048 44416 2100
rect 46664 2048 46716 2100
rect 49884 2048 49936 2100
rect 9680 1980 9732 2032
rect 14832 1980 14884 2032
rect 41328 1980 41380 2032
rect 43904 1980 43956 2032
rect 44272 1980 44324 2032
rect 48228 1980 48280 2032
rect 10324 1912 10376 1964
rect 15384 1912 15436 1964
rect 40960 1912 41012 1964
rect 48504 1912 48556 1964
rect 12164 1844 12216 1896
rect 16304 1844 16356 1896
rect 45100 1844 45152 1896
rect 47400 1844 47452 1896
rect 11704 1776 11756 1828
rect 12992 1776 13044 1828
rect 41236 1776 41288 1828
rect 42708 1776 42760 1828
rect 45560 1776 45612 1828
rect 49148 1776 49200 1828
rect 49608 1776 49660 1828
rect 11428 1708 11480 1760
rect 12900 1708 12952 1760
rect 16120 1708 16172 1760
rect 16396 1708 16448 1760
rect 47216 1708 47268 1760
rect 47860 1708 47912 1760
rect 10692 1640 10744 1692
rect 12808 1640 12860 1692
rect 48964 1572 49016 1624
rect 52368 1572 52420 1624
rect 13912 1368 13964 1420
rect 14648 1368 14700 1420
rect 17684 1368 17736 1420
rect 11612 1164 11664 1216
rect 14188 1164 14240 1216
rect 15016 1164 15068 1216
rect 14740 1096 14792 1148
rect 14740 892 14792 944
rect 15016 892 15068 944
rect 15108 892 15160 944
<< metal2 >>
rect 3790 59200 3846 60000
rect 4342 59200 4398 60000
rect 4894 59200 4950 60000
rect 5446 59200 5502 60000
rect 5998 59200 6054 60000
rect 6550 59200 6606 60000
rect 7102 59200 7158 60000
rect 7654 59200 7710 60000
rect 8206 59200 8262 60000
rect 8758 59200 8814 60000
rect 9310 59200 9366 60000
rect 9862 59200 9918 60000
rect 10414 59200 10470 60000
rect 10966 59200 11022 60000
rect 11518 59200 11574 60000
rect 12070 59200 12126 60000
rect 12622 59200 12678 60000
rect 13174 59200 13230 60000
rect 13726 59200 13782 60000
rect 14278 59200 14334 60000
rect 14830 59200 14886 60000
rect 15382 59200 15438 60000
rect 15934 59200 15990 60000
rect 16486 59200 16542 60000
rect 17038 59200 17094 60000
rect 17590 59200 17646 60000
rect 18142 59200 18198 60000
rect 18694 59200 18750 60000
rect 19246 59200 19302 60000
rect 19798 59200 19854 60000
rect 20350 59200 20406 60000
rect 20902 59200 20958 60000
rect 21454 59200 21510 60000
rect 22006 59200 22062 60000
rect 22558 59200 22614 60000
rect 23110 59200 23166 60000
rect 23662 59200 23718 60000
rect 24214 59200 24270 60000
rect 24766 59200 24822 60000
rect 25318 59200 25374 60000
rect 25870 59200 25926 60000
rect 26422 59200 26478 60000
rect 26974 59200 27030 60000
rect 27526 59200 27582 60000
rect 28078 59200 28134 60000
rect 28630 59200 28686 60000
rect 29182 59200 29238 60000
rect 29734 59200 29790 60000
rect 30286 59200 30342 60000
rect 30838 59200 30894 60000
rect 31390 59200 31446 60000
rect 31942 59200 31998 60000
rect 32494 59200 32550 60000
rect 33046 59200 33102 60000
rect 33598 59200 33654 60000
rect 34150 59200 34206 60000
rect 34702 59200 34758 60000
rect 35254 59200 35310 60000
rect 35806 59200 35862 60000
rect 36358 59200 36414 60000
rect 36910 59200 36966 60000
rect 37462 59200 37518 60000
rect 38014 59200 38070 60000
rect 38566 59200 38622 60000
rect 39118 59200 39174 60000
rect 39670 59200 39726 60000
rect 39776 59214 39988 59242
rect 4356 57458 4384 59200
rect 4908 57458 4936 59200
rect 6012 57458 6040 59200
rect 6564 57458 6592 59200
rect 7668 57458 7696 59200
rect 8220 57458 8248 59200
rect 9324 57458 9352 59200
rect 9876 57458 9904 59200
rect 10980 57458 11008 59200
rect 11532 57458 11560 59200
rect 12636 57458 12664 59200
rect 13188 57458 13216 59200
rect 14292 57458 14320 59200
rect 14844 57458 14872 59200
rect 15948 57458 15976 59200
rect 4344 57452 4396 57458
rect 4344 57394 4396 57400
rect 4896 57452 4948 57458
rect 4896 57394 4948 57400
rect 6000 57452 6052 57458
rect 6000 57394 6052 57400
rect 6552 57452 6604 57458
rect 6552 57394 6604 57400
rect 7656 57452 7708 57458
rect 7656 57394 7708 57400
rect 8208 57452 8260 57458
rect 8208 57394 8260 57400
rect 9312 57452 9364 57458
rect 9312 57394 9364 57400
rect 9864 57452 9916 57458
rect 9864 57394 9916 57400
rect 10968 57452 11020 57458
rect 10968 57394 11020 57400
rect 11520 57452 11572 57458
rect 11520 57394 11572 57400
rect 12624 57452 12676 57458
rect 12624 57394 12676 57400
rect 13176 57452 13228 57458
rect 13176 57394 13228 57400
rect 14280 57452 14332 57458
rect 14280 57394 14332 57400
rect 14832 57452 14884 57458
rect 14832 57394 14884 57400
rect 15936 57452 15988 57458
rect 15936 57394 15988 57400
rect 16500 57390 16528 59200
rect 17604 57458 17632 59200
rect 18156 57458 18184 59200
rect 19260 57458 19288 59200
rect 19812 58290 19840 59200
rect 19812 58262 20024 58290
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 19996 57458 20024 58262
rect 20916 57458 20944 59200
rect 21468 57458 21496 59200
rect 22572 57458 22600 59200
rect 23124 57458 23152 59200
rect 17592 57452 17644 57458
rect 17592 57394 17644 57400
rect 18144 57452 18196 57458
rect 18144 57394 18196 57400
rect 19248 57452 19300 57458
rect 19248 57394 19300 57400
rect 19984 57452 20036 57458
rect 19984 57394 20036 57400
rect 20904 57452 20956 57458
rect 20904 57394 20956 57400
rect 21456 57452 21508 57458
rect 21456 57394 21508 57400
rect 22560 57452 22612 57458
rect 22560 57394 22612 57400
rect 23112 57452 23164 57458
rect 23112 57394 23164 57400
rect 16488 57384 16540 57390
rect 16488 57326 16540 57332
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 24228 57050 24256 59200
rect 24780 57440 24808 59200
rect 25884 57458 25912 59200
rect 26436 57458 26464 59200
rect 27540 57458 27568 59200
rect 28092 57458 28120 59200
rect 29196 57458 29224 59200
rect 29748 57458 29776 59200
rect 30852 57458 30880 59200
rect 31404 57458 31432 59200
rect 32508 57458 32536 59200
rect 24860 57452 24912 57458
rect 24780 57412 24860 57440
rect 24860 57394 24912 57400
rect 25872 57452 25924 57458
rect 25872 57394 25924 57400
rect 26424 57452 26476 57458
rect 26424 57394 26476 57400
rect 27528 57452 27580 57458
rect 27528 57394 27580 57400
rect 28080 57452 28132 57458
rect 28080 57394 28132 57400
rect 29184 57452 29236 57458
rect 29184 57394 29236 57400
rect 29736 57452 29788 57458
rect 29736 57394 29788 57400
rect 30840 57452 30892 57458
rect 30840 57394 30892 57400
rect 31392 57452 31444 57458
rect 31392 57394 31444 57400
rect 32496 57452 32548 57458
rect 33060 57440 33088 59200
rect 34164 57458 34192 59200
rect 34716 57458 34744 59200
rect 33140 57452 33192 57458
rect 33060 57412 33140 57440
rect 32496 57394 32548 57400
rect 33140 57394 33192 57400
rect 34152 57452 34204 57458
rect 34152 57394 34204 57400
rect 34704 57452 34756 57458
rect 34704 57394 34756 57400
rect 35820 57390 35848 59200
rect 36372 57458 36400 59200
rect 37476 57458 37504 59200
rect 38028 57458 38056 59200
rect 39132 57458 39160 59200
rect 39684 59106 39712 59200
rect 39776 59106 39804 59214
rect 39684 59078 39804 59106
rect 36360 57452 36412 57458
rect 36360 57394 36412 57400
rect 37464 57452 37516 57458
rect 37464 57394 37516 57400
rect 38016 57452 38068 57458
rect 38016 57394 38068 57400
rect 39120 57452 39172 57458
rect 39960 57440 39988 59214
rect 40222 59200 40278 60000
rect 40774 59200 40830 60000
rect 41326 59200 41382 60000
rect 41878 59200 41934 60000
rect 42430 59200 42486 60000
rect 42982 59200 43038 60000
rect 43534 59200 43590 60000
rect 44086 59200 44142 60000
rect 44638 59200 44694 60000
rect 45190 59200 45246 60000
rect 45742 59200 45798 60000
rect 46294 59200 46350 60000
rect 46846 59200 46902 60000
rect 47398 59200 47454 60000
rect 47950 59200 48006 60000
rect 48502 59200 48558 60000
rect 49054 59200 49110 60000
rect 49606 59200 49662 60000
rect 50158 59200 50214 60000
rect 50710 59200 50766 60000
rect 51262 59200 51318 60000
rect 51814 59200 51870 60000
rect 52366 59200 52422 60000
rect 52918 59200 52974 60000
rect 53470 59200 53526 60000
rect 54022 59200 54078 60000
rect 54574 59200 54630 60000
rect 55126 59200 55182 60000
rect 55678 59200 55734 60000
rect 56230 59200 56286 60000
rect 56336 59214 56548 59242
rect 40788 57458 40816 59200
rect 40040 57452 40092 57458
rect 39960 57412 40040 57440
rect 39120 57394 39172 57400
rect 40040 57394 40092 57400
rect 40776 57452 40828 57458
rect 41340 57440 41368 59200
rect 42444 57458 42472 59200
rect 42996 57458 43024 59200
rect 42432 57452 42484 57458
rect 41340 57412 41460 57440
rect 40776 57394 40828 57400
rect 35808 57384 35860 57390
rect 35808 57326 35860 57332
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 41432 57050 41460 57412
rect 42432 57394 42484 57400
rect 42984 57452 43036 57458
rect 44100 57440 44128 59200
rect 44652 57458 44680 59200
rect 45756 57458 45784 59200
rect 46308 57458 46336 59200
rect 47412 57458 47440 59200
rect 47964 57458 47992 59200
rect 49068 57458 49096 59200
rect 49620 57474 49648 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 49620 57458 49740 57474
rect 50724 57458 50752 59200
rect 51276 57458 51304 59200
rect 52380 57474 52408 59200
rect 52380 57458 52500 57474
rect 52932 57458 52960 59200
rect 54036 57458 54064 59200
rect 44180 57452 44232 57458
rect 44100 57412 44180 57440
rect 42984 57394 43036 57400
rect 44180 57394 44232 57400
rect 44640 57452 44692 57458
rect 44640 57394 44692 57400
rect 45744 57452 45796 57458
rect 45744 57394 45796 57400
rect 46296 57452 46348 57458
rect 46296 57394 46348 57400
rect 47400 57452 47452 57458
rect 47400 57394 47452 57400
rect 47952 57452 48004 57458
rect 47952 57394 48004 57400
rect 49056 57452 49108 57458
rect 49620 57452 49752 57458
rect 49620 57446 49700 57452
rect 49056 57394 49108 57400
rect 49700 57394 49752 57400
rect 50712 57452 50764 57458
rect 50712 57394 50764 57400
rect 51264 57452 51316 57458
rect 52380 57452 52512 57458
rect 52380 57446 52460 57452
rect 51264 57394 51316 57400
rect 52460 57394 52512 57400
rect 52920 57452 52972 57458
rect 52920 57394 52972 57400
rect 54024 57452 54076 57458
rect 54024 57394 54076 57400
rect 54588 57322 54616 59200
rect 55692 57458 55720 59200
rect 56244 59106 56272 59200
rect 56336 59106 56364 59214
rect 56244 59078 56364 59106
rect 56520 57882 56548 59214
rect 56782 59200 56838 60000
rect 57334 59200 57390 60000
rect 57886 59200 57942 60000
rect 58438 59200 58494 60000
rect 58990 59200 59046 60000
rect 59542 59200 59598 60000
rect 60094 59200 60150 60000
rect 60646 59200 60702 60000
rect 61198 59200 61254 60000
rect 61750 59200 61806 60000
rect 62302 59200 62358 60000
rect 62854 59200 62910 60000
rect 63406 59200 63462 60000
rect 63958 59200 64014 60000
rect 64510 59200 64566 60000
rect 65062 59200 65118 60000
rect 65614 59200 65670 60000
rect 66166 59200 66222 60000
rect 56520 57854 56640 57882
rect 56612 57458 56640 57854
rect 57348 57458 57376 59200
rect 57900 57474 57928 59200
rect 57900 57458 58020 57474
rect 59004 57458 59032 59200
rect 59556 57458 59584 59200
rect 60660 57474 60688 59200
rect 60660 57458 60780 57474
rect 61212 57458 61240 59200
rect 62316 57458 62344 59200
rect 55680 57452 55732 57458
rect 55680 57394 55732 57400
rect 56600 57452 56652 57458
rect 56600 57394 56652 57400
rect 57336 57452 57388 57458
rect 57900 57452 58032 57458
rect 57900 57446 57980 57452
rect 57336 57394 57388 57400
rect 57980 57394 58032 57400
rect 58992 57452 59044 57458
rect 58992 57394 59044 57400
rect 59544 57452 59596 57458
rect 60660 57452 60792 57458
rect 60660 57446 60740 57452
rect 59544 57394 59596 57400
rect 60740 57394 60792 57400
rect 61200 57452 61252 57458
rect 61200 57394 61252 57400
rect 62304 57452 62356 57458
rect 62304 57394 62356 57400
rect 62868 57390 62896 59200
rect 63972 57458 64000 59200
rect 63960 57452 64012 57458
rect 63960 57394 64012 57400
rect 62856 57384 62908 57390
rect 62856 57326 62908 57332
rect 54576 57316 54628 57322
rect 54576 57258 54628 57264
rect 64524 57050 64552 59200
rect 65628 57458 65656 59200
rect 66180 57474 66208 59200
rect 66180 57458 66300 57474
rect 65616 57452 65668 57458
rect 66180 57452 66312 57458
rect 66180 57446 66260 57452
rect 65616 57394 65668 57400
rect 66260 57394 66312 57400
rect 65654 57148 65962 57157
rect 65654 57146 65660 57148
rect 65716 57146 65740 57148
rect 65796 57146 65820 57148
rect 65876 57146 65900 57148
rect 65956 57146 65962 57148
rect 65716 57094 65718 57146
rect 65898 57094 65900 57146
rect 65654 57092 65660 57094
rect 65716 57092 65740 57094
rect 65796 57092 65820 57094
rect 65876 57092 65900 57094
rect 65956 57092 65962 57094
rect 65654 57083 65962 57092
rect 24216 57044 24268 57050
rect 24216 56986 24268 56992
rect 41420 57044 41472 57050
rect 41420 56986 41472 56992
rect 64512 57044 64564 57050
rect 64512 56986 64564 56992
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 67364 56364 67416 56370
rect 67364 56306 67416 56312
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 65654 56060 65962 56069
rect 65654 56058 65660 56060
rect 65716 56058 65740 56060
rect 65796 56058 65820 56060
rect 65876 56058 65900 56060
rect 65956 56058 65962 56060
rect 65716 56006 65718 56058
rect 65898 56006 65900 56058
rect 65654 56004 65660 56006
rect 65716 56004 65740 56006
rect 65796 56004 65820 56006
rect 65876 56004 65900 56006
rect 65956 56004 65962 56006
rect 65654 55995 65962 56004
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 65654 54972 65962 54981
rect 65654 54970 65660 54972
rect 65716 54970 65740 54972
rect 65796 54970 65820 54972
rect 65876 54970 65900 54972
rect 65956 54970 65962 54972
rect 65716 54918 65718 54970
rect 65898 54918 65900 54970
rect 65654 54916 65660 54918
rect 65716 54916 65740 54918
rect 65796 54916 65820 54918
rect 65876 54916 65900 54918
rect 65956 54916 65962 54918
rect 65654 54907 65962 54916
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 65654 53884 65962 53893
rect 65654 53882 65660 53884
rect 65716 53882 65740 53884
rect 65796 53882 65820 53884
rect 65876 53882 65900 53884
rect 65956 53882 65962 53884
rect 65716 53830 65718 53882
rect 65898 53830 65900 53882
rect 65654 53828 65660 53830
rect 65716 53828 65740 53830
rect 65796 53828 65820 53830
rect 65876 53828 65900 53830
rect 65956 53828 65962 53830
rect 65654 53819 65962 53828
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 65654 52796 65962 52805
rect 65654 52794 65660 52796
rect 65716 52794 65740 52796
rect 65796 52794 65820 52796
rect 65876 52794 65900 52796
rect 65956 52794 65962 52796
rect 65716 52742 65718 52794
rect 65898 52742 65900 52794
rect 65654 52740 65660 52742
rect 65716 52740 65740 52742
rect 65796 52740 65820 52742
rect 65876 52740 65900 52742
rect 65956 52740 65962 52742
rect 65654 52731 65962 52740
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 65654 51708 65962 51717
rect 65654 51706 65660 51708
rect 65716 51706 65740 51708
rect 65796 51706 65820 51708
rect 65876 51706 65900 51708
rect 65956 51706 65962 51708
rect 65716 51654 65718 51706
rect 65898 51654 65900 51706
rect 65654 51652 65660 51654
rect 65716 51652 65740 51654
rect 65796 51652 65820 51654
rect 65876 51652 65900 51654
rect 65956 51652 65962 51654
rect 65654 51643 65962 51652
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 65654 50620 65962 50629
rect 65654 50618 65660 50620
rect 65716 50618 65740 50620
rect 65796 50618 65820 50620
rect 65876 50618 65900 50620
rect 65956 50618 65962 50620
rect 65716 50566 65718 50618
rect 65898 50566 65900 50618
rect 65654 50564 65660 50566
rect 65716 50564 65740 50566
rect 65796 50564 65820 50566
rect 65876 50564 65900 50566
rect 65956 50564 65962 50566
rect 65654 50555 65962 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 65654 49532 65962 49541
rect 65654 49530 65660 49532
rect 65716 49530 65740 49532
rect 65796 49530 65820 49532
rect 65876 49530 65900 49532
rect 65956 49530 65962 49532
rect 65716 49478 65718 49530
rect 65898 49478 65900 49530
rect 65654 49476 65660 49478
rect 65716 49476 65740 49478
rect 65796 49476 65820 49478
rect 65876 49476 65900 49478
rect 65956 49476 65962 49478
rect 65654 49467 65962 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 65654 48444 65962 48453
rect 65654 48442 65660 48444
rect 65716 48442 65740 48444
rect 65796 48442 65820 48444
rect 65876 48442 65900 48444
rect 65956 48442 65962 48444
rect 65716 48390 65718 48442
rect 65898 48390 65900 48442
rect 65654 48388 65660 48390
rect 65716 48388 65740 48390
rect 65796 48388 65820 48390
rect 65876 48388 65900 48390
rect 65956 48388 65962 48390
rect 65654 48379 65962 48388
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 65654 47356 65962 47365
rect 65654 47354 65660 47356
rect 65716 47354 65740 47356
rect 65796 47354 65820 47356
rect 65876 47354 65900 47356
rect 65956 47354 65962 47356
rect 65716 47302 65718 47354
rect 65898 47302 65900 47354
rect 65654 47300 65660 47302
rect 65716 47300 65740 47302
rect 65796 47300 65820 47302
rect 65876 47300 65900 47302
rect 65956 47300 65962 47302
rect 65654 47291 65962 47300
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 65654 46268 65962 46277
rect 65654 46266 65660 46268
rect 65716 46266 65740 46268
rect 65796 46266 65820 46268
rect 65876 46266 65900 46268
rect 65956 46266 65962 46268
rect 65716 46214 65718 46266
rect 65898 46214 65900 46266
rect 65654 46212 65660 46214
rect 65716 46212 65740 46214
rect 65796 46212 65820 46214
rect 65876 46212 65900 46214
rect 65956 46212 65962 46214
rect 65654 46203 65962 46212
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 43996 45484 44048 45490
rect 43996 45426 44048 45432
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 44008 35894 44036 45426
rect 67376 45354 67404 56306
rect 67548 56160 67600 56166
rect 67546 56128 67548 56137
rect 67600 56128 67602 56137
rect 67546 56063 67602 56072
rect 67456 48748 67508 48754
rect 67456 48690 67508 48696
rect 67364 45348 67416 45354
rect 67364 45290 67416 45296
rect 65654 45180 65962 45189
rect 65654 45178 65660 45180
rect 65716 45178 65740 45180
rect 65796 45178 65820 45180
rect 65876 45178 65900 45180
rect 65956 45178 65962 45180
rect 65716 45126 65718 45178
rect 65898 45126 65900 45178
rect 65654 45124 65660 45126
rect 65716 45124 65740 45126
rect 65796 45124 65820 45126
rect 65876 45124 65900 45126
rect 65956 45124 65962 45126
rect 65654 45115 65962 45124
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 65654 44092 65962 44101
rect 65654 44090 65660 44092
rect 65716 44090 65740 44092
rect 65796 44090 65820 44092
rect 65876 44090 65900 44092
rect 65956 44090 65962 44092
rect 65716 44038 65718 44090
rect 65898 44038 65900 44090
rect 65654 44036 65660 44038
rect 65716 44036 65740 44038
rect 65796 44036 65820 44038
rect 65876 44036 65900 44038
rect 65956 44036 65962 44038
rect 65654 44027 65962 44036
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 65654 43004 65962 43013
rect 65654 43002 65660 43004
rect 65716 43002 65740 43004
rect 65796 43002 65820 43004
rect 65876 43002 65900 43004
rect 65956 43002 65962 43004
rect 65716 42950 65718 43002
rect 65898 42950 65900 43002
rect 65654 42948 65660 42950
rect 65716 42948 65740 42950
rect 65796 42948 65820 42950
rect 65876 42948 65900 42950
rect 65956 42948 65962 42950
rect 65654 42939 65962 42948
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 65654 41916 65962 41925
rect 65654 41914 65660 41916
rect 65716 41914 65740 41916
rect 65796 41914 65820 41916
rect 65876 41914 65900 41916
rect 65956 41914 65962 41916
rect 65716 41862 65718 41914
rect 65898 41862 65900 41914
rect 65654 41860 65660 41862
rect 65716 41860 65740 41862
rect 65796 41860 65820 41862
rect 65876 41860 65900 41862
rect 65956 41860 65962 41862
rect 65654 41851 65962 41860
rect 67272 41472 67324 41478
rect 67272 41414 67324 41420
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 65654 40828 65962 40837
rect 65654 40826 65660 40828
rect 65716 40826 65740 40828
rect 65796 40826 65820 40828
rect 65876 40826 65900 40828
rect 65956 40826 65962 40828
rect 65716 40774 65718 40826
rect 65898 40774 65900 40826
rect 65654 40772 65660 40774
rect 65716 40772 65740 40774
rect 65796 40772 65820 40774
rect 65876 40772 65900 40774
rect 65956 40772 65962 40774
rect 65654 40763 65962 40772
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 65654 39740 65962 39749
rect 65654 39738 65660 39740
rect 65716 39738 65740 39740
rect 65796 39738 65820 39740
rect 65876 39738 65900 39740
rect 65956 39738 65962 39740
rect 65716 39686 65718 39738
rect 65898 39686 65900 39738
rect 65654 39684 65660 39686
rect 65716 39684 65740 39686
rect 65796 39684 65820 39686
rect 65876 39684 65900 39686
rect 65956 39684 65962 39686
rect 65654 39675 65962 39684
rect 67180 39432 67232 39438
rect 67180 39374 67232 39380
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 65654 38652 65962 38661
rect 65654 38650 65660 38652
rect 65716 38650 65740 38652
rect 65796 38650 65820 38652
rect 65876 38650 65900 38652
rect 65956 38650 65962 38652
rect 65716 38598 65718 38650
rect 65898 38598 65900 38650
rect 65654 38596 65660 38598
rect 65716 38596 65740 38598
rect 65796 38596 65820 38598
rect 65876 38596 65900 38598
rect 65956 38596 65962 38598
rect 65654 38587 65962 38596
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 65654 37564 65962 37573
rect 65654 37562 65660 37564
rect 65716 37562 65740 37564
rect 65796 37562 65820 37564
rect 65876 37562 65900 37564
rect 65956 37562 65962 37564
rect 65716 37510 65718 37562
rect 65898 37510 65900 37562
rect 65654 37508 65660 37510
rect 65716 37508 65740 37510
rect 65796 37508 65820 37510
rect 65876 37508 65900 37510
rect 65956 37508 65962 37510
rect 65654 37499 65962 37508
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 65654 36476 65962 36485
rect 65654 36474 65660 36476
rect 65716 36474 65740 36476
rect 65796 36474 65820 36476
rect 65876 36474 65900 36476
rect 65956 36474 65962 36476
rect 65716 36422 65718 36474
rect 65898 36422 65900 36474
rect 65654 36420 65660 36422
rect 65716 36420 65740 36422
rect 65796 36420 65820 36422
rect 65876 36420 65900 36422
rect 65956 36420 65962 36422
rect 65654 36411 65962 36420
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 44008 35866 44128 35894
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 27620 34400 27672 34406
rect 27620 34342 27672 34348
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 26884 34128 26936 34134
rect 26884 34070 26936 34076
rect 26896 33998 26924 34070
rect 27252 34060 27304 34066
rect 27252 34002 27304 34008
rect 26884 33992 26936 33998
rect 26804 33940 26884 33946
rect 26804 33934 26936 33940
rect 26804 33918 26924 33934
rect 27068 33924 27120 33930
rect 12900 33856 12952 33862
rect 12900 33798 12952 33804
rect 7472 33516 7524 33522
rect 7472 33458 7524 33464
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 7104 32428 7156 32434
rect 7104 32370 7156 32376
rect 6368 32224 6420 32230
rect 6368 32166 6420 32172
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 5264 31816 5316 31822
rect 5264 31758 5316 31764
rect 5276 31226 5304 31758
rect 5540 31748 5592 31754
rect 5540 31690 5592 31696
rect 5276 31210 5488 31226
rect 5276 31204 5500 31210
rect 5276 31198 5448 31204
rect 5448 31146 5500 31152
rect 5172 31136 5224 31142
rect 5172 31078 5224 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 5080 30796 5132 30802
rect 5080 30738 5132 30744
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4988 29640 5040 29646
rect 5092 29594 5120 30738
rect 5184 30734 5212 31078
rect 5460 30802 5488 31146
rect 5552 30938 5580 31690
rect 5632 31680 5684 31686
rect 5632 31622 5684 31628
rect 5644 31482 5672 31622
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 5540 30932 5592 30938
rect 5540 30874 5592 30880
rect 5448 30796 5500 30802
rect 5448 30738 5500 30744
rect 6380 30734 6408 32166
rect 7116 32026 7144 32370
rect 7104 32020 7156 32026
rect 7104 31962 7156 31968
rect 7012 31884 7064 31890
rect 7012 31826 7064 31832
rect 7024 31754 7052 31826
rect 7288 31816 7340 31822
rect 7288 31758 7340 31764
rect 7024 31726 7144 31754
rect 6460 31680 6512 31686
rect 6460 31622 6512 31628
rect 6472 31346 6500 31622
rect 7116 31482 7144 31726
rect 7104 31476 7156 31482
rect 7104 31418 7156 31424
rect 6460 31340 6512 31346
rect 6460 31282 6512 31288
rect 7116 30802 7144 31418
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 5172 30728 5224 30734
rect 5172 30670 5224 30676
rect 6368 30728 6420 30734
rect 6368 30670 6420 30676
rect 7012 29708 7064 29714
rect 7012 29650 7064 29656
rect 5040 29588 5120 29594
rect 4988 29582 5120 29588
rect 6736 29640 6788 29646
rect 6736 29582 6788 29588
rect 5000 29566 5120 29582
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 5092 27470 5120 29566
rect 5264 29572 5316 29578
rect 5264 29514 5316 29520
rect 5276 29306 5304 29514
rect 6748 29306 6776 29582
rect 5264 29300 5316 29306
rect 5264 29242 5316 29248
rect 6736 29300 6788 29306
rect 6736 29242 6788 29248
rect 6184 29232 6236 29238
rect 6184 29174 6236 29180
rect 5908 28076 5960 28082
rect 5908 28018 5960 28024
rect 4804 27464 4856 27470
rect 4804 27406 4856 27412
rect 5080 27464 5132 27470
rect 5080 27406 5132 27412
rect 4712 27328 4764 27334
rect 4712 27270 4764 27276
rect 4620 27056 4672 27062
rect 4620 26998 4672 27004
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25294 4660 26998
rect 4724 26994 4752 27270
rect 4712 26988 4764 26994
rect 4712 26930 4764 26936
rect 4816 26586 4844 27406
rect 5092 26994 5120 27406
rect 5080 26988 5132 26994
rect 5080 26930 5132 26936
rect 5172 26784 5224 26790
rect 5172 26726 5224 26732
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 5184 26382 5212 26726
rect 5724 26512 5776 26518
rect 5724 26454 5776 26460
rect 5448 26444 5500 26450
rect 5448 26386 5500 26392
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 4896 25900 4948 25906
rect 4896 25842 4948 25848
rect 4712 25696 4764 25702
rect 4712 25638 4764 25644
rect 4620 25288 4672 25294
rect 4620 25230 4672 25236
rect 4724 25226 4752 25638
rect 4908 25498 4936 25842
rect 4896 25492 4948 25498
rect 4896 25434 4948 25440
rect 4712 25220 4764 25226
rect 4712 25162 4764 25168
rect 5184 24818 5212 26318
rect 5460 25378 5488 26386
rect 5736 26042 5764 26454
rect 5724 26036 5776 26042
rect 5724 25978 5776 25984
rect 5460 25362 5580 25378
rect 5460 25356 5592 25362
rect 5460 25350 5540 25356
rect 5172 24812 5224 24818
rect 5172 24754 5224 24760
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4724 24274 4752 24550
rect 4712 24268 4764 24274
rect 4712 24210 4764 24216
rect 5356 24064 5408 24070
rect 5356 24006 5408 24012
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 5368 23118 5396 24006
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 5368 22234 5396 22578
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5368 21690 5396 22170
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5460 21418 5488 25350
rect 5540 25298 5592 25304
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 5644 23798 5672 25094
rect 5632 23792 5684 23798
rect 5632 23734 5684 23740
rect 5724 23588 5776 23594
rect 5724 23530 5776 23536
rect 5736 23118 5764 23530
rect 5816 23520 5868 23526
rect 5816 23462 5868 23468
rect 5828 23118 5856 23462
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5724 23112 5776 23118
rect 5724 23054 5776 23060
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 5552 22778 5580 23054
rect 5920 22964 5948 28018
rect 6000 27396 6052 27402
rect 6000 27338 6052 27344
rect 6012 26586 6040 27338
rect 6000 26580 6052 26586
rect 6000 26522 6052 26528
rect 5644 22936 5948 22964
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 5644 22094 5672 22936
rect 5908 22500 5960 22506
rect 5908 22442 5960 22448
rect 5552 22066 5672 22094
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 5552 20262 5580 22066
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5828 21690 5856 21966
rect 5920 21690 5948 22442
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5540 20256 5592 20262
rect 5540 20198 5592 20204
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 5552 19854 5580 20198
rect 5724 19916 5776 19922
rect 5724 19858 5776 19864
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 4620 19780 4672 19786
rect 4620 19722 4672 19728
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4448 19258 4476 19314
rect 4632 19258 4660 19722
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 4448 19230 4660 19258
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16794 4660 19230
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 5000 18970 5028 19110
rect 4988 18964 5040 18970
rect 4988 18906 5040 18912
rect 5460 18358 5488 19654
rect 5552 18970 5580 19790
rect 5736 19514 5764 19858
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5736 19242 5764 19450
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5736 18766 5764 19178
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 6196 18630 6224 29174
rect 7024 29170 7052 29650
rect 7012 29164 7064 29170
rect 7012 29106 7064 29112
rect 7024 28218 7052 29106
rect 7116 29102 7144 30738
rect 7104 29096 7156 29102
rect 7104 29038 7156 29044
rect 7012 28212 7064 28218
rect 7012 28154 7064 28160
rect 6460 28008 6512 28014
rect 6460 27950 6512 27956
rect 6472 27674 6500 27950
rect 6460 27668 6512 27674
rect 6460 27610 6512 27616
rect 6368 26920 6420 26926
rect 6368 26862 6420 26868
rect 6380 25974 6408 26862
rect 6472 26738 6500 27610
rect 6920 27328 6972 27334
rect 6920 27270 6972 27276
rect 6932 27062 6960 27270
rect 6920 27056 6972 27062
rect 6920 26998 6972 27004
rect 6552 26784 6604 26790
rect 6472 26732 6552 26738
rect 6472 26726 6604 26732
rect 6472 26710 6592 26726
rect 7116 26450 7144 29038
rect 7300 26518 7328 31758
rect 7484 31686 7512 33458
rect 12532 33448 12584 33454
rect 12532 33390 12584 33396
rect 9772 33380 9824 33386
rect 9772 33322 9824 33328
rect 9784 32978 9812 33322
rect 11152 33312 11204 33318
rect 11152 33254 11204 33260
rect 9772 32972 9824 32978
rect 9772 32914 9824 32920
rect 11164 32910 11192 33254
rect 12544 33046 12572 33390
rect 12912 33046 12940 33798
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 13176 33652 13228 33658
rect 13176 33594 13228 33600
rect 13188 33386 13216 33594
rect 14280 33584 14332 33590
rect 14280 33526 14332 33532
rect 13268 33516 13320 33522
rect 13268 33458 13320 33464
rect 13176 33380 13228 33386
rect 13176 33322 13228 33328
rect 12532 33040 12584 33046
rect 12532 32982 12584 32988
rect 12900 33040 12952 33046
rect 12900 32982 12952 32988
rect 12912 32910 12940 32982
rect 12992 32972 13044 32978
rect 12992 32914 13044 32920
rect 11152 32904 11204 32910
rect 11152 32846 11204 32852
rect 12900 32904 12952 32910
rect 12900 32846 12952 32852
rect 10232 32768 10284 32774
rect 10232 32710 10284 32716
rect 9036 32428 9088 32434
rect 9036 32370 9088 32376
rect 7472 31680 7524 31686
rect 7472 31622 7524 31628
rect 7484 30938 7512 31622
rect 8392 31340 8444 31346
rect 8392 31282 8444 31288
rect 8300 31204 8352 31210
rect 8300 31146 8352 31152
rect 7472 30932 7524 30938
rect 7472 30874 7524 30880
rect 8312 30734 8340 31146
rect 8404 30938 8432 31282
rect 9048 31210 9076 32370
rect 9680 32224 9732 32230
rect 9680 32166 9732 32172
rect 9036 31204 9088 31210
rect 9036 31146 9088 31152
rect 9692 31142 9720 32166
rect 10244 31346 10272 32710
rect 12808 32360 12860 32366
rect 12808 32302 12860 32308
rect 12072 31816 12124 31822
rect 12072 31758 12124 31764
rect 9772 31340 9824 31346
rect 9772 31282 9824 31288
rect 9956 31340 10008 31346
rect 9956 31282 10008 31288
rect 10232 31340 10284 31346
rect 10232 31282 10284 31288
rect 8484 31136 8536 31142
rect 8484 31078 8536 31084
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 8496 30938 8524 31078
rect 8392 30932 8444 30938
rect 8392 30874 8444 30880
rect 8484 30932 8536 30938
rect 8484 30874 8536 30880
rect 8300 30728 8352 30734
rect 8300 30670 8352 30676
rect 7932 30660 7984 30666
rect 7932 30602 7984 30608
rect 7380 27464 7432 27470
rect 7380 27406 7432 27412
rect 7392 26586 7420 27406
rect 7748 27396 7800 27402
rect 7748 27338 7800 27344
rect 7760 27130 7788 27338
rect 7748 27124 7800 27130
rect 7748 27066 7800 27072
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 7288 26512 7340 26518
rect 7288 26454 7340 26460
rect 7104 26444 7156 26450
rect 7104 26386 7156 26392
rect 7564 26444 7616 26450
rect 7564 26386 7616 26392
rect 6920 26308 6972 26314
rect 6920 26250 6972 26256
rect 6368 25968 6420 25974
rect 6368 25910 6420 25916
rect 6644 24744 6696 24750
rect 6644 24686 6696 24692
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6564 23662 6592 24142
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 6368 23044 6420 23050
rect 6368 22986 6420 22992
rect 6380 22778 6408 22986
rect 6368 22772 6420 22778
rect 6368 22714 6420 22720
rect 6656 22098 6684 24686
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6748 23730 6776 24006
rect 6736 23724 6788 23730
rect 6736 23666 6788 23672
rect 6644 22092 6696 22098
rect 6644 22034 6696 22040
rect 6656 21010 6684 22034
rect 6932 21010 6960 26250
rect 7576 25430 7604 26386
rect 7760 26314 7788 27066
rect 7748 26308 7800 26314
rect 7748 26250 7800 26256
rect 7944 26042 7972 30602
rect 9784 30394 9812 31282
rect 9772 30388 9824 30394
rect 9772 30330 9824 30336
rect 9968 29782 9996 31282
rect 12084 30734 12112 31758
rect 12624 31748 12676 31754
rect 12624 31690 12676 31696
rect 12636 31482 12664 31690
rect 12624 31476 12676 31482
rect 12624 31418 12676 31424
rect 12072 30728 12124 30734
rect 12072 30670 12124 30676
rect 11704 30660 11756 30666
rect 11704 30602 11756 30608
rect 11716 30394 11744 30602
rect 12164 30592 12216 30598
rect 12164 30534 12216 30540
rect 11704 30388 11756 30394
rect 11704 30330 11756 30336
rect 11152 30252 11204 30258
rect 11152 30194 11204 30200
rect 11796 30252 11848 30258
rect 11796 30194 11848 30200
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 9956 29776 10008 29782
rect 9956 29718 10008 29724
rect 9128 29640 9180 29646
rect 9128 29582 9180 29588
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 9140 28762 9168 29582
rect 10324 29164 10376 29170
rect 10324 29106 10376 29112
rect 9588 29096 9640 29102
rect 9588 29038 9640 29044
rect 9128 28756 9180 28762
rect 9128 28698 9180 28704
rect 9600 28558 9628 29038
rect 10336 28762 10364 29106
rect 10324 28756 10376 28762
rect 10324 28698 10376 28704
rect 9680 28620 9732 28626
rect 9680 28562 9732 28568
rect 9588 28552 9640 28558
rect 9588 28494 9640 28500
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 8300 27872 8352 27878
rect 8300 27814 8352 27820
rect 8312 26994 8340 27814
rect 8760 27464 8812 27470
rect 8760 27406 8812 27412
rect 8772 27130 8800 27406
rect 9220 27396 9272 27402
rect 9220 27338 9272 27344
rect 8760 27124 8812 27130
rect 8760 27066 8812 27072
rect 8300 26988 8352 26994
rect 8300 26930 8352 26936
rect 8312 26314 8340 26930
rect 9128 26784 9180 26790
rect 9128 26726 9180 26732
rect 9140 26518 9168 26726
rect 9232 26586 9260 27338
rect 9324 27334 9352 28358
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 9220 26580 9272 26586
rect 9220 26522 9272 26528
rect 9128 26512 9180 26518
rect 9128 26454 9180 26460
rect 8300 26308 8352 26314
rect 8300 26250 8352 26256
rect 7932 26036 7984 26042
rect 7932 25978 7984 25984
rect 7564 25424 7616 25430
rect 7564 25366 7616 25372
rect 7944 25294 7972 25978
rect 7932 25288 7984 25294
rect 7932 25230 7984 25236
rect 7944 24818 7972 25230
rect 7380 24812 7432 24818
rect 7932 24812 7984 24818
rect 7380 24754 7432 24760
rect 7852 24772 7932 24800
rect 7392 23866 7420 24754
rect 7852 24274 7880 24772
rect 7932 24754 7984 24760
rect 9128 24608 9180 24614
rect 9128 24550 9180 24556
rect 9140 24410 9168 24550
rect 9128 24404 9180 24410
rect 9128 24346 9180 24352
rect 7840 24268 7892 24274
rect 7840 24210 7892 24216
rect 9140 24206 9168 24346
rect 8024 24200 8076 24206
rect 8024 24142 8076 24148
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7380 23860 7432 23866
rect 7380 23802 7432 23808
rect 7576 23730 7604 24006
rect 8036 23730 8064 24142
rect 8116 24132 8168 24138
rect 8116 24074 8168 24080
rect 8300 24132 8352 24138
rect 8300 24074 8352 24080
rect 8128 23866 8156 24074
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 8312 23730 8340 24074
rect 8852 24064 8904 24070
rect 8852 24006 8904 24012
rect 8864 23730 8892 24006
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 8024 23724 8076 23730
rect 8024 23666 8076 23672
rect 8300 23724 8352 23730
rect 8300 23666 8352 23672
rect 8852 23724 8904 23730
rect 8852 23666 8904 23672
rect 8312 23322 8340 23666
rect 9128 23520 9180 23526
rect 9128 23462 9180 23468
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 7932 22432 7984 22438
rect 7932 22374 7984 22380
rect 7944 21554 7972 22374
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8220 21554 8248 21898
rect 7104 21548 7156 21554
rect 7104 21490 7156 21496
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 8208 21548 8260 21554
rect 8208 21490 8260 21496
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 7024 21078 7052 21422
rect 7012 21072 7064 21078
rect 7012 21014 7064 21020
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 7116 20874 7144 21490
rect 7564 21412 7616 21418
rect 7564 21354 7616 21360
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 6276 20868 6328 20874
rect 6276 20810 6328 20816
rect 7104 20868 7156 20874
rect 7104 20810 7156 20816
rect 6288 20602 6316 20810
rect 7012 20800 7064 20806
rect 7012 20742 7064 20748
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 7024 20466 7052 20742
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 7392 20398 7420 21286
rect 7576 21010 7604 21354
rect 7564 21004 7616 21010
rect 7564 20946 7616 20952
rect 7380 20392 7432 20398
rect 7380 20334 7432 20340
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7116 19718 7144 19790
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 6564 19378 6592 19654
rect 7116 19446 7144 19654
rect 7104 19440 7156 19446
rect 7104 19382 7156 19388
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 7116 18834 7144 19382
rect 7380 19372 7432 19378
rect 7380 19314 7432 19320
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6460 18624 6512 18630
rect 6460 18566 6512 18572
rect 5448 18352 5500 18358
rect 5448 18294 5500 18300
rect 5460 17746 5488 18294
rect 6472 17814 6500 18566
rect 7392 18426 7420 19314
rect 7380 18420 7432 18426
rect 7380 18362 7432 18368
rect 6460 17808 6512 17814
rect 6460 17750 6512 17756
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5736 17202 5764 17614
rect 6472 17338 6500 17750
rect 7392 17746 7420 18362
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4356 16114 4384 16594
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15570 4660 16730
rect 4724 16522 4752 16934
rect 5736 16794 5764 17138
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 6932 16658 6960 17478
rect 6920 16652 6972 16658
rect 6920 16594 6972 16600
rect 7024 16590 7052 17478
rect 7484 17134 7512 18022
rect 7576 17270 7604 20946
rect 7944 20058 7972 21490
rect 8220 20942 8248 21490
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8220 19854 8248 20334
rect 8312 19990 8340 20946
rect 8404 20466 8432 21286
rect 8956 21146 8984 21422
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 9140 20602 9168 23462
rect 9220 20800 9272 20806
rect 9220 20742 9272 20748
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 9232 20466 9260 20742
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 9036 20460 9088 20466
rect 9036 20402 9088 20408
rect 9220 20460 9272 20466
rect 9220 20402 9272 20408
rect 8300 19984 8352 19990
rect 8300 19926 8352 19932
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7760 18290 7788 18566
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8128 17746 8156 18158
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 7668 17338 7696 17682
rect 8220 17626 8248 19790
rect 8312 19378 8340 19926
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8496 18426 8524 19858
rect 9048 19718 9076 20402
rect 9324 20398 9352 27270
rect 9600 26994 9628 28494
rect 9692 27062 9720 28562
rect 10980 28218 11008 29582
rect 11072 29034 11100 30126
rect 11164 29646 11192 30194
rect 11808 29850 11836 30194
rect 11796 29844 11848 29850
rect 11796 29786 11848 29792
rect 11152 29640 11204 29646
rect 11152 29582 11204 29588
rect 11796 29640 11848 29646
rect 11796 29582 11848 29588
rect 11704 29504 11756 29510
rect 11704 29446 11756 29452
rect 11716 29170 11744 29446
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 11704 29164 11756 29170
rect 11704 29106 11756 29112
rect 11060 29028 11112 29034
rect 11060 28970 11112 28976
rect 9956 28212 10008 28218
rect 9956 28154 10008 28160
rect 10968 28212 11020 28218
rect 10968 28154 11020 28160
rect 9968 27538 9996 28154
rect 11072 28082 11100 28970
rect 11164 28490 11192 29106
rect 11716 28694 11744 29106
rect 11704 28688 11756 28694
rect 11704 28630 11756 28636
rect 11612 28552 11664 28558
rect 11612 28494 11664 28500
rect 11152 28484 11204 28490
rect 11152 28426 11204 28432
rect 11060 28076 11112 28082
rect 11060 28018 11112 28024
rect 11164 27606 11192 28426
rect 11244 28008 11296 28014
rect 11244 27950 11296 27956
rect 11152 27600 11204 27606
rect 11152 27542 11204 27548
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 10232 27328 10284 27334
rect 10232 27270 10284 27276
rect 10244 27062 10272 27270
rect 9680 27056 9732 27062
rect 9680 26998 9732 27004
rect 10232 27056 10284 27062
rect 10232 26998 10284 27004
rect 9588 26988 9640 26994
rect 9588 26930 9640 26936
rect 9496 25900 9548 25906
rect 9496 25842 9548 25848
rect 9508 25498 9536 25842
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9496 21412 9548 21418
rect 9496 21354 9548 21360
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 9416 20942 9444 21286
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9508 20874 9536 21354
rect 9496 20868 9548 20874
rect 9496 20810 9548 20816
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 9220 20324 9272 20330
rect 9220 20266 9272 20272
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8128 17610 8248 17626
rect 8116 17604 8248 17610
rect 8168 17598 8248 17604
rect 8116 17546 8168 17552
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5184 15706 5212 16050
rect 6920 16040 6972 16046
rect 6840 15988 6920 15994
rect 6840 15982 6972 15988
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 6840 15966 6960 15982
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 5460 15502 5488 15914
rect 6460 15700 6512 15706
rect 6460 15642 6512 15648
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 6380 14618 6408 15370
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4724 12306 4752 13262
rect 4908 12986 4936 13874
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 5000 13326 5028 13670
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6104 12986 6132 13126
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6104 12714 6132 12922
rect 6472 12782 6500 15642
rect 6840 15638 6868 15966
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 6828 15632 6880 15638
rect 6828 15574 6880 15580
rect 7024 15162 7052 15642
rect 7116 15570 7144 17070
rect 7484 16250 7512 17070
rect 7668 16590 7696 17274
rect 8128 16658 8156 17546
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 7656 16584 7708 16590
rect 7656 16526 7708 16532
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7472 16244 7524 16250
rect 7472 16186 7524 16192
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7760 15706 7788 16050
rect 7852 16046 7880 16390
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7748 15700 7800 15706
rect 7748 15642 7800 15648
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6564 14414 6592 14758
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 7392 14278 7420 14894
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6748 13326 6776 13806
rect 7116 13802 7144 14214
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 6092 12708 6144 12714
rect 6092 12650 6144 12656
rect 4712 12300 4764 12306
rect 4712 12242 4764 12248
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4724 11218 4752 12242
rect 5644 12238 5672 12650
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5264 12164 5316 12170
rect 5264 12106 5316 12112
rect 5276 11898 5304 12106
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4724 7954 4752 11154
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 5184 10810 5212 11018
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 6472 10674 6500 12718
rect 7116 12170 7144 12786
rect 7392 12306 7420 14214
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7668 13530 7696 13670
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7668 12986 7696 13466
rect 7760 13326 7788 13738
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7656 12980 7708 12986
rect 7656 12922 7708 12928
rect 7760 12918 7788 13262
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7748 12912 7800 12918
rect 7748 12854 7800 12860
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 6748 11762 6776 12038
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 7300 11558 7328 12038
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 11354 7328 11494
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6748 10810 6776 11154
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4724 6866 4752 7890
rect 5368 7886 5396 8230
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5368 6866 5396 7278
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 5356 6860 5408 6866
rect 5356 6802 5408 6808
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 5368 5778 5396 6802
rect 6380 6798 6408 7142
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6472 6254 6500 10610
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6552 10124 6604 10130
rect 6552 10066 6604 10072
rect 6564 9518 6592 10066
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6656 8634 6684 9522
rect 6840 8634 6868 10406
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 6656 8090 6684 8570
rect 7392 8430 7420 12242
rect 7852 11762 7880 13126
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7944 11218 7972 12310
rect 8128 11898 8156 16594
rect 9048 16250 9076 16594
rect 9232 16590 9260 20266
rect 9508 19854 9536 20810
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9220 16584 9272 16590
rect 9220 16526 9272 16532
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8208 15360 8260 15366
rect 8208 15302 8260 15308
rect 8220 14414 8248 15302
rect 8312 15026 8340 15438
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8588 14822 8616 15846
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8312 12442 8340 12718
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8312 11762 8340 12378
rect 8404 11830 8432 13194
rect 8668 12776 8720 12782
rect 8588 12724 8668 12730
rect 8588 12718 8720 12724
rect 8588 12702 8708 12718
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8116 11688 8168 11694
rect 8036 11636 8116 11642
rect 8036 11630 8168 11636
rect 8036 11614 8156 11630
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 8036 10962 8064 11614
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 11098 8156 11494
rect 8404 11354 8432 11766
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8404 11234 8432 11290
rect 8312 11206 8432 11234
rect 8496 11218 8524 12582
rect 8588 12170 8616 12702
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8680 12442 8708 12582
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8680 12238 8708 12378
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8484 11212 8536 11218
rect 8128 11070 8248 11098
rect 8036 10934 8156 10962
rect 8128 10674 8156 10934
rect 8220 10674 8248 11070
rect 8312 10742 8340 11206
rect 8484 11154 8536 11160
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7668 10266 7696 10406
rect 7656 10260 7708 10266
rect 7656 10202 7708 10208
rect 8128 10130 8156 10610
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 8128 9110 8156 10066
rect 8220 10062 8248 10610
rect 8404 10538 8432 11086
rect 8588 11082 8616 12106
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8772 11762 8800 12038
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8576 11076 8628 11082
rect 8576 11018 8628 11024
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 9140 10198 9168 16458
rect 9324 12306 9352 19654
rect 9600 19310 9628 26930
rect 9692 26586 9720 26998
rect 10692 26920 10744 26926
rect 10692 26862 10744 26868
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 10232 26784 10284 26790
rect 10232 26726 10284 26732
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9784 26450 9812 26726
rect 9772 26444 9824 26450
rect 9772 26386 9824 26392
rect 10244 26382 10272 26726
rect 10704 26586 10732 26862
rect 10692 26580 10744 26586
rect 10692 26522 10744 26528
rect 10232 26376 10284 26382
rect 10232 26318 10284 26324
rect 10600 26308 10652 26314
rect 10600 26250 10652 26256
rect 10508 26036 10560 26042
rect 10508 25978 10560 25984
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9876 24954 9904 25230
rect 10520 24954 10548 25978
rect 10612 25906 10640 26250
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10692 24880 10744 24886
rect 10692 24822 10744 24828
rect 9772 24676 9824 24682
rect 9772 24618 9824 24624
rect 9784 24070 9812 24618
rect 10704 24070 10732 24822
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 10692 24064 10744 24070
rect 10692 24006 10744 24012
rect 9784 23730 9812 24006
rect 10140 23792 10192 23798
rect 10140 23734 10192 23740
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 10152 23594 10180 23734
rect 10704 23730 10732 24006
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 10692 23724 10744 23730
rect 10692 23666 10744 23672
rect 10140 23588 10192 23594
rect 10140 23530 10192 23536
rect 10416 23520 10468 23526
rect 10416 23462 10468 23468
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9784 20942 9812 21830
rect 10060 21554 10088 21966
rect 10244 21554 10272 21966
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 9588 19304 9640 19310
rect 9588 19246 9640 19252
rect 10336 18630 10364 20402
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10428 17678 10456 23462
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 10704 22030 10732 22170
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10784 21548 10836 21554
rect 10784 21490 10836 21496
rect 10796 21146 10824 21490
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10600 20256 10652 20262
rect 10600 20198 10652 20204
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 10612 19310 10640 20198
rect 10796 19786 10824 20198
rect 10784 19780 10836 19786
rect 10784 19722 10836 19728
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10428 17134 10456 17614
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10508 16992 10560 16998
rect 10508 16934 10560 16940
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9692 15434 9720 16662
rect 10520 16046 10548 16934
rect 10612 16454 10640 19246
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10796 17202 10824 17478
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10796 17066 10824 17138
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10612 15502 10640 16050
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 9680 15428 9732 15434
rect 9680 15370 9732 15376
rect 10140 15360 10192 15366
rect 10140 15302 10192 15308
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9968 14618 9996 14962
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10152 14414 10180 15302
rect 10612 15162 10640 15438
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10140 14408 10192 14414
rect 10140 14350 10192 14356
rect 10796 13938 10824 17002
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10888 13870 10916 23802
rect 11072 22778 11100 27406
rect 11256 27334 11284 27950
rect 11624 27674 11652 28494
rect 11808 28218 11836 29582
rect 12176 29578 12204 30534
rect 12164 29572 12216 29578
rect 12164 29514 12216 29520
rect 12072 28552 12124 28558
rect 12072 28494 12124 28500
rect 11980 28484 12032 28490
rect 11980 28426 12032 28432
rect 11992 28218 12020 28426
rect 11796 28212 11848 28218
rect 11796 28154 11848 28160
rect 11980 28212 12032 28218
rect 11980 28154 12032 28160
rect 12084 28082 12112 28494
rect 12176 28082 12204 29514
rect 12532 29164 12584 29170
rect 12532 29106 12584 29112
rect 12440 29028 12492 29034
rect 12440 28970 12492 28976
rect 12452 28490 12480 28970
rect 12440 28484 12492 28490
rect 12440 28426 12492 28432
rect 12072 28076 12124 28082
rect 12072 28018 12124 28024
rect 12164 28076 12216 28082
rect 12164 28018 12216 28024
rect 12176 27946 12204 28018
rect 11704 27940 11756 27946
rect 11704 27882 11756 27888
rect 12164 27940 12216 27946
rect 12164 27882 12216 27888
rect 11612 27668 11664 27674
rect 11612 27610 11664 27616
rect 11716 27470 11744 27882
rect 11704 27464 11756 27470
rect 11704 27406 11756 27412
rect 11244 27328 11296 27334
rect 11244 27270 11296 27276
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 11164 23322 11192 24142
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 11072 22234 11100 22714
rect 11060 22228 11112 22234
rect 11060 22170 11112 22176
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 11072 21010 11100 21422
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 11072 19718 11100 20946
rect 11256 20942 11284 27270
rect 12544 27146 12572 29106
rect 12820 28762 12848 32302
rect 12624 28756 12676 28762
rect 12624 28698 12676 28704
rect 12808 28756 12860 28762
rect 12808 28698 12860 28704
rect 12636 28626 12664 28698
rect 12624 28620 12676 28626
rect 12624 28562 12676 28568
rect 12808 27872 12860 27878
rect 12808 27814 12860 27820
rect 12452 27118 12572 27146
rect 12256 26920 12308 26926
rect 12256 26862 12308 26868
rect 12268 26586 12296 26862
rect 12348 26852 12400 26858
rect 12348 26794 12400 26800
rect 12360 26586 12388 26794
rect 11980 26580 12032 26586
rect 11980 26522 12032 26528
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 12348 26580 12400 26586
rect 12348 26522 12400 26528
rect 11992 26382 12020 26522
rect 11980 26376 12032 26382
rect 12256 26376 12308 26382
rect 11980 26318 12032 26324
rect 12084 26324 12256 26330
rect 12084 26318 12308 26324
rect 12084 26314 12296 26318
rect 12072 26308 12296 26314
rect 12124 26302 12296 26308
rect 12072 26250 12124 26256
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 11888 25152 11940 25158
rect 11888 25094 11940 25100
rect 11428 24744 11480 24750
rect 11624 24698 11652 25094
rect 11900 24818 11928 25094
rect 11888 24812 11940 24818
rect 11888 24754 11940 24760
rect 11480 24692 11652 24698
rect 11428 24686 11652 24692
rect 11440 24670 11652 24686
rect 11520 24200 11572 24206
rect 11520 24142 11572 24148
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11348 23798 11376 24006
rect 11336 23792 11388 23798
rect 11336 23734 11388 23740
rect 11532 23662 11560 24142
rect 11520 23656 11572 23662
rect 11520 23598 11572 23604
rect 11532 23254 11560 23598
rect 11428 23248 11480 23254
rect 11428 23190 11480 23196
rect 11520 23248 11572 23254
rect 11520 23190 11572 23196
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 11256 20602 11284 20878
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 10980 17746 11008 18634
rect 10968 17740 11020 17746
rect 10968 17682 11020 17688
rect 10980 16726 11008 17682
rect 11072 17270 11100 19314
rect 11164 18902 11192 19858
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 11164 16250 11192 16730
rect 11440 16590 11468 23190
rect 11532 22098 11560 23190
rect 11624 22098 11652 24670
rect 11704 24268 11756 24274
rect 11704 24210 11756 24216
rect 11716 23186 11744 24210
rect 11900 23798 11928 24754
rect 11888 23792 11940 23798
rect 11888 23734 11940 23740
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 11520 22092 11572 22098
rect 11520 22034 11572 22040
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11532 21554 11560 22034
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11716 21146 11744 23122
rect 11704 21140 11756 21146
rect 11704 21082 11756 21088
rect 11612 20800 11664 20806
rect 11612 20742 11664 20748
rect 11624 20602 11652 20742
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11992 20058 12020 20402
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11532 19378 11560 19790
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11532 18290 11560 19314
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11624 18358 11652 18566
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11440 15366 11468 16390
rect 11532 16182 11560 18226
rect 11808 17882 11836 18702
rect 11796 17876 11848 17882
rect 11796 17818 11848 17824
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11808 17134 11836 17478
rect 11796 17128 11848 17134
rect 11796 17070 11848 17076
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11808 16590 11836 16934
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11520 16176 11572 16182
rect 11520 16118 11572 16124
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 11992 15502 12020 16118
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11072 15162 11100 15302
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 11440 14958 11468 15302
rect 11428 14952 11480 14958
rect 11428 14894 11480 14900
rect 12084 14074 12112 26250
rect 12452 26042 12480 27118
rect 12820 27062 12848 27814
rect 12808 27056 12860 27062
rect 12808 26998 12860 27004
rect 12820 26858 12848 26998
rect 12808 26852 12860 26858
rect 12808 26794 12860 26800
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12912 25498 12940 32846
rect 13004 32026 13032 32914
rect 13188 32434 13216 33322
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 13280 32366 13308 33458
rect 14096 33312 14148 33318
rect 14096 33254 14148 33260
rect 13820 32768 13872 32774
rect 13820 32710 13872 32716
rect 13832 32434 13860 32710
rect 14108 32434 14136 33254
rect 14292 32910 14320 33526
rect 16212 33516 16264 33522
rect 16212 33458 16264 33464
rect 22192 33516 22244 33522
rect 22192 33458 22244 33464
rect 25964 33516 26016 33522
rect 25964 33458 26016 33464
rect 16028 33312 16080 33318
rect 16028 33254 16080 33260
rect 14280 32904 14332 32910
rect 14280 32846 14332 32852
rect 14464 32904 14516 32910
rect 14464 32846 14516 32852
rect 15016 32904 15068 32910
rect 15016 32846 15068 32852
rect 14476 32434 14504 32846
rect 15028 32774 15056 32846
rect 16040 32842 16068 33254
rect 16224 33114 16252 33458
rect 16212 33108 16264 33114
rect 16212 33050 16264 33056
rect 19340 33040 19392 33046
rect 19340 32982 19392 32988
rect 19352 32910 19380 32982
rect 22204 32910 22232 33458
rect 23664 33448 23716 33454
rect 23664 33390 23716 33396
rect 16396 32904 16448 32910
rect 16396 32846 16448 32852
rect 19340 32904 19392 32910
rect 19340 32846 19392 32852
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 16028 32836 16080 32842
rect 16028 32778 16080 32784
rect 15016 32768 15068 32774
rect 15016 32710 15068 32716
rect 13820 32428 13872 32434
rect 13820 32370 13872 32376
rect 14096 32428 14148 32434
rect 14096 32370 14148 32376
rect 14464 32428 14516 32434
rect 14464 32370 14516 32376
rect 13268 32360 13320 32366
rect 13268 32302 13320 32308
rect 14280 32224 14332 32230
rect 14280 32166 14332 32172
rect 12992 32020 13044 32026
rect 12992 31962 13044 31968
rect 13636 32020 13688 32026
rect 13636 31962 13688 31968
rect 13648 31822 13676 31962
rect 13636 31816 13688 31822
rect 13636 31758 13688 31764
rect 13648 31482 13676 31758
rect 13636 31476 13688 31482
rect 13636 31418 13688 31424
rect 13728 31272 13780 31278
rect 13728 31214 13780 31220
rect 13820 31272 13872 31278
rect 13820 31214 13872 31220
rect 13740 30666 13768 31214
rect 13728 30660 13780 30666
rect 13728 30602 13780 30608
rect 13832 30122 13860 31214
rect 14188 31136 14240 31142
rect 14188 31078 14240 31084
rect 13820 30116 13872 30122
rect 13820 30058 13872 30064
rect 13832 29714 13860 30058
rect 13820 29708 13872 29714
rect 13820 29650 13872 29656
rect 13544 28552 13596 28558
rect 13544 28494 13596 28500
rect 12992 28076 13044 28082
rect 12992 28018 13044 28024
rect 13004 27334 13032 28018
rect 13556 27878 13584 28494
rect 13544 27872 13596 27878
rect 13544 27814 13596 27820
rect 12992 27328 13044 27334
rect 12992 27270 13044 27276
rect 13004 26586 13032 27270
rect 13176 26988 13228 26994
rect 13176 26930 13228 26936
rect 12992 26580 13044 26586
rect 12992 26522 13044 26528
rect 13188 26314 13216 26930
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 13176 26308 13228 26314
rect 13176 26250 13228 26256
rect 12900 25492 12952 25498
rect 12900 25434 12952 25440
rect 12912 24886 12940 25434
rect 13096 25242 13124 26250
rect 13176 25900 13228 25906
rect 13176 25842 13228 25848
rect 13188 25430 13216 25842
rect 13176 25424 13228 25430
rect 13176 25366 13228 25372
rect 13096 25214 13216 25242
rect 12900 24880 12952 24886
rect 12900 24822 12952 24828
rect 12808 24812 12860 24818
rect 12808 24754 12860 24760
rect 12820 24410 12848 24754
rect 12900 24744 12952 24750
rect 12900 24686 12952 24692
rect 12808 24404 12860 24410
rect 12808 24346 12860 24352
rect 12912 23866 12940 24686
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12452 22642 12480 22918
rect 12544 22778 12572 23666
rect 12912 23050 12940 23802
rect 12900 23044 12952 23050
rect 12900 22986 12952 22992
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12912 22642 12940 22986
rect 13096 22710 13124 24550
rect 13084 22704 13136 22710
rect 13084 22646 13136 22652
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 13188 22094 13216 25214
rect 13360 24132 13412 24138
rect 13360 24074 13412 24080
rect 13372 23866 13400 24074
rect 13360 23860 13412 23866
rect 13360 23802 13412 23808
rect 13188 22066 13400 22094
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12544 21486 12572 21966
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12176 20058 12204 20334
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 12268 19922 12296 20946
rect 12544 20942 12572 21422
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12360 19854 12388 20538
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12544 17610 12572 18090
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12360 17134 12388 17478
rect 12544 17202 12572 17546
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12176 15978 12204 16390
rect 12164 15972 12216 15978
rect 12164 15914 12216 15920
rect 12360 15162 12388 17070
rect 12636 17066 12664 17206
rect 12728 17202 12756 18566
rect 12912 18222 12940 18838
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12912 18086 12940 18158
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12912 17678 12940 18022
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 13372 17542 13400 22066
rect 13556 20874 13584 27814
rect 13832 26790 13860 29650
rect 13912 29504 13964 29510
rect 13912 29446 13964 29452
rect 13924 27010 13952 29446
rect 14004 29300 14056 29306
rect 14004 29242 14056 29248
rect 14016 28558 14044 29242
rect 14096 28756 14148 28762
rect 14096 28698 14148 28704
rect 14004 28552 14056 28558
rect 14004 28494 14056 28500
rect 14108 27130 14136 28698
rect 14200 28626 14228 31078
rect 14292 29102 14320 32166
rect 14476 32026 14504 32370
rect 14740 32360 14792 32366
rect 14740 32302 14792 32308
rect 14464 32020 14516 32026
rect 14464 31962 14516 31968
rect 14556 29300 14608 29306
rect 14556 29242 14608 29248
rect 14280 29096 14332 29102
rect 14280 29038 14332 29044
rect 14188 28620 14240 28626
rect 14188 28562 14240 28568
rect 14292 28150 14320 29038
rect 14568 28762 14596 29242
rect 14556 28756 14608 28762
rect 14556 28698 14608 28704
rect 14752 28626 14780 32302
rect 14924 31272 14976 31278
rect 14924 31214 14976 31220
rect 14936 31142 14964 31214
rect 14924 31136 14976 31142
rect 14922 31104 14924 31113
rect 14976 31104 14978 31113
rect 14922 31039 14978 31048
rect 14740 28620 14792 28626
rect 14740 28562 14792 28568
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14384 28218 14412 28494
rect 14372 28212 14424 28218
rect 14372 28154 14424 28160
rect 14280 28144 14332 28150
rect 14280 28086 14332 28092
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14096 27124 14148 27130
rect 14096 27066 14148 27072
rect 13924 26982 14228 27010
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 14004 26784 14056 26790
rect 14004 26726 14056 26732
rect 13636 26308 13688 26314
rect 13636 26250 13688 26256
rect 13820 26308 13872 26314
rect 13820 26250 13872 26256
rect 13544 20868 13596 20874
rect 13544 20810 13596 20816
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13556 18154 13584 18566
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12636 16794 12664 17002
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12440 16720 12492 16726
rect 12440 16662 12492 16668
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12452 14890 12480 16662
rect 12808 16176 12860 16182
rect 12808 16118 12860 16124
rect 12532 15428 12584 15434
rect 12532 15370 12584 15376
rect 12544 15162 12572 15370
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12440 14884 12492 14890
rect 12440 14826 12492 14832
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12544 14618 12572 14758
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9508 11558 9536 12038
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 9508 10130 9536 10950
rect 9600 10810 9628 10950
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8312 9450 8340 9930
rect 8956 9722 8984 10066
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8116 9104 8168 9110
rect 8116 9046 8168 9052
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7478 7880 7686
rect 7840 7472 7892 7478
rect 7840 7414 7892 7420
rect 7944 7410 7972 8366
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 7196 7404 7248 7410
rect 7196 7346 7248 7352
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7208 7002 7236 7346
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7944 6866 7972 7346
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7668 6390 7696 6598
rect 8312 6458 8340 8026
rect 8404 6798 8432 9658
rect 9048 9654 9076 9998
rect 9036 9648 9088 9654
rect 9036 9590 9088 9596
rect 9048 8634 9076 9590
rect 9140 9450 9168 9998
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9232 7546 9260 7822
rect 9324 7546 9352 9522
rect 9784 9042 9812 13670
rect 10612 12850 10640 13738
rect 11704 13728 11756 13734
rect 11704 13670 11756 13676
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11428 13252 11480 13258
rect 11428 13194 11480 13200
rect 11440 12986 11468 13194
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10428 12442 10456 12786
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10428 11898 10456 12174
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 11072 11694 11100 12038
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 11060 11688 11112 11694
rect 11060 11630 11112 11636
rect 10704 9518 10732 11630
rect 11072 11121 11100 11630
rect 11256 11354 11284 11698
rect 11532 11694 11560 13262
rect 11716 12850 11744 13670
rect 12084 13530 12112 14010
rect 12544 14006 12572 14554
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 12636 12714 12664 13738
rect 12820 13258 12848 16118
rect 13452 15088 13504 15094
rect 13452 15030 13504 15036
rect 13464 14618 13492 15030
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12716 12912 12768 12918
rect 12716 12854 12768 12860
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12728 12442 12756 12854
rect 12820 12442 12848 13194
rect 13084 12708 13136 12714
rect 13084 12650 13136 12656
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12808 12436 12860 12442
rect 12808 12378 12860 12384
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11992 11830 12020 12038
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11058 11112 11114 11121
rect 11058 11047 11114 11056
rect 11532 10606 11560 11630
rect 12268 11354 12296 12174
rect 12624 11620 12676 11626
rect 12624 11562 12676 11568
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12636 11150 12664 11562
rect 13096 11218 13124 12650
rect 13464 12434 13492 14554
rect 13464 12406 13584 12434
rect 13452 11280 13504 11286
rect 13452 11222 13504 11228
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 10692 9512 10744 9518
rect 10692 9454 10744 9460
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9600 8090 9628 8366
rect 9692 8362 9720 8910
rect 9784 8566 9812 8978
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9968 8090 9996 8842
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10796 8242 10824 8298
rect 10796 8214 10916 8242
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10888 7818 10916 8214
rect 10980 8022 11008 9454
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10888 7546 10916 7754
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 9324 6730 9352 7278
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9324 6458 9352 6666
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6380 5370 6408 5578
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6932 5234 6960 6054
rect 7668 5914 7696 6326
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 8312 5846 8340 6394
rect 10060 6322 10088 6598
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 9508 5710 9536 6054
rect 10336 5710 10364 6598
rect 10428 6254 10456 6802
rect 10520 6458 10548 7210
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10980 6458 11008 6734
rect 10508 6452 10560 6458
rect 10508 6394 10560 6400
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 9140 5234 9168 5646
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5234 9444 5510
rect 10520 5370 10548 6394
rect 11440 6390 11468 7822
rect 11532 6390 11560 10542
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11428 6384 11480 6390
rect 11428 6326 11480 6332
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11072 5778 11100 6190
rect 11440 5846 11468 6326
rect 11532 6254 11560 6326
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11520 6248 11572 6254
rect 11520 6190 11572 6196
rect 11532 5914 11560 6190
rect 11624 5914 11652 6258
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 9876 4758 9904 5170
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10428 4758 10456 5034
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 8666 4176 8722 4185
rect 8666 4111 8668 4120
rect 8720 4111 8722 4120
rect 8668 4082 8720 4088
rect 8116 3936 8168 3942
rect 10324 3936 10376 3942
rect 8116 3878 8168 3884
rect 10322 3904 10324 3913
rect 10376 3904 10378 3913
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 8128 3534 8156 3878
rect 10322 3839 10378 3848
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8390 3496 8446 3505
rect 8390 3431 8392 3440
rect 8444 3431 8446 3440
rect 10692 3460 10744 3466
rect 8392 3402 8444 3408
rect 10692 3402 10744 3408
rect 11336 3460 11388 3466
rect 11336 3402 11388 3408
rect 9956 3392 10008 3398
rect 8482 3360 8538 3369
rect 9956 3334 10008 3340
rect 8482 3295 8538 3304
rect 8496 3126 8524 3295
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 9680 2440 9732 2446
rect 9968 2417 9996 3334
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10244 3058 10272 3130
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10152 2825 10180 2994
rect 10138 2816 10194 2825
rect 10138 2751 10194 2760
rect 10324 2440 10376 2446
rect 9680 2382 9732 2388
rect 9954 2408 10010 2417
rect 8220 2106 8248 2382
rect 8208 2100 8260 2106
rect 8208 2042 8260 2048
rect 9692 2038 9720 2382
rect 10324 2382 10376 2388
rect 9954 2343 10010 2352
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 10336 1970 10364 2382
rect 10324 1964 10376 1970
rect 10324 1906 10376 1912
rect 10704 1698 10732 3402
rect 10874 3088 10930 3097
rect 10874 3023 10930 3032
rect 10888 2854 10916 3023
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10980 2650 11008 2926
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11348 2582 11376 3402
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 10692 1692 10744 1698
rect 10692 1634 10744 1640
rect 10980 1465 11008 2382
rect 11440 1766 11468 4558
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11624 3738 11652 4490
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11428 1760 11480 1766
rect 11428 1702 11480 1708
rect 10966 1456 11022 1465
rect 10966 1391 11022 1400
rect 11624 1222 11652 3538
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 11716 1834 11744 2314
rect 11704 1828 11756 1834
rect 11704 1770 11756 1776
rect 11612 1216 11664 1222
rect 11612 1158 11664 1164
rect 11808 762 11836 10406
rect 12176 10266 12204 10610
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12912 10062 12940 10678
rect 13096 10130 13124 11154
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11992 7478 12020 8502
rect 12268 8430 12296 8774
rect 12348 8492 12400 8498
rect 12348 8434 12400 8440
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11900 2009 11928 3470
rect 11992 2378 12020 7142
rect 12360 6798 12388 8434
rect 12728 8430 12756 9522
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12636 7274 12664 7822
rect 12624 7268 12676 7274
rect 12624 7210 12676 7216
rect 13096 6866 13124 10066
rect 13464 9586 13492 11222
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13280 8022 13308 9454
rect 13556 8401 13584 12406
rect 13648 9450 13676 26250
rect 13832 25770 13860 26250
rect 13820 25764 13872 25770
rect 13820 25706 13872 25712
rect 13728 24880 13780 24886
rect 13728 24822 13780 24828
rect 13740 22982 13768 24822
rect 13832 24070 13860 25706
rect 14016 25498 14044 26726
rect 14096 25900 14148 25906
rect 14096 25842 14148 25848
rect 14004 25492 14056 25498
rect 14004 25434 14056 25440
rect 14108 25158 14136 25842
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 13924 24206 13952 24686
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13832 23050 13860 24006
rect 13924 23118 13952 24142
rect 14108 23866 14136 25094
rect 14096 23860 14148 23866
rect 14096 23802 14148 23808
rect 14004 23724 14056 23730
rect 14004 23666 14056 23672
rect 14016 23322 14044 23666
rect 14004 23316 14056 23322
rect 14004 23258 14056 23264
rect 14108 23186 14136 23802
rect 14096 23180 14148 23186
rect 14096 23122 14148 23128
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 13820 23044 13872 23050
rect 13820 22986 13872 22992
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13820 22092 13872 22098
rect 13820 22034 13872 22040
rect 13728 15360 13780 15366
rect 13728 15302 13780 15308
rect 13740 12986 13768 15302
rect 13832 14006 13860 22034
rect 13924 21010 13952 23054
rect 14200 22642 14228 26982
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14292 26518 14320 26726
rect 14280 26512 14332 26518
rect 14280 26454 14332 26460
rect 14292 25838 14320 26454
rect 14752 25838 14780 27406
rect 14280 25832 14332 25838
rect 14280 25774 14332 25780
rect 14740 25832 14792 25838
rect 14740 25774 14792 25780
rect 14188 22636 14240 22642
rect 14188 22578 14240 22584
rect 14004 22500 14056 22506
rect 14004 22442 14056 22448
rect 14016 22166 14044 22442
rect 14004 22160 14056 22166
rect 14004 22102 14056 22108
rect 13912 21004 13964 21010
rect 13912 20946 13964 20952
rect 14016 20602 14044 22102
rect 14200 21894 14228 22578
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14200 20913 14228 21830
rect 14292 21146 14320 25774
rect 14924 25696 14976 25702
rect 14924 25638 14976 25644
rect 14464 25220 14516 25226
rect 14464 25162 14516 25168
rect 14476 23186 14504 25162
rect 14936 24614 14964 25638
rect 14924 24608 14976 24614
rect 14924 24550 14976 24556
rect 14936 24274 14964 24550
rect 14924 24268 14976 24274
rect 14924 24210 14976 24216
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14464 23180 14516 23186
rect 14464 23122 14516 23128
rect 14476 22094 14504 23122
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 22710 14596 22918
rect 14660 22778 14688 24142
rect 15028 24138 15056 32710
rect 16040 32434 16068 32778
rect 15476 32428 15528 32434
rect 15476 32370 15528 32376
rect 16028 32428 16080 32434
rect 16028 32370 16080 32376
rect 15292 32224 15344 32230
rect 15292 32166 15344 32172
rect 15304 31754 15332 32166
rect 15292 31748 15344 31754
rect 15292 31690 15344 31696
rect 15384 31748 15436 31754
rect 15384 31690 15436 31696
rect 15396 29646 15424 31690
rect 15488 31482 15516 32370
rect 16408 32026 16436 32846
rect 18236 32768 18288 32774
rect 18236 32710 18288 32716
rect 18248 32570 18276 32710
rect 18236 32564 18288 32570
rect 18236 32506 18288 32512
rect 18696 32428 18748 32434
rect 18696 32370 18748 32376
rect 17408 32360 17460 32366
rect 17408 32302 17460 32308
rect 16396 32020 16448 32026
rect 16396 31962 16448 31968
rect 16408 31482 16436 31962
rect 16580 31952 16632 31958
rect 16580 31894 16632 31900
rect 15476 31476 15528 31482
rect 15476 31418 15528 31424
rect 16396 31476 16448 31482
rect 16396 31418 16448 31424
rect 16592 30938 16620 31894
rect 17420 31482 17448 32302
rect 17592 32224 17644 32230
rect 17592 32166 17644 32172
rect 17604 31754 17632 32166
rect 18144 31816 18196 31822
rect 18144 31758 18196 31764
rect 17592 31748 17644 31754
rect 17592 31690 17644 31696
rect 17224 31476 17276 31482
rect 17224 31418 17276 31424
rect 17408 31476 17460 31482
rect 17408 31418 17460 31424
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 16948 31204 17000 31210
rect 16948 31146 17000 31152
rect 15936 30932 15988 30938
rect 15936 30874 15988 30880
rect 16580 30932 16632 30938
rect 16580 30874 16632 30880
rect 15476 30728 15528 30734
rect 15476 30670 15528 30676
rect 15488 30394 15516 30670
rect 15568 30592 15620 30598
rect 15568 30534 15620 30540
rect 15476 30388 15528 30394
rect 15476 30330 15528 30336
rect 15580 29646 15608 30534
rect 15844 30184 15896 30190
rect 15844 30126 15896 30132
rect 15384 29640 15436 29646
rect 15384 29582 15436 29588
rect 15568 29640 15620 29646
rect 15568 29582 15620 29588
rect 15108 29504 15160 29510
rect 15108 29446 15160 29452
rect 15120 29170 15148 29446
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 15120 28540 15148 29106
rect 15200 28552 15252 28558
rect 15120 28512 15200 28540
rect 15200 28494 15252 28500
rect 15212 28218 15240 28494
rect 15200 28212 15252 28218
rect 15120 28172 15200 28200
rect 15120 27538 15148 28172
rect 15200 28154 15252 28160
rect 15292 28076 15344 28082
rect 15212 28036 15292 28064
rect 15108 27532 15160 27538
rect 15108 27474 15160 27480
rect 15212 27470 15240 28036
rect 15292 28018 15344 28024
rect 15200 27464 15252 27470
rect 15200 27406 15252 27412
rect 15212 26586 15240 27406
rect 15200 26580 15252 26586
rect 15200 26522 15252 26528
rect 15396 26450 15424 29582
rect 15856 29170 15884 30126
rect 15948 29238 15976 30874
rect 16960 30666 16988 31146
rect 16948 30660 17000 30666
rect 16948 30602 17000 30608
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 16684 29850 16712 30194
rect 16960 30054 16988 30602
rect 17052 30326 17080 31282
rect 17132 31272 17184 31278
rect 17132 31214 17184 31220
rect 17144 30802 17172 31214
rect 17132 30796 17184 30802
rect 17132 30738 17184 30744
rect 17040 30320 17092 30326
rect 17040 30262 17092 30268
rect 16948 30048 17000 30054
rect 16948 29990 17000 29996
rect 16672 29844 16724 29850
rect 16672 29786 16724 29792
rect 16684 29646 16712 29786
rect 16672 29640 16724 29646
rect 16672 29582 16724 29588
rect 15936 29232 15988 29238
rect 15936 29174 15988 29180
rect 15844 29164 15896 29170
rect 15844 29106 15896 29112
rect 15568 27940 15620 27946
rect 15568 27882 15620 27888
rect 15580 27334 15608 27882
rect 15568 27328 15620 27334
rect 15568 27270 15620 27276
rect 15568 26784 15620 26790
rect 15568 26726 15620 26732
rect 15384 26444 15436 26450
rect 15384 26386 15436 26392
rect 15396 26042 15424 26386
rect 15580 26246 15608 26726
rect 15660 26308 15712 26314
rect 15660 26250 15712 26256
rect 15568 26240 15620 26246
rect 15568 26182 15620 26188
rect 15384 26036 15436 26042
rect 15384 25978 15436 25984
rect 15580 25906 15608 26182
rect 15672 26042 15700 26250
rect 15660 26036 15712 26042
rect 15660 25978 15712 25984
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15948 25650 15976 29174
rect 16684 29170 16712 29582
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16672 28960 16724 28966
rect 16672 28902 16724 28908
rect 16684 28694 16712 28902
rect 16672 28688 16724 28694
rect 16672 28630 16724 28636
rect 16762 28656 16818 28665
rect 16762 28591 16818 28600
rect 16776 28558 16804 28591
rect 16764 28552 16816 28558
rect 16764 28494 16816 28500
rect 16580 25900 16632 25906
rect 16580 25842 16632 25848
rect 16488 25832 16540 25838
rect 16488 25774 16540 25780
rect 15856 25622 15976 25650
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15304 24614 15332 25094
rect 15292 24608 15344 24614
rect 15292 24550 15344 24556
rect 15304 24342 15332 24550
rect 15292 24336 15344 24342
rect 15292 24278 15344 24284
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 15200 23724 15252 23730
rect 15200 23666 15252 23672
rect 14648 22772 14700 22778
rect 14648 22714 14700 22720
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14476 22066 14596 22094
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14186 20904 14242 20913
rect 14186 20839 14242 20848
rect 14188 20800 14240 20806
rect 14188 20742 14240 20748
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 14200 20534 14228 20742
rect 14188 20528 14240 20534
rect 14188 20470 14240 20476
rect 14200 19990 14228 20470
rect 14188 19984 14240 19990
rect 14188 19926 14240 19932
rect 14476 19922 14504 20946
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14188 17536 14240 17542
rect 14186 17504 14188 17513
rect 14240 17504 14242 17513
rect 14186 17439 14242 17448
rect 14096 15904 14148 15910
rect 14096 15846 14148 15852
rect 14108 15026 14136 15846
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13832 12918 13860 13942
rect 14108 13258 14136 14962
rect 14476 14906 14504 14962
rect 14384 14878 14504 14906
rect 14384 14414 14412 14878
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14384 13938 14412 14350
rect 14372 13932 14424 13938
rect 14372 13874 14424 13880
rect 14096 13252 14148 13258
rect 14096 13194 14148 13200
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 14108 12850 14136 13194
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 14108 12434 14136 12786
rect 14108 12406 14320 12434
rect 13728 10804 13780 10810
rect 13728 10746 13780 10752
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13740 9382 13768 10746
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14108 8634 14136 9046
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 13542 8392 13598 8401
rect 13542 8327 13598 8336
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13268 8016 13320 8022
rect 13268 7958 13320 7964
rect 13740 7954 13768 8298
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 13912 7200 13964 7206
rect 13912 7142 13964 7148
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13924 6798 13952 7142
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 12072 6656 12124 6662
rect 12072 6598 12124 6604
rect 12084 5710 12112 6598
rect 12360 6458 12388 6734
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12164 6112 12216 6118
rect 12164 6054 12216 6060
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12072 5160 12124 5166
rect 12072 5102 12124 5108
rect 12084 4622 12112 5102
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12084 4282 12112 4558
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12176 3738 12204 6054
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12254 5128 12310 5137
rect 12452 5098 12480 5646
rect 12820 5642 12848 6598
rect 13648 6322 13676 6598
rect 14016 6390 14044 6666
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 14108 5710 14136 7210
rect 13268 5704 13320 5710
rect 14096 5704 14148 5710
rect 13268 5646 13320 5652
rect 13924 5664 14096 5692
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12254 5063 12310 5072
rect 12440 5092 12492 5098
rect 12268 4486 12296 5063
rect 12440 5034 12492 5040
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12072 3528 12124 3534
rect 12070 3496 12072 3505
rect 12124 3496 12126 3505
rect 12126 3454 12204 3482
rect 12070 3431 12126 3440
rect 12072 2984 12124 2990
rect 12070 2952 12072 2961
rect 12124 2952 12126 2961
rect 12070 2887 12126 2896
rect 11980 2372 12032 2378
rect 11980 2314 12032 2320
rect 11886 2000 11942 2009
rect 11886 1935 11942 1944
rect 12176 1902 12204 3454
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12268 2990 12296 3334
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12360 2582 12388 4966
rect 12452 2666 12480 5034
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12636 3398 12664 4966
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12728 4622 12756 4762
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12820 4468 12848 5578
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12728 4440 12848 4468
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12728 3194 12756 4440
rect 12806 4176 12862 4185
rect 12806 4111 12808 4120
rect 12860 4111 12862 4120
rect 12808 4082 12860 4088
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12820 3738 12848 3946
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12912 3534 12940 5510
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 12714 2680 12770 2689
rect 12452 2638 12664 2666
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12164 1896 12216 1902
rect 12164 1838 12216 1844
rect 12268 870 12388 898
rect 12268 762 12296 870
rect 12360 800 12388 870
rect 12452 800 12480 2450
rect 12544 800 12572 2518
rect 12636 800 12664 2638
rect 12714 2615 12770 2624
rect 12728 2514 12756 2615
rect 12716 2508 12768 2514
rect 12716 2450 12768 2456
rect 12716 2100 12768 2106
rect 12716 2042 12768 2048
rect 12728 800 12756 2042
rect 12992 1828 13044 1834
rect 12992 1770 13044 1776
rect 12900 1760 12952 1766
rect 12900 1702 12952 1708
rect 12808 1692 12860 1698
rect 12808 1634 12860 1640
rect 12820 800 12848 1634
rect 12912 800 12940 1702
rect 13004 800 13032 1770
rect 13096 800 13124 2790
rect 13188 800 13216 5170
rect 13280 4690 13308 5646
rect 13360 5160 13412 5166
rect 13360 5102 13412 5108
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13280 800 13308 4626
rect 13372 3534 13400 5102
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13464 4010 13492 4558
rect 13728 4208 13780 4214
rect 13728 4150 13780 4156
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13372 800 13400 2994
rect 13464 800 13492 3674
rect 13556 2553 13584 4082
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13542 2544 13598 2553
rect 13542 2479 13598 2488
rect 13648 800 13676 3470
rect 13740 800 13768 4150
rect 13832 800 13860 4966
rect 13924 3482 13952 5664
rect 14096 5646 14148 5652
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14016 3602 14044 5510
rect 14004 3596 14056 3602
rect 14004 3538 14056 3544
rect 14108 3534 14136 5510
rect 14188 4752 14240 4758
rect 14188 4694 14240 4700
rect 14292 4706 14320 12406
rect 14384 4826 14412 13874
rect 14568 13326 14596 22066
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 14740 21344 14792 21350
rect 14740 21286 14792 21292
rect 14752 20942 14780 21286
rect 14740 20936 14792 20942
rect 15016 20936 15068 20942
rect 14740 20878 14792 20884
rect 15014 20904 15016 20913
rect 15068 20904 15070 20913
rect 15014 20839 15070 20848
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14844 19854 14872 20198
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 19446 14688 19654
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 15120 17610 15148 21830
rect 15212 20534 15240 23666
rect 15396 22166 15424 25094
rect 15660 24064 15712 24070
rect 15660 24006 15712 24012
rect 15672 23118 15700 24006
rect 15856 23730 15884 25622
rect 16500 25362 16528 25774
rect 16488 25356 16540 25362
rect 16488 25298 16540 25304
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15948 24818 15976 25094
rect 16500 24954 16528 25298
rect 16488 24948 16540 24954
rect 16488 24890 16540 24896
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 16120 24200 16172 24206
rect 16120 24142 16172 24148
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 16132 23594 16160 24142
rect 16396 24132 16448 24138
rect 16396 24074 16448 24080
rect 16408 23594 16436 24074
rect 16120 23588 16172 23594
rect 16120 23530 16172 23536
rect 16396 23588 16448 23594
rect 16396 23530 16448 23536
rect 16500 23526 16528 24890
rect 16592 24410 16620 25842
rect 16868 25498 16896 29106
rect 16856 25492 16908 25498
rect 16856 25434 16908 25440
rect 16868 25294 16896 25434
rect 16856 25288 16908 25294
rect 16856 25230 16908 25236
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16764 24608 16816 24614
rect 16764 24550 16816 24556
rect 16580 24404 16632 24410
rect 16580 24346 16632 24352
rect 16776 24206 16804 24550
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 16500 22166 16528 23462
rect 16776 23322 16804 23598
rect 16764 23316 16816 23322
rect 16764 23258 16816 23264
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 16776 22166 16804 22714
rect 15384 22160 15436 22166
rect 15384 22102 15436 22108
rect 16488 22160 16540 22166
rect 16488 22102 16540 22108
rect 16764 22160 16816 22166
rect 16764 22102 16816 22108
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15200 20528 15252 20534
rect 15200 20470 15252 20476
rect 15304 20330 15332 21490
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 15396 18426 15424 22102
rect 16776 21978 16804 22102
rect 16868 22030 16896 25094
rect 16960 22094 16988 29990
rect 17038 28520 17094 28529
rect 17038 28455 17040 28464
rect 17092 28455 17094 28464
rect 17040 28426 17092 28432
rect 17132 28416 17184 28422
rect 17132 28358 17184 28364
rect 17144 27878 17172 28358
rect 17132 27872 17184 27878
rect 17132 27814 17184 27820
rect 17040 27396 17092 27402
rect 17040 27338 17092 27344
rect 17052 27062 17080 27338
rect 17040 27056 17092 27062
rect 17040 26998 17092 27004
rect 17132 26988 17184 26994
rect 17132 26930 17184 26936
rect 17144 26042 17172 26930
rect 17132 26036 17184 26042
rect 17132 25978 17184 25984
rect 17040 25968 17092 25974
rect 17040 25910 17092 25916
rect 17052 24886 17080 25910
rect 17040 24880 17092 24886
rect 17040 24822 17092 24828
rect 17052 22658 17080 24822
rect 17236 24818 17264 31418
rect 18156 31362 18184 31758
rect 18156 31346 18276 31362
rect 18156 31340 18288 31346
rect 18156 31334 18236 31340
rect 18236 31282 18288 31288
rect 18420 31340 18472 31346
rect 18420 31282 18472 31288
rect 17316 31136 17368 31142
rect 17316 31078 17368 31084
rect 17328 30734 17356 31078
rect 17960 30864 18012 30870
rect 17960 30806 18012 30812
rect 17316 30728 17368 30734
rect 17316 30670 17368 30676
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17316 27396 17368 27402
rect 17316 27338 17368 27344
rect 17328 27130 17356 27338
rect 17316 27124 17368 27130
rect 17316 27066 17368 27072
rect 17512 27010 17540 28358
rect 17684 27872 17736 27878
rect 17684 27814 17736 27820
rect 17328 26982 17540 27010
rect 17224 24812 17276 24818
rect 17224 24754 17276 24760
rect 17132 23792 17184 23798
rect 17132 23734 17184 23740
rect 17144 22778 17172 23734
rect 17236 23730 17264 24754
rect 17224 23724 17276 23730
rect 17224 23666 17276 23672
rect 17236 22778 17264 23666
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17224 22772 17276 22778
rect 17224 22714 17276 22720
rect 17052 22630 17172 22658
rect 16960 22066 17080 22094
rect 16592 21950 16804 21978
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16948 21956 17000 21962
rect 16028 20868 16080 20874
rect 16028 20810 16080 20816
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15856 20534 15884 20742
rect 15844 20528 15896 20534
rect 15844 20470 15896 20476
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15488 19718 15516 20402
rect 15844 20392 15896 20398
rect 15844 20334 15896 20340
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15488 19514 15516 19654
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15856 18340 15884 20334
rect 15936 19780 15988 19786
rect 15936 19722 15988 19728
rect 15948 19514 15976 19722
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15856 18312 15976 18340
rect 15948 18222 15976 18312
rect 15936 18216 15988 18222
rect 15936 18158 15988 18164
rect 15752 18148 15804 18154
rect 15752 18090 15804 18096
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15108 17604 15160 17610
rect 15108 17546 15160 17552
rect 15292 17604 15344 17610
rect 15292 17546 15344 17552
rect 15120 16250 15148 17546
rect 15304 17338 15332 17546
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15396 17202 15424 18022
rect 15764 17678 15792 18090
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15764 16590 15792 17614
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15108 16244 15160 16250
rect 15108 16186 15160 16192
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15304 15502 15332 15846
rect 15764 15706 15792 16526
rect 15948 16046 15976 18158
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14752 13870 14780 14894
rect 15200 14272 15252 14278
rect 15200 14214 15252 14220
rect 15212 14074 15240 14214
rect 15200 14068 15252 14074
rect 15252 14028 15332 14056
rect 15200 14010 15252 14016
rect 14922 13968 14978 13977
rect 14922 13903 14924 13912
rect 14976 13903 14978 13912
rect 14924 13874 14976 13880
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14752 13530 14780 13806
rect 14740 13524 14792 13530
rect 14936 13512 14964 13874
rect 14936 13484 15056 13512
rect 14740 13466 14792 13472
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14752 12434 14780 13466
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14660 12406 14780 12434
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14464 7336 14516 7342
rect 14464 7278 14516 7284
rect 14476 6730 14504 7278
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14568 5574 14596 9862
rect 14660 7954 14688 12406
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14752 11218 14780 11494
rect 14844 11354 14872 12038
rect 14936 11626 14964 12582
rect 15028 12170 15056 13484
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 12374 15240 12786
rect 15304 12782 15332 14028
rect 15488 13870 15516 14962
rect 15764 14482 15792 15642
rect 15948 15094 15976 15982
rect 15936 15088 15988 15094
rect 15936 15030 15988 15036
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 15764 12918 15792 13262
rect 15752 12912 15804 12918
rect 15752 12854 15804 12860
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15016 12164 15068 12170
rect 15016 12106 15068 12112
rect 15292 12164 15344 12170
rect 15292 12106 15344 12112
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 15304 11558 15332 12106
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14752 8974 14780 9386
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14752 8650 14780 8910
rect 14752 8622 14872 8650
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14660 7342 14688 7890
rect 14752 7818 14780 8434
rect 14844 8090 14872 8622
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14936 7886 14964 8910
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14752 7478 14780 7754
rect 14740 7472 14792 7478
rect 14740 7414 14792 7420
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14752 6458 14780 7414
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 15212 6361 15240 6666
rect 15198 6352 15254 6361
rect 15198 6287 15200 6296
rect 15252 6287 15254 6296
rect 15200 6258 15252 6264
rect 15304 6202 15332 11494
rect 15672 10674 15700 11630
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15672 10130 15700 10610
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15396 9042 15424 9590
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15396 8498 15424 8978
rect 15476 8900 15528 8906
rect 15476 8842 15528 8848
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15488 7410 15516 8842
rect 15672 8838 15700 9522
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15672 8430 15700 8774
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15212 6174 15332 6202
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14936 5137 14964 5170
rect 14922 5128 14978 5137
rect 14922 5063 14978 5072
rect 15016 5092 15068 5098
rect 15016 5034 15068 5040
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14200 3738 14228 4694
rect 14292 4678 14504 4706
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14292 4282 14320 4558
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14292 3738 14320 4218
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14096 3528 14148 3534
rect 13924 3454 14044 3482
rect 14096 3470 14148 3476
rect 13910 3360 13966 3369
rect 13910 3295 13966 3304
rect 13924 3058 13952 3295
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13910 2816 13966 2825
rect 13910 2751 13966 2760
rect 13924 1426 13952 2751
rect 13912 1420 13964 1426
rect 13912 1362 13964 1368
rect 14016 800 14044 3454
rect 14108 2990 14136 3470
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14200 2854 14228 3674
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14292 3058 14320 3538
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14108 800 14136 2790
rect 14188 1216 14240 1222
rect 14188 1158 14240 1164
rect 14200 800 14228 1158
rect 14384 800 14412 3946
rect 14476 2922 14504 4678
rect 14832 4548 14884 4554
rect 14832 4490 14884 4496
rect 14648 4208 14700 4214
rect 14648 4150 14700 4156
rect 14556 3936 14608 3942
rect 14660 3913 14688 4150
rect 14738 4040 14794 4049
rect 14738 3975 14794 3984
rect 14752 3942 14780 3975
rect 14844 3942 14872 4490
rect 14924 4004 14976 4010
rect 14924 3946 14976 3952
rect 14740 3936 14792 3942
rect 14556 3878 14608 3884
rect 14646 3904 14702 3913
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14462 2816 14518 2825
rect 14462 2751 14518 2760
rect 14476 800 14504 2751
rect 14568 800 14596 3878
rect 14740 3878 14792 3884
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 14646 3839 14702 3848
rect 14660 2825 14688 3839
rect 14936 3738 14964 3946
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14646 2816 14702 2825
rect 14646 2751 14702 2760
rect 14646 2680 14702 2689
rect 14646 2615 14648 2624
rect 14700 2615 14702 2624
rect 14648 2586 14700 2592
rect 14752 2310 14780 2994
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14648 1420 14700 1426
rect 14648 1362 14700 1368
rect 14660 800 14688 1362
rect 14752 1154 14780 2246
rect 14832 2032 14884 2038
rect 14832 1974 14884 1980
rect 14922 2000 14978 2009
rect 14740 1148 14792 1154
rect 14740 1090 14792 1096
rect 14740 944 14792 950
rect 14740 886 14792 892
rect 14752 800 14780 886
rect 14844 800 14872 1974
rect 14922 1935 14978 1944
rect 14936 800 14964 1935
rect 15028 1222 15056 5034
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 15120 3194 15148 4490
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15212 3126 15240 6174
rect 15396 5710 15424 7278
rect 15488 6662 15516 7346
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 4146 15332 5578
rect 15764 5234 15792 12854
rect 16040 12442 16068 20810
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16132 19378 16160 20198
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16396 18692 16448 18698
rect 16396 18634 16448 18640
rect 16408 18290 16436 18634
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16408 17882 16436 18226
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16500 17513 16528 17546
rect 16486 17504 16542 17513
rect 16486 17439 16542 17448
rect 16592 17270 16620 21950
rect 16948 21898 17000 21904
rect 16764 21888 16816 21894
rect 16764 21830 16816 21836
rect 16776 21554 16804 21830
rect 16764 21548 16816 21554
rect 16764 21490 16816 21496
rect 16960 21350 16988 21898
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 16948 21344 17000 21350
rect 16948 21286 17000 21292
rect 16868 20942 16896 21286
rect 16960 21146 16988 21286
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 16856 20936 16908 20942
rect 16856 20878 16908 20884
rect 16948 20596 17000 20602
rect 16948 20538 17000 20544
rect 16764 20324 16816 20330
rect 16764 20266 16816 20272
rect 16776 19310 16804 20266
rect 16960 20262 16988 20538
rect 16948 20256 17000 20262
rect 16948 20198 17000 20204
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16960 17882 16988 18702
rect 16948 17876 17000 17882
rect 16948 17818 17000 17824
rect 16580 17264 16632 17270
rect 17052 17241 17080 22066
rect 17144 20602 17172 22630
rect 17236 22234 17264 22714
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17328 22114 17356 26982
rect 17592 24812 17644 24818
rect 17592 24754 17644 24760
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17512 23798 17540 24142
rect 17500 23792 17552 23798
rect 17500 23734 17552 23740
rect 17604 23730 17632 24754
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 17696 23610 17724 27814
rect 17868 26920 17920 26926
rect 17868 26862 17920 26868
rect 17880 24750 17908 26862
rect 17972 26518 18000 30806
rect 18052 30660 18104 30666
rect 18052 30602 18104 30608
rect 18064 30394 18092 30602
rect 18144 30592 18196 30598
rect 18144 30534 18196 30540
rect 18052 30388 18104 30394
rect 18052 30330 18104 30336
rect 18156 30326 18184 30534
rect 18144 30320 18196 30326
rect 18144 30262 18196 30268
rect 18248 29238 18276 31282
rect 18432 30938 18460 31282
rect 18708 30938 18736 32370
rect 19352 32026 19380 32846
rect 23676 32842 23704 33390
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 23664 32836 23716 32842
rect 23664 32778 23716 32784
rect 20168 32768 20220 32774
rect 20168 32710 20220 32716
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19340 32020 19392 32026
rect 19340 31962 19392 31968
rect 19156 31816 19208 31822
rect 19156 31758 19208 31764
rect 18972 31340 19024 31346
rect 18972 31282 19024 31288
rect 18420 30932 18472 30938
rect 18420 30874 18472 30880
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18984 30326 19012 31282
rect 18972 30320 19024 30326
rect 18972 30262 19024 30268
rect 18328 29640 18380 29646
rect 18328 29582 18380 29588
rect 18236 29232 18288 29238
rect 18236 29174 18288 29180
rect 18248 27470 18276 29174
rect 18340 28966 18368 29582
rect 19064 29164 19116 29170
rect 19064 29106 19116 29112
rect 18328 28960 18380 28966
rect 18328 28902 18380 28908
rect 18340 28558 18368 28902
rect 19076 28558 19104 29106
rect 18328 28552 18380 28558
rect 18328 28494 18380 28500
rect 19064 28552 19116 28558
rect 19064 28494 19116 28500
rect 18340 28422 18368 28494
rect 18328 28416 18380 28422
rect 18328 28358 18380 28364
rect 19076 27878 19104 28494
rect 19064 27872 19116 27878
rect 19064 27814 19116 27820
rect 18236 27464 18288 27470
rect 18236 27406 18288 27412
rect 17960 26512 18012 26518
rect 18012 26460 18092 26466
rect 17960 26454 18092 26460
rect 17972 26438 18092 26454
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17880 24274 17908 24686
rect 17972 24410 18000 26318
rect 18064 25974 18092 26438
rect 18248 25974 18276 27406
rect 18420 27328 18472 27334
rect 18420 27270 18472 27276
rect 18328 26988 18380 26994
rect 18328 26930 18380 26936
rect 18052 25968 18104 25974
rect 18052 25910 18104 25916
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 18340 25498 18368 26930
rect 18328 25492 18380 25498
rect 18328 25434 18380 25440
rect 17960 24404 18012 24410
rect 17960 24346 18012 24352
rect 18144 24336 18196 24342
rect 18144 24278 18196 24284
rect 17868 24268 17920 24274
rect 17868 24210 17920 24216
rect 17236 22086 17356 22114
rect 17512 23582 17724 23610
rect 17236 21622 17264 22086
rect 17224 21616 17276 21622
rect 17224 21558 17276 21564
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 17144 19990 17172 20538
rect 17132 19984 17184 19990
rect 17132 19926 17184 19932
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 17144 18290 17172 18566
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 16580 17206 16632 17212
rect 17038 17232 17094 17241
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 16132 13530 16160 14282
rect 16408 14006 16436 14037
rect 16396 14000 16448 14006
rect 16500 13954 16528 16730
rect 16592 15434 16620 17206
rect 16856 17196 16908 17202
rect 17038 17167 17094 17176
rect 16856 17138 16908 17144
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16522 16712 16934
rect 16672 16516 16724 16522
rect 16672 16458 16724 16464
rect 16868 15706 16896 17138
rect 17040 16720 17092 16726
rect 17040 16662 17092 16668
rect 17052 16454 17080 16662
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 16948 16108 17000 16114
rect 16948 16050 17000 16056
rect 16856 15700 16908 15706
rect 16856 15642 16908 15648
rect 16764 15632 16816 15638
rect 16764 15574 16816 15580
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16776 14414 16804 15574
rect 16960 15366 16988 16050
rect 17052 15502 17080 16390
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16960 14414 16988 15302
rect 17236 15026 17264 15506
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17236 14550 17264 14962
rect 17224 14544 17276 14550
rect 17224 14486 17276 14492
rect 16764 14408 16816 14414
rect 16764 14350 16816 14356
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16776 14074 16804 14350
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 17236 14006 17264 14486
rect 16448 13948 16528 13954
rect 16396 13942 16528 13948
rect 17224 14000 17276 14006
rect 17224 13942 17276 13948
rect 16408 13926 16528 13942
rect 16408 13530 16436 13926
rect 16488 13796 16540 13802
rect 16488 13738 16540 13744
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16212 13388 16264 13394
rect 16212 13330 16264 13336
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 16120 10192 16172 10198
rect 16120 10134 16172 10140
rect 16132 9722 16160 10134
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15948 9178 15976 9522
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16132 8566 16160 9046
rect 16120 8560 16172 8566
rect 16120 8502 16172 8508
rect 16224 7936 16252 13330
rect 16500 13326 16528 13738
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 16316 12238 16344 12582
rect 16408 12374 16436 12650
rect 17328 12434 17356 17478
rect 17420 16402 17448 17750
rect 17512 16538 17540 23582
rect 17684 23248 17736 23254
rect 17684 23190 17736 23196
rect 17696 22094 17724 23190
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 17788 22506 17816 23054
rect 17776 22500 17828 22506
rect 17776 22442 17828 22448
rect 17696 22066 17816 22094
rect 17788 21486 17816 22066
rect 17880 21622 17908 24210
rect 18156 24206 18184 24278
rect 18144 24200 18196 24206
rect 18144 24142 18196 24148
rect 18052 23656 18104 23662
rect 18052 23598 18104 23604
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 17972 22098 18000 22578
rect 18064 22574 18092 23598
rect 18142 23488 18198 23497
rect 18142 23423 18198 23432
rect 18052 22568 18104 22574
rect 18052 22510 18104 22516
rect 18064 22098 18092 22510
rect 17960 22092 18012 22098
rect 17960 22034 18012 22040
rect 18052 22092 18104 22098
rect 18052 22034 18104 22040
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17880 20942 17908 21558
rect 17972 21146 18000 22034
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 17868 20936 17920 20942
rect 17868 20878 17920 20884
rect 17972 20754 18000 21082
rect 18052 20868 18104 20874
rect 18052 20810 18104 20816
rect 17880 20726 18000 20754
rect 17880 17678 17908 20726
rect 18064 19990 18092 20810
rect 18156 20330 18184 23423
rect 18328 23112 18380 23118
rect 18328 23054 18380 23060
rect 18340 21894 18368 23054
rect 18432 22778 18460 27270
rect 18880 26376 18932 26382
rect 18880 26318 18932 26324
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18604 24744 18656 24750
rect 18604 24686 18656 24692
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18524 24206 18552 24550
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18524 23730 18552 24006
rect 18616 23798 18644 24686
rect 18708 24342 18736 25230
rect 18696 24336 18748 24342
rect 18696 24278 18748 24284
rect 18604 23792 18656 23798
rect 18604 23734 18656 23740
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 18420 22772 18472 22778
rect 18420 22714 18472 22720
rect 18604 22704 18656 22710
rect 18604 22646 18656 22652
rect 18512 22432 18564 22438
rect 18512 22374 18564 22380
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 18052 19984 18104 19990
rect 18052 19926 18104 19932
rect 17868 17672 17920 17678
rect 17868 17614 17920 17620
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17696 16726 17724 17070
rect 17880 17066 17908 17614
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17684 16720 17736 16726
rect 17684 16662 17736 16668
rect 17512 16510 17724 16538
rect 17880 16522 17908 17002
rect 18236 16992 18288 16998
rect 18236 16934 18288 16940
rect 18248 16794 18276 16934
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 17420 16374 17632 16402
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17236 12406 17356 12434
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16316 11694 16344 12174
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16592 10606 16620 12174
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16684 11558 16712 12038
rect 16776 11898 16804 12174
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16592 10198 16620 10542
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16684 9654 16712 11494
rect 16764 11280 16816 11286
rect 16764 11222 16816 11228
rect 16776 11014 16804 11222
rect 16868 11218 16896 11698
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 16764 11008 16816 11014
rect 16764 10950 16816 10956
rect 16776 10810 16804 10950
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16960 10130 16988 11018
rect 17144 10266 17172 11018
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16500 8906 16528 8978
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 16580 8492 16632 8498
rect 16580 8434 16632 8440
rect 16948 8492 17000 8498
rect 16948 8434 17000 8440
rect 16132 7908 16252 7936
rect 15936 7744 15988 7750
rect 15936 7686 15988 7692
rect 15948 5642 15976 7686
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15764 4842 15792 5170
rect 15936 5160 15988 5166
rect 15936 5102 15988 5108
rect 15844 5024 15896 5030
rect 15844 4966 15896 4972
rect 15672 4826 15792 4842
rect 15660 4820 15792 4826
rect 15712 4814 15792 4820
rect 15660 4762 15712 4768
rect 15752 4752 15804 4758
rect 15752 4694 15804 4700
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15304 3641 15332 3674
rect 15290 3632 15346 3641
rect 15290 3567 15346 3576
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15198 2952 15254 2961
rect 15198 2887 15200 2896
rect 15252 2887 15254 2896
rect 15200 2858 15252 2864
rect 15304 2854 15332 3567
rect 15396 3534 15424 4150
rect 15488 4146 15516 4422
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15488 3602 15516 4082
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15396 2990 15424 3470
rect 15488 2990 15516 3538
rect 15580 3194 15608 3878
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15476 2984 15528 2990
rect 15476 2926 15528 2932
rect 15580 2854 15608 3130
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15106 2680 15162 2689
rect 15106 2615 15162 2624
rect 15120 2582 15148 2615
rect 15108 2576 15160 2582
rect 15108 2518 15160 2524
rect 15198 2544 15254 2553
rect 15198 2479 15254 2488
rect 15292 2508 15344 2514
rect 15016 1216 15068 1222
rect 15016 1158 15068 1164
rect 15016 944 15068 950
rect 15016 886 15068 892
rect 15108 944 15160 950
rect 15108 886 15160 892
rect 15028 800 15056 886
rect 15120 800 15148 886
rect 15212 800 15240 2479
rect 15292 2450 15344 2456
rect 15304 800 15332 2450
rect 15382 2408 15438 2417
rect 15438 2352 15608 2360
rect 15382 2343 15384 2352
rect 15436 2332 15608 2352
rect 15384 2314 15436 2320
rect 15384 1964 15436 1970
rect 15384 1906 15436 1912
rect 15396 800 15424 1906
rect 15580 800 15608 2332
rect 15672 800 15700 4626
rect 15764 4146 15792 4694
rect 15856 4282 15884 4966
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15764 3738 15792 3878
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15856 800 15884 2246
rect 15948 800 15976 5102
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 16040 4690 16068 5034
rect 16028 4684 16080 4690
rect 16028 4626 16080 4632
rect 16132 3398 16160 7908
rect 16592 6866 16620 8434
rect 16960 8090 16988 8434
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16672 7336 16724 7342
rect 16672 7278 16724 7284
rect 16684 6934 16712 7278
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16672 6928 16724 6934
rect 16672 6870 16724 6876
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16776 6798 16804 7210
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16212 4616 16264 4622
rect 16212 4558 16264 4564
rect 16224 4214 16252 4558
rect 16212 4208 16264 4214
rect 16212 4150 16264 4156
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 16210 3088 16266 3097
rect 16210 3023 16266 3032
rect 16026 2680 16082 2689
rect 16026 2615 16028 2624
rect 16080 2615 16082 2624
rect 16028 2586 16080 2592
rect 16120 1760 16172 1766
rect 16120 1702 16172 1708
rect 16132 800 16160 1702
rect 16224 800 16252 3023
rect 16408 2378 16436 6734
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16500 3738 16528 4082
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16486 3632 16542 3641
rect 16486 3567 16488 3576
rect 16540 3567 16542 3576
rect 16488 3538 16540 3544
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16500 3194 16528 3402
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16592 2774 16620 6054
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16684 4146 16712 4626
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16776 3942 16804 6190
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16868 4282 16896 4558
rect 16948 4548 17000 4554
rect 16948 4490 17000 4496
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16764 3936 16816 3942
rect 16764 3878 16816 3884
rect 16868 3346 16896 4014
rect 16960 4010 16988 4490
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16500 2746 16620 2774
rect 16684 3318 16896 3346
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 16304 1896 16356 1902
rect 16304 1838 16356 1844
rect 16316 1034 16344 1838
rect 16408 1766 16436 2314
rect 16396 1760 16448 1766
rect 16396 1702 16448 1708
rect 16316 1006 16436 1034
rect 16408 800 16436 1006
rect 16500 800 16528 2746
rect 16684 898 16712 3318
rect 17236 2774 17264 12406
rect 17408 6452 17460 6458
rect 17408 6394 17460 6400
rect 17420 6254 17448 6394
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17512 3738 17540 14010
rect 17604 6866 17632 16374
rect 17696 9654 17724 16510
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 18156 16046 18184 16526
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18156 14958 18184 15982
rect 18144 14952 18196 14958
rect 18144 14894 18196 14900
rect 18248 13530 18276 16186
rect 18340 14550 18368 21830
rect 18524 21622 18552 22374
rect 18616 21894 18644 22646
rect 18708 22642 18736 24278
rect 18696 22636 18748 22642
rect 18696 22578 18748 22584
rect 18892 22506 18920 26318
rect 18880 22500 18932 22506
rect 18880 22442 18932 22448
rect 18604 21888 18656 21894
rect 18604 21830 18656 21836
rect 18512 21616 18564 21622
rect 18512 21558 18564 21564
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18524 19854 18552 20334
rect 18512 19848 18564 19854
rect 18512 19790 18564 19796
rect 18616 17542 18644 21830
rect 18892 21010 18920 22442
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18800 20602 18828 20742
rect 18788 20596 18840 20602
rect 18788 20538 18840 20544
rect 18892 20466 18920 20946
rect 18984 20806 19012 21286
rect 18972 20800 19024 20806
rect 18972 20742 19024 20748
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18788 19984 18840 19990
rect 18788 19926 18840 19932
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18708 18766 18736 19654
rect 18800 19378 18828 19926
rect 18880 19780 18932 19786
rect 18880 19722 18932 19728
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18892 19174 18920 19722
rect 18880 19168 18932 19174
rect 18880 19110 18932 19116
rect 18892 18970 18920 19110
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18984 18426 19012 20742
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18892 16794 18920 18226
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 17202 19012 18022
rect 18972 17196 19024 17202
rect 18972 17138 19024 17144
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18432 14618 18460 14962
rect 18420 14612 18472 14618
rect 18420 14554 18472 14560
rect 18328 14544 18380 14550
rect 18328 14486 18380 14492
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17880 12918 17908 13330
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17788 12306 17816 12718
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17880 11830 17908 12854
rect 18248 12850 18276 13466
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18524 11898 18552 14350
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 17868 11824 17920 11830
rect 17868 11766 17920 11772
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17880 8566 17908 11766
rect 17868 8560 17920 8566
rect 17868 8502 17920 8508
rect 17880 7954 17908 8502
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17604 6458 17632 6802
rect 17592 6452 17644 6458
rect 17592 6394 17644 6400
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17316 2916 17368 2922
rect 17316 2858 17368 2864
rect 16776 2746 17264 2774
rect 16776 2650 16804 2746
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 17038 1456 17094 1465
rect 17038 1391 17094 1400
rect 16684 870 16804 898
rect 16776 800 16804 870
rect 17052 800 17080 1391
rect 17328 800 17356 2858
rect 17500 2576 17552 2582
rect 17498 2544 17500 2553
rect 17552 2544 17554 2553
rect 17498 2479 17554 2488
rect 17604 800 17632 5646
rect 17880 5166 17908 7890
rect 17972 6322 18000 11834
rect 18616 11286 18644 12854
rect 18696 12844 18748 12850
rect 18696 12786 18748 12792
rect 18708 12102 18736 12786
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 18708 10198 18736 12038
rect 18696 10192 18748 10198
rect 18696 10134 18748 10140
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18064 8362 18092 10066
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18248 8838 18276 8910
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18052 8356 18104 8362
rect 18052 8298 18104 8304
rect 18064 7750 18092 8298
rect 18248 7818 18276 8774
rect 18236 7812 18288 7818
rect 18236 7754 18288 7760
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18248 7478 18276 7754
rect 18236 7472 18288 7478
rect 18236 7414 18288 7420
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18064 6458 18092 6734
rect 18052 6452 18104 6458
rect 18052 6394 18104 6400
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18524 6225 18552 6258
rect 18510 6216 18566 6225
rect 18510 6151 18566 6160
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 17868 5160 17920 5166
rect 17868 5102 17920 5108
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 17788 2774 17816 4966
rect 17880 4690 17908 5102
rect 17868 4684 17920 4690
rect 17868 4626 17920 4632
rect 17972 4146 18000 5238
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17788 2746 17908 2774
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17696 2106 17724 2382
rect 17684 2100 17736 2106
rect 17684 2042 17736 2048
rect 17696 1426 17724 2042
rect 17684 1420 17736 1426
rect 17684 1362 17736 1368
rect 17880 800 17908 2746
rect 18156 800 18184 5646
rect 18616 5030 18644 5714
rect 18696 5704 18748 5710
rect 18696 5646 18748 5652
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18248 3398 18276 4082
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 18432 800 18460 4966
rect 18616 4146 18644 4966
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18708 800 18736 5646
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18984 800 19012 4694
rect 19076 3126 19104 27814
rect 19168 26450 19196 31758
rect 19984 31680 20036 31686
rect 19984 31622 20036 31628
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19996 31346 20024 31622
rect 20180 31482 20208 32710
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 23388 32428 23440 32434
rect 23388 32370 23440 32376
rect 22744 32224 22796 32230
rect 22744 32166 22796 32172
rect 22284 32020 22336 32026
rect 22284 31962 22336 31968
rect 20628 31816 20680 31822
rect 20628 31758 20680 31764
rect 20168 31476 20220 31482
rect 20168 31418 20220 31424
rect 19984 31340 20036 31346
rect 19984 31282 20036 31288
rect 19432 30660 19484 30666
rect 19432 30602 19484 30608
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19248 29640 19300 29646
rect 19248 29582 19300 29588
rect 19260 28762 19288 29582
rect 19248 28756 19300 28762
rect 19248 28698 19300 28704
rect 19248 28416 19300 28422
rect 19248 28358 19300 28364
rect 19260 28082 19288 28358
rect 19352 28098 19380 30534
rect 19444 30122 19472 30602
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19432 30116 19484 30122
rect 19432 30058 19484 30064
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 20088 29578 20116 29990
rect 20076 29572 20128 29578
rect 20076 29514 20128 29520
rect 19432 29504 19484 29510
rect 19432 29446 19484 29452
rect 19444 29170 19472 29446
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 29164 19484 29170
rect 19432 29106 19484 29112
rect 19984 28960 20036 28966
rect 19984 28902 20036 28908
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19248 28076 19300 28082
rect 19352 28070 19564 28098
rect 19248 28018 19300 28024
rect 19260 27674 19288 28018
rect 19432 28008 19484 28014
rect 19432 27950 19484 27956
rect 19248 27668 19300 27674
rect 19248 27610 19300 27616
rect 19444 27606 19472 27950
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 19340 27396 19392 27402
rect 19340 27338 19392 27344
rect 19156 26444 19208 26450
rect 19156 26386 19208 26392
rect 19168 24750 19196 26386
rect 19352 25770 19380 27338
rect 19444 26042 19472 27542
rect 19536 27402 19564 28070
rect 19996 27946 20024 28902
rect 20088 28558 20116 29514
rect 20076 28552 20128 28558
rect 20076 28494 20128 28500
rect 20180 28218 20208 31418
rect 20260 30796 20312 30802
rect 20260 30738 20312 30744
rect 20272 28626 20300 30738
rect 20640 30734 20668 31758
rect 20996 31748 21048 31754
rect 20996 31690 21048 31696
rect 21008 31482 21036 31690
rect 22192 31680 22244 31686
rect 22192 31622 22244 31628
rect 20996 31476 21048 31482
rect 20996 31418 21048 31424
rect 22204 31414 22232 31622
rect 22296 31482 22324 31962
rect 22756 31754 22784 32166
rect 22744 31748 22796 31754
rect 22744 31690 22796 31696
rect 23216 31482 23244 32370
rect 23400 32026 23428 32370
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 23676 31958 23704 32778
rect 25332 32434 25360 32846
rect 25320 32428 25372 32434
rect 25320 32370 25372 32376
rect 25976 32026 26004 33458
rect 26332 33380 26384 33386
rect 26332 33322 26384 33328
rect 26056 33312 26108 33318
rect 26056 33254 26108 33260
rect 26068 33114 26096 33254
rect 26056 33108 26108 33114
rect 26056 33050 26108 33056
rect 26344 32978 26372 33322
rect 26332 32972 26384 32978
rect 26332 32914 26384 32920
rect 26804 32910 26832 33918
rect 27068 33866 27120 33872
rect 27080 33454 27108 33866
rect 27068 33448 27120 33454
rect 27068 33390 27120 33396
rect 27080 33114 27108 33390
rect 27068 33108 27120 33114
rect 27068 33050 27120 33056
rect 26792 32904 26844 32910
rect 26792 32846 26844 32852
rect 26424 32768 26476 32774
rect 26424 32710 26476 32716
rect 26436 32434 26464 32710
rect 26804 32570 26832 32846
rect 26792 32564 26844 32570
rect 26792 32506 26844 32512
rect 26424 32428 26476 32434
rect 26424 32370 26476 32376
rect 25964 32020 26016 32026
rect 25964 31962 26016 31968
rect 23664 31952 23716 31958
rect 23664 31894 23716 31900
rect 23676 31482 23704 31894
rect 24308 31748 24360 31754
rect 24308 31690 24360 31696
rect 24492 31748 24544 31754
rect 24492 31690 24544 31696
rect 24320 31634 24348 31690
rect 24320 31606 24440 31634
rect 22284 31476 22336 31482
rect 22284 31418 22336 31424
rect 23204 31476 23256 31482
rect 23204 31418 23256 31424
rect 23664 31476 23716 31482
rect 23664 31418 23716 31424
rect 22192 31408 22244 31414
rect 22192 31350 22244 31356
rect 22204 30938 22232 31350
rect 22744 31272 22796 31278
rect 22744 31214 22796 31220
rect 22192 30932 22244 30938
rect 22192 30874 22244 30880
rect 20628 30728 20680 30734
rect 20628 30670 20680 30676
rect 20536 30320 20588 30326
rect 20536 30262 20588 30268
rect 20640 30274 20668 30670
rect 21088 30660 21140 30666
rect 21088 30602 21140 30608
rect 21100 30394 21128 30602
rect 21916 30592 21968 30598
rect 21916 30534 21968 30540
rect 21088 30388 21140 30394
rect 21088 30330 21140 30336
rect 20260 28620 20312 28626
rect 20260 28562 20312 28568
rect 20168 28212 20220 28218
rect 20168 28154 20220 28160
rect 20180 28082 20208 28154
rect 20168 28076 20220 28082
rect 20088 28036 20168 28064
rect 19984 27940 20036 27946
rect 19984 27882 20036 27888
rect 19524 27396 19576 27402
rect 19524 27338 19576 27344
rect 19984 27328 20036 27334
rect 19984 27270 20036 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 27062 20024 27270
rect 19984 27056 20036 27062
rect 19984 26998 20036 27004
rect 19984 26784 20036 26790
rect 19984 26726 20036 26732
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 26036 19484 26042
rect 19432 25978 19484 25984
rect 19800 26036 19852 26042
rect 19800 25978 19852 25984
rect 19430 25936 19486 25945
rect 19812 25906 19840 25978
rect 19430 25871 19432 25880
rect 19484 25871 19486 25880
rect 19800 25900 19852 25906
rect 19432 25842 19484 25848
rect 19800 25842 19852 25848
rect 19340 25764 19392 25770
rect 19340 25706 19392 25712
rect 19444 25650 19472 25842
rect 19352 25622 19472 25650
rect 19156 24744 19208 24750
rect 19156 24686 19208 24692
rect 19352 24256 19380 25622
rect 19996 25362 20024 26726
rect 20088 26314 20116 28036
rect 20168 28018 20220 28024
rect 20168 27396 20220 27402
rect 20168 27338 20220 27344
rect 20076 26308 20128 26314
rect 20076 26250 20128 26256
rect 19984 25356 20036 25362
rect 19984 25298 20036 25304
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19444 24886 19472 25094
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19432 24880 19484 24886
rect 19432 24822 19484 24828
rect 20088 24818 20116 25230
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20180 24614 20208 27338
rect 20272 25786 20300 28562
rect 20352 27600 20404 27606
rect 20352 27542 20404 27548
rect 20364 27130 20392 27542
rect 20444 27532 20496 27538
rect 20444 27474 20496 27480
rect 20352 27124 20404 27130
rect 20352 27066 20404 27072
rect 20364 26450 20392 27066
rect 20352 26444 20404 26450
rect 20352 26386 20404 26392
rect 20364 25974 20392 26386
rect 20352 25968 20404 25974
rect 20456 25945 20484 27474
rect 20548 27033 20576 30262
rect 20640 30246 20760 30274
rect 20732 29170 20760 30246
rect 21928 30190 21956 30534
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 21916 30184 21968 30190
rect 21916 30126 21968 30132
rect 20720 29164 20772 29170
rect 20720 29106 20772 29112
rect 21732 29164 21784 29170
rect 21732 29106 21784 29112
rect 21744 28626 21772 29106
rect 21732 28620 21784 28626
rect 21732 28562 21784 28568
rect 21088 28484 21140 28490
rect 21272 28484 21324 28490
rect 21140 28444 21220 28472
rect 21088 28426 21140 28432
rect 20904 28416 20956 28422
rect 20904 28358 20956 28364
rect 20916 27470 20944 28358
rect 20904 27464 20956 27470
rect 20904 27406 20956 27412
rect 20812 27396 20864 27402
rect 20812 27338 20864 27344
rect 20534 27024 20590 27033
rect 20590 26994 20668 27010
rect 20590 26988 20680 26994
rect 20590 26982 20628 26988
rect 20534 26959 20590 26968
rect 20548 26899 20576 26959
rect 20628 26930 20680 26936
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 20352 25910 20404 25916
rect 20442 25936 20498 25945
rect 20442 25871 20498 25880
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 20272 25758 20392 25786
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 19260 24228 19380 24256
rect 19260 24154 19288 24228
rect 19168 24126 19288 24154
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 19340 24132 19392 24138
rect 19168 23594 19196 24126
rect 19340 24074 19392 24080
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19156 23588 19208 23594
rect 19156 23530 19208 23536
rect 19168 20398 19196 23530
rect 19260 23322 19288 23598
rect 19248 23316 19300 23322
rect 19248 23258 19300 23264
rect 19352 23118 19380 24074
rect 19444 23866 19472 24142
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23860 19484 23866
rect 19432 23802 19484 23808
rect 19984 23724 20036 23730
rect 19984 23666 20036 23672
rect 19524 23180 19576 23186
rect 19444 23140 19524 23168
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19444 21010 19472 23140
rect 19524 23122 19576 23128
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19524 22772 19576 22778
rect 19524 22714 19576 22720
rect 19536 22681 19564 22714
rect 19522 22672 19578 22681
rect 19522 22607 19578 22616
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21004 19484 21010
rect 19432 20946 19484 20952
rect 19444 20534 19472 20946
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19432 20528 19484 20534
rect 19432 20470 19484 20476
rect 19156 20392 19208 20398
rect 19156 20334 19208 20340
rect 19168 19854 19196 20334
rect 19892 20324 19944 20330
rect 19892 20266 19944 20272
rect 19248 20256 19300 20262
rect 19248 20198 19300 20204
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19260 18970 19288 20198
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19156 18760 19208 18766
rect 19156 18702 19208 18708
rect 19168 18290 19196 18702
rect 19260 18426 19288 18906
rect 19352 18834 19380 20198
rect 19800 19848 19852 19854
rect 19536 19796 19800 19802
rect 19536 19790 19852 19796
rect 19536 19786 19840 19790
rect 19904 19786 19932 20266
rect 19996 19922 20024 23666
rect 20180 23186 20208 24550
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 20168 23180 20220 23186
rect 20168 23122 20220 23128
rect 20272 22710 20300 23258
rect 20260 22704 20312 22710
rect 20260 22646 20312 22652
rect 20168 22636 20220 22642
rect 20168 22578 20220 22584
rect 20180 21350 20208 22578
rect 20272 21690 20300 22646
rect 20260 21684 20312 21690
rect 20260 21626 20312 21632
rect 20364 21554 20392 25758
rect 20444 25696 20496 25702
rect 20444 25638 20496 25644
rect 20456 24614 20484 25638
rect 20548 25226 20576 25842
rect 20536 25220 20588 25226
rect 20536 25162 20588 25168
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20456 24206 20484 24550
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20168 21344 20220 21350
rect 20168 21286 20220 21292
rect 20180 21146 20208 21286
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19524 19780 19840 19786
rect 19576 19774 19840 19780
rect 19892 19780 19944 19786
rect 19524 19722 19576 19728
rect 19892 19722 19944 19728
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 19446 19472 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 19446 20024 19858
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 20088 19378 20116 19654
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20180 19258 20208 21082
rect 20088 19230 20208 19258
rect 19432 19168 19484 19174
rect 19432 19110 19484 19116
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19340 18692 19392 18698
rect 19340 18634 19392 18640
rect 19352 18426 19380 18634
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19156 18284 19208 18290
rect 19156 18226 19208 18232
rect 19444 17338 19472 19110
rect 19984 18624 20036 18630
rect 19984 18566 20036 18572
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 17332 19484 17338
rect 19432 17274 19484 17280
rect 19996 17270 20024 18566
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19168 16726 19196 17138
rect 19156 16720 19208 16726
rect 19156 16662 19208 16668
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19352 15502 19380 16458
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19352 14906 19380 15302
rect 19444 15026 19472 17138
rect 19996 16590 20024 17206
rect 20088 17202 20116 19230
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19260 14878 19380 14906
rect 19260 14414 19288 14878
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19352 14278 19380 14758
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19168 13938 19196 14214
rect 19352 14074 19380 14214
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19168 12918 19196 13466
rect 19156 12912 19208 12918
rect 19156 12854 19208 12860
rect 19352 12850 19380 13670
rect 19444 13258 19472 14418
rect 19628 14414 19656 14758
rect 19616 14408 19668 14414
rect 19668 14356 19840 14362
rect 19616 14350 19840 14356
rect 19628 14346 19840 14350
rect 19628 14340 19852 14346
rect 19628 14334 19800 14340
rect 19800 14282 19852 14288
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 19904 13734 19932 13874
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19432 13252 19484 13258
rect 19432 13194 19484 13200
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19628 12646 19656 12786
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19260 11762 19288 12038
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19352 9178 19380 12582
rect 19996 12442 20024 15438
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19444 11354 19472 12174
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20088 11778 20116 16390
rect 20180 12986 20208 17138
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20168 12776 20220 12782
rect 20168 12718 20220 12724
rect 20180 12442 20208 12718
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20088 11750 20208 11778
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19812 11354 19840 11494
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19996 11150 20024 11494
rect 20076 11212 20128 11218
rect 20076 11154 20128 11160
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19984 11008 20036 11014
rect 19984 10950 20036 10956
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19996 10146 20024 10950
rect 19904 10118 20024 10146
rect 19904 9994 19932 10118
rect 20088 10010 20116 11154
rect 19892 9988 19944 9994
rect 19892 9930 19944 9936
rect 19996 9982 20116 10010
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19340 9172 19392 9178
rect 19340 9114 19392 9120
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8480 20024 9982
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 20088 9586 20116 9862
rect 20076 9580 20128 9586
rect 20076 9522 20128 9528
rect 20180 8974 20208 11750
rect 20272 10538 20300 17682
rect 20364 12968 20392 19110
rect 20456 17882 20484 24142
rect 20548 23730 20576 25162
rect 20732 24954 20760 26862
rect 20824 26518 20852 27338
rect 20812 26512 20864 26518
rect 20812 26454 20864 26460
rect 20720 24948 20772 24954
rect 20720 24890 20772 24896
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 21100 23866 21128 24074
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20536 23588 20588 23594
rect 20536 23530 20588 23536
rect 20548 23050 20576 23530
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 20536 23044 20588 23050
rect 20536 22986 20588 22992
rect 20548 22642 20576 22986
rect 20628 22976 20680 22982
rect 20628 22918 20680 22924
rect 20536 22636 20588 22642
rect 20536 22578 20588 22584
rect 20548 19258 20576 22578
rect 20640 22030 20668 22918
rect 20824 22642 20852 23054
rect 20904 23044 20956 23050
rect 20904 22986 20956 22992
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20732 20602 20760 22102
rect 20824 21690 20852 22578
rect 20916 22234 20944 22986
rect 21088 22432 21140 22438
rect 21088 22374 21140 22380
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 21100 22030 21128 22374
rect 21088 22024 21140 22030
rect 21088 21966 21140 21972
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 20824 20942 20852 21626
rect 21192 21622 21220 28444
rect 21272 28426 21324 28432
rect 21284 28218 21312 28426
rect 21928 28404 21956 30126
rect 22204 29646 22232 30194
rect 22756 30190 22784 31214
rect 24412 30802 24440 31606
rect 24504 31482 24532 31690
rect 25976 31482 26004 31962
rect 24492 31476 24544 31482
rect 24492 31418 24544 31424
rect 25964 31476 26016 31482
rect 25964 31418 26016 31424
rect 25504 31340 25556 31346
rect 25504 31282 25556 31288
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 24400 30796 24452 30802
rect 24400 30738 24452 30744
rect 22744 30184 22796 30190
rect 22744 30126 22796 30132
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 22008 28960 22060 28966
rect 22008 28902 22060 28908
rect 22020 28558 22048 28902
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 21928 28376 22048 28404
rect 21272 28212 21324 28218
rect 21272 28154 21324 28160
rect 22020 27538 22048 28376
rect 22112 28218 22140 29106
rect 22468 28416 22520 28422
rect 22468 28358 22520 28364
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 22480 28082 22508 28358
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 22756 28014 22784 30126
rect 24412 30054 24440 30738
rect 25516 30734 25544 31282
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 24676 30728 24728 30734
rect 24676 30670 24728 30676
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 24492 30592 24544 30598
rect 24492 30534 24544 30540
rect 24504 30326 24532 30534
rect 24492 30320 24544 30326
rect 24492 30262 24544 30268
rect 24400 30048 24452 30054
rect 24400 29990 24452 29996
rect 23848 29504 23900 29510
rect 23848 29446 23900 29452
rect 23112 28416 23164 28422
rect 23112 28358 23164 28364
rect 23124 28218 23152 28358
rect 23860 28218 23888 29446
rect 24412 28558 24440 29990
rect 24688 29850 24716 30670
rect 24768 30048 24820 30054
rect 24768 29990 24820 29996
rect 24676 29844 24728 29850
rect 24676 29786 24728 29792
rect 24780 29578 24808 29990
rect 24768 29572 24820 29578
rect 24768 29514 24820 29520
rect 24584 29164 24636 29170
rect 24584 29106 24636 29112
rect 24400 28552 24452 28558
rect 24400 28494 24452 28500
rect 23112 28212 23164 28218
rect 23112 28154 23164 28160
rect 23848 28212 23900 28218
rect 23848 28154 23900 28160
rect 22744 28008 22796 28014
rect 22744 27950 22796 27956
rect 22560 27668 22612 27674
rect 22560 27610 22612 27616
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 22020 25906 22048 27474
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 21456 24948 21508 24954
rect 21456 24890 21508 24896
rect 21468 22030 21496 24890
rect 21916 24812 21968 24818
rect 21916 24754 21968 24760
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21836 24138 21864 24550
rect 21824 24132 21876 24138
rect 21824 24074 21876 24080
rect 21928 22982 21956 24754
rect 22572 24750 22600 27610
rect 22652 27464 22704 27470
rect 22652 27406 22704 27412
rect 22664 26586 22692 27406
rect 23124 26926 23152 28154
rect 23860 28082 23888 28154
rect 23848 28076 23900 28082
rect 23848 28018 23900 28024
rect 24216 28008 24268 28014
rect 24216 27950 24268 27956
rect 23204 27532 23256 27538
rect 23204 27474 23256 27480
rect 23216 27130 23244 27474
rect 23296 27328 23348 27334
rect 23296 27270 23348 27276
rect 23664 27328 23716 27334
rect 23664 27270 23716 27276
rect 23204 27124 23256 27130
rect 23204 27066 23256 27072
rect 23112 26920 23164 26926
rect 23112 26862 23164 26868
rect 22744 26852 22796 26858
rect 22744 26794 22796 26800
rect 22652 26580 22704 26586
rect 22652 26522 22704 26528
rect 22756 25974 22784 26794
rect 22744 25968 22796 25974
rect 22744 25910 22796 25916
rect 22756 25838 22784 25910
rect 23124 25906 23152 26862
rect 23216 26450 23244 27066
rect 23204 26444 23256 26450
rect 23204 26386 23256 26392
rect 23308 26382 23336 27270
rect 23676 26994 23704 27270
rect 24228 27130 24256 27950
rect 24412 27606 24440 28494
rect 24596 28218 24624 29106
rect 24676 28960 24728 28966
rect 24676 28902 24728 28908
rect 24688 28558 24716 28902
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24584 28212 24636 28218
rect 24584 28154 24636 28160
rect 24400 27600 24452 27606
rect 24400 27542 24452 27548
rect 24780 27470 24808 29514
rect 25412 29504 25464 29510
rect 25412 29446 25464 29452
rect 25424 28694 25452 29446
rect 25412 28688 25464 28694
rect 25412 28630 25464 28636
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 24860 28212 24912 28218
rect 24860 28154 24912 28160
rect 24768 27464 24820 27470
rect 24768 27406 24820 27412
rect 24216 27124 24268 27130
rect 24216 27066 24268 27072
rect 23664 26988 23716 26994
rect 23664 26930 23716 26936
rect 23572 26512 23624 26518
rect 23572 26454 23624 26460
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 22744 25832 22796 25838
rect 22744 25774 22796 25780
rect 22756 25498 22784 25774
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 22560 24744 22612 24750
rect 22560 24686 22612 24692
rect 22572 24274 22600 24686
rect 22100 24268 22152 24274
rect 22100 24210 22152 24216
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22112 23186 22140 24210
rect 22848 23866 22876 25298
rect 23124 25294 23152 25842
rect 23020 25288 23072 25294
rect 23020 25230 23072 25236
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23032 23866 23060 25230
rect 23296 24608 23348 24614
rect 23296 24550 23348 24556
rect 22836 23860 22888 23866
rect 22836 23802 22888 23808
rect 23020 23860 23072 23866
rect 23020 23802 23072 23808
rect 23308 23644 23336 24550
rect 23584 24342 23612 26454
rect 23572 24336 23624 24342
rect 23572 24278 23624 24284
rect 23388 24132 23440 24138
rect 23388 24074 23440 24080
rect 23400 23798 23428 24074
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23388 23656 23440 23662
rect 23308 23616 23388 23644
rect 23388 23598 23440 23604
rect 23400 23254 23428 23598
rect 23676 23526 23704 26930
rect 24872 26450 24900 28154
rect 25056 28082 25084 28358
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 24952 26920 25004 26926
rect 24952 26862 25004 26868
rect 24860 26444 24912 26450
rect 24860 26386 24912 26392
rect 24492 26240 24544 26246
rect 24492 26182 24544 26188
rect 24504 25906 24532 26182
rect 24216 25900 24268 25906
rect 24216 25842 24268 25848
rect 24492 25900 24544 25906
rect 24492 25842 24544 25848
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24228 25498 24256 25842
rect 24216 25492 24268 25498
rect 24216 25434 24268 25440
rect 24504 24818 24532 25842
rect 24688 25294 24716 25842
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24872 25362 24900 25638
rect 24860 25356 24912 25362
rect 24860 25298 24912 25304
rect 24964 25294 24992 26862
rect 24676 25288 24728 25294
rect 24676 25230 24728 25236
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 24492 24812 24544 24818
rect 24492 24754 24544 24760
rect 24768 24608 24820 24614
rect 24768 24550 24820 24556
rect 24780 24342 24808 24550
rect 24768 24336 24820 24342
rect 24768 24278 24820 24284
rect 25056 24274 25084 28018
rect 25412 27328 25464 27334
rect 25412 27270 25464 27276
rect 25136 26988 25188 26994
rect 25136 26930 25188 26936
rect 25148 26450 25176 26930
rect 25136 26444 25188 26450
rect 25136 26386 25188 26392
rect 25148 25226 25176 26386
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 25136 25220 25188 25226
rect 25136 25162 25188 25168
rect 25044 24268 25096 24274
rect 25044 24210 25096 24216
rect 24584 24132 24636 24138
rect 24584 24074 24636 24080
rect 24596 23866 24624 24074
rect 23756 23860 23808 23866
rect 23756 23802 23808 23808
rect 24584 23860 24636 23866
rect 24584 23802 24636 23808
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 23388 23248 23440 23254
rect 23388 23190 23440 23196
rect 22100 23180 22152 23186
rect 22100 23122 22152 23128
rect 21916 22976 21968 22982
rect 21916 22918 21968 22924
rect 21548 22636 21600 22642
rect 21548 22578 21600 22584
rect 21560 22234 21588 22578
rect 22112 22574 22140 23122
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22100 22568 22152 22574
rect 22100 22510 22152 22516
rect 22284 22568 22336 22574
rect 22284 22510 22336 22516
rect 21548 22228 21600 22234
rect 21548 22170 21600 22176
rect 22296 22098 22324 22510
rect 22284 22092 22336 22098
rect 22284 22034 22336 22040
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21284 21690 21312 21966
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21824 21684 21876 21690
rect 21824 21626 21876 21632
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 21180 21616 21232 21622
rect 21180 21558 21232 21564
rect 21364 21616 21416 21622
rect 21364 21558 21416 21564
rect 20996 21548 21048 21554
rect 20996 21490 21048 21496
rect 20904 21344 20956 21350
rect 20904 21286 20956 21292
rect 20916 21010 20944 21286
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 20812 20936 20864 20942
rect 20812 20878 20864 20884
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20824 19990 20852 20878
rect 20916 20330 20944 20946
rect 21008 20534 21036 21490
rect 20996 20528 21048 20534
rect 20996 20470 21048 20476
rect 20904 20324 20956 20330
rect 20904 20266 20956 20272
rect 20916 19990 20944 20266
rect 20812 19984 20864 19990
rect 20812 19926 20864 19932
rect 20904 19984 20956 19990
rect 20904 19926 20956 19932
rect 20628 19712 20680 19718
rect 20628 19654 20680 19660
rect 20640 19514 20668 19654
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20996 19440 21048 19446
rect 20996 19382 21048 19388
rect 20548 19230 20668 19258
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20548 18766 20576 19110
rect 20536 18760 20588 18766
rect 20536 18702 20588 18708
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20456 16250 20484 17818
rect 20640 17678 20668 19230
rect 20812 19236 20864 19242
rect 20812 19178 20864 19184
rect 20904 19236 20956 19242
rect 20904 19178 20956 19184
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20640 17202 20668 17614
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20640 15366 20668 15397
rect 20628 15360 20680 15366
rect 20732 15314 20760 18362
rect 20824 18222 20852 19178
rect 20812 18216 20864 18222
rect 20812 18158 20864 18164
rect 20916 18154 20944 19178
rect 20904 18148 20956 18154
rect 20904 18090 20956 18096
rect 21008 18086 21036 19382
rect 21100 19310 21128 21558
rect 21180 21480 21232 21486
rect 21180 21422 21232 21428
rect 21192 21146 21220 21422
rect 21180 21140 21232 21146
rect 21180 21082 21232 21088
rect 21376 20874 21404 21558
rect 21836 21350 21864 21626
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 21364 20868 21416 20874
rect 21364 20810 21416 20816
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22112 20210 22140 20470
rect 22204 20398 22232 21898
rect 22296 20942 22324 22034
rect 22848 22030 22876 23054
rect 23400 22778 23428 23190
rect 23480 23044 23532 23050
rect 23480 22986 23532 22992
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 23492 22506 23520 22986
rect 23480 22500 23532 22506
rect 23480 22442 23532 22448
rect 23492 22030 23520 22442
rect 22836 22024 22888 22030
rect 22836 21966 22888 21972
rect 23480 22024 23532 22030
rect 23480 21966 23532 21972
rect 23676 21690 23704 23462
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 22928 21548 22980 21554
rect 22928 21490 22980 21496
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22468 20868 22520 20874
rect 22468 20810 22520 20816
rect 22192 20392 22244 20398
rect 22192 20334 22244 20340
rect 22284 20256 22336 20262
rect 22112 20182 22232 20210
rect 22284 20198 22336 20204
rect 22204 20058 22232 20182
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 20996 18080 21048 18086
rect 20996 18022 21048 18028
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20824 17338 20852 17614
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 21008 17184 21036 18022
rect 21100 17814 21128 19246
rect 21088 17808 21140 17814
rect 21088 17750 21140 17756
rect 21192 17542 21220 19314
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21284 17678 21312 18702
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21088 17196 21140 17202
rect 21008 17156 21088 17184
rect 21088 17138 21140 17144
rect 20680 15308 20760 15314
rect 20628 15302 20760 15308
rect 20640 15286 20760 15302
rect 20640 15162 20668 15286
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20548 14618 20576 14962
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20548 13870 20576 14418
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20364 12940 20484 12968
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20364 10810 20392 12786
rect 20456 12646 20484 12940
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20456 11898 20484 12106
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20548 11218 20576 13806
rect 20732 12850 20760 14010
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20640 10690 20668 12038
rect 20732 11558 20760 12786
rect 20824 11762 20852 13806
rect 20916 13530 20944 14350
rect 20996 14272 21048 14278
rect 20996 14214 21048 14220
rect 21008 13938 21036 14214
rect 20996 13932 21048 13938
rect 20996 13874 21048 13880
rect 21100 13734 21128 17138
rect 21284 15026 21312 17614
rect 22204 16658 22232 19994
rect 22296 19854 22324 20198
rect 22480 20058 22508 20810
rect 22940 20806 22968 21490
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 22928 20800 22980 20806
rect 22928 20742 22980 20748
rect 22836 20392 22888 20398
rect 22836 20334 22888 20340
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22560 17604 22612 17610
rect 22560 17546 22612 17552
rect 22572 17338 22600 17546
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 22284 17196 22336 17202
rect 22284 17138 22336 17144
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21652 15094 21680 16526
rect 22204 15706 22232 16594
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22296 15502 22324 17138
rect 22756 17105 22784 18362
rect 22742 17096 22798 17105
rect 22742 17031 22798 17040
rect 22848 16454 22876 20334
rect 22940 19446 22968 20742
rect 23584 20602 23612 21082
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 23388 20256 23440 20262
rect 23388 20198 23440 20204
rect 23020 19848 23072 19854
rect 23020 19790 23072 19796
rect 22928 19440 22980 19446
rect 22928 19382 22980 19388
rect 23032 19310 23060 19790
rect 23400 19378 23428 20198
rect 23768 20058 23796 23802
rect 24676 22976 24728 22982
rect 24676 22918 24728 22924
rect 24308 22228 24360 22234
rect 24308 22170 24360 22176
rect 24320 21894 24348 22170
rect 24400 22092 24452 22098
rect 24400 22034 24452 22040
rect 24308 21888 24360 21894
rect 24308 21830 24360 21836
rect 23756 20052 23808 20058
rect 23756 19994 23808 20000
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23020 19304 23072 19310
rect 23020 19246 23072 19252
rect 23032 18698 23060 19246
rect 23020 18692 23072 18698
rect 23020 18634 23072 18640
rect 23032 17814 23060 18634
rect 23400 18290 23428 19314
rect 23676 18426 23704 19450
rect 24320 19242 24348 21830
rect 24412 19378 24440 22034
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 24504 21350 24532 21966
rect 24688 21962 24716 22918
rect 24676 21956 24728 21962
rect 24676 21898 24728 21904
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24768 21344 24820 21350
rect 24768 21286 24820 21292
rect 24504 21146 24532 21286
rect 24492 21140 24544 21146
rect 24492 21082 24544 21088
rect 24780 20874 24808 21286
rect 25056 21078 25084 24210
rect 25134 22536 25190 22545
rect 25134 22471 25136 22480
rect 25188 22471 25190 22480
rect 25136 22442 25188 22448
rect 25044 21072 25096 21078
rect 24964 21032 25044 21060
rect 24768 20868 24820 20874
rect 24768 20810 24820 20816
rect 24780 20466 24808 20810
rect 24768 20460 24820 20466
rect 24768 20402 24820 20408
rect 24964 20262 24992 21032
rect 25044 21014 25096 21020
rect 24952 20256 25004 20262
rect 24952 20198 25004 20204
rect 25240 19446 25268 26318
rect 25424 25838 25452 27270
rect 25792 27130 25820 31214
rect 27172 30870 27200 31282
rect 27160 30864 27212 30870
rect 27160 30806 27212 30812
rect 25964 30660 26016 30666
rect 25964 30602 26016 30608
rect 25976 30394 26004 30602
rect 25964 30388 26016 30394
rect 25964 30330 26016 30336
rect 26240 27872 26292 27878
rect 26240 27814 26292 27820
rect 26252 27402 26280 27814
rect 26240 27396 26292 27402
rect 26240 27338 26292 27344
rect 25780 27124 25832 27130
rect 25780 27066 25832 27072
rect 25872 26852 25924 26858
rect 25872 26794 25924 26800
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 25412 25832 25464 25838
rect 25412 25774 25464 25780
rect 25516 25498 25544 25842
rect 25596 25764 25648 25770
rect 25596 25706 25648 25712
rect 25504 25492 25556 25498
rect 25504 25434 25556 25440
rect 25608 25294 25636 25706
rect 25596 25288 25648 25294
rect 25596 25230 25648 25236
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25516 21486 25544 21898
rect 25504 21480 25556 21486
rect 25504 21422 25556 21428
rect 25608 21146 25636 25230
rect 25688 25152 25740 25158
rect 25688 25094 25740 25100
rect 25700 24750 25728 25094
rect 25688 24744 25740 24750
rect 25688 24686 25740 24692
rect 25700 23866 25728 24686
rect 25780 24268 25832 24274
rect 25780 24210 25832 24216
rect 25688 23860 25740 23866
rect 25688 23802 25740 23808
rect 25792 23730 25820 24210
rect 25780 23724 25832 23730
rect 25780 23666 25832 23672
rect 25884 22778 25912 26794
rect 27264 25498 27292 34002
rect 27632 33862 27660 34342
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 29092 34128 29144 34134
rect 29092 34070 29144 34076
rect 27896 34060 27948 34066
rect 27896 34002 27948 34008
rect 29000 34060 29052 34066
rect 29000 34002 29052 34008
rect 27436 33856 27488 33862
rect 27436 33798 27488 33804
rect 27620 33856 27672 33862
rect 27620 33798 27672 33804
rect 27448 32910 27476 33798
rect 27436 32904 27488 32910
rect 27436 32846 27488 32852
rect 27632 32298 27660 33798
rect 27710 33552 27766 33561
rect 27908 33522 27936 34002
rect 28172 33856 28224 33862
rect 28172 33798 28224 33804
rect 28816 33856 28868 33862
rect 28816 33798 28868 33804
rect 28184 33590 28212 33798
rect 28172 33584 28224 33590
rect 28172 33526 28224 33532
rect 27710 33487 27712 33496
rect 27764 33487 27766 33496
rect 27897 33516 27949 33522
rect 27712 33458 27764 33464
rect 27897 33458 27949 33464
rect 28080 33516 28132 33522
rect 28080 33458 28132 33464
rect 28448 33516 28500 33522
rect 28448 33458 28500 33464
rect 28092 33386 28120 33458
rect 28080 33380 28132 33386
rect 28080 33322 28132 33328
rect 28264 33380 28316 33386
rect 28460 33368 28488 33458
rect 28828 33454 28856 33798
rect 28908 33584 28960 33590
rect 28906 33552 28908 33561
rect 28960 33552 28962 33561
rect 28906 33487 28962 33496
rect 28816 33448 28868 33454
rect 28816 33390 28868 33396
rect 28316 33340 28488 33368
rect 28264 33322 28316 33328
rect 28356 32904 28408 32910
rect 28356 32846 28408 32852
rect 28632 32904 28684 32910
rect 28632 32846 28684 32852
rect 27896 32428 27948 32434
rect 27896 32370 27948 32376
rect 27620 32292 27672 32298
rect 27620 32234 27672 32240
rect 27632 32026 27660 32234
rect 27620 32020 27672 32026
rect 27620 31962 27672 31968
rect 27908 31890 27936 32370
rect 27896 31884 27948 31890
rect 27896 31826 27948 31832
rect 27436 31748 27488 31754
rect 27436 31690 27488 31696
rect 27448 31210 27476 31690
rect 28368 31482 28396 32846
rect 28644 32570 28672 32846
rect 28632 32564 28684 32570
rect 28632 32506 28684 32512
rect 28828 32450 28856 33390
rect 29012 32910 29040 34002
rect 29104 33522 29132 34070
rect 31208 33652 31260 33658
rect 31208 33594 31260 33600
rect 32404 33652 32456 33658
rect 32404 33594 32456 33600
rect 29092 33516 29144 33522
rect 29092 33458 29144 33464
rect 31220 33386 31248 33594
rect 31116 33380 31168 33386
rect 31116 33322 31168 33328
rect 31208 33380 31260 33386
rect 31208 33322 31260 33328
rect 29000 32904 29052 32910
rect 29000 32846 29052 32852
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 28736 32422 28856 32450
rect 29012 32434 29040 32846
rect 29000 32428 29052 32434
rect 28736 32366 28764 32422
rect 29000 32370 29052 32376
rect 29748 32366 29776 32846
rect 28724 32360 28776 32366
rect 28724 32302 28776 32308
rect 29736 32360 29788 32366
rect 29736 32302 29788 32308
rect 28448 31680 28500 31686
rect 28448 31622 28500 31628
rect 28816 31680 28868 31686
rect 28816 31622 28868 31628
rect 28460 31482 28488 31622
rect 28356 31476 28408 31482
rect 28356 31418 28408 31424
rect 28448 31476 28500 31482
rect 28448 31418 28500 31424
rect 28828 31414 28856 31622
rect 29748 31482 29776 32302
rect 29736 31476 29788 31482
rect 29736 31418 29788 31424
rect 28816 31408 28868 31414
rect 28816 31350 28868 31356
rect 28356 31272 28408 31278
rect 28356 31214 28408 31220
rect 27436 31204 27488 31210
rect 27436 31146 27488 31152
rect 27448 30734 27476 31146
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27448 30138 27476 30670
rect 27528 30592 27580 30598
rect 27528 30534 27580 30540
rect 27896 30592 27948 30598
rect 27896 30534 27948 30540
rect 27540 30258 27568 30534
rect 27908 30326 27936 30534
rect 27896 30320 27948 30326
rect 27896 30262 27948 30268
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 27908 30190 27936 30262
rect 28368 30258 28396 31214
rect 29644 30660 29696 30666
rect 29644 30602 29696 30608
rect 29000 30592 29052 30598
rect 29000 30534 29052 30540
rect 28356 30252 28408 30258
rect 28356 30194 28408 30200
rect 28816 30252 28868 30258
rect 28816 30194 28868 30200
rect 27896 30184 27948 30190
rect 27448 30110 27568 30138
rect 27896 30126 27948 30132
rect 27540 29714 27568 30110
rect 28368 29714 28396 30194
rect 28828 29850 28856 30194
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 27528 29708 27580 29714
rect 27528 29650 27580 29656
rect 28356 29708 28408 29714
rect 28356 29650 28408 29656
rect 27540 28014 27568 29650
rect 29012 29646 29040 30534
rect 29656 30054 29684 30602
rect 30840 30252 30892 30258
rect 30840 30194 30892 30200
rect 29644 30048 29696 30054
rect 29644 29990 29696 29996
rect 30656 30048 30708 30054
rect 30656 29990 30708 29996
rect 29000 29640 29052 29646
rect 29000 29582 29052 29588
rect 29656 28558 29684 29990
rect 30472 29708 30524 29714
rect 30472 29650 30524 29656
rect 30484 29238 30512 29650
rect 30668 29578 30696 29990
rect 30656 29572 30708 29578
rect 30656 29514 30708 29520
rect 30472 29232 30524 29238
rect 30472 29174 30524 29180
rect 30196 28960 30248 28966
rect 30196 28902 30248 28908
rect 29644 28552 29696 28558
rect 29644 28494 29696 28500
rect 28816 28484 28868 28490
rect 28816 28426 28868 28432
rect 28264 28416 28316 28422
rect 28264 28358 28316 28364
rect 28276 28014 28304 28358
rect 28356 28076 28408 28082
rect 28356 28018 28408 28024
rect 27344 28008 27396 28014
rect 27344 27950 27396 27956
rect 27528 28008 27580 28014
rect 27528 27950 27580 27956
rect 28264 28008 28316 28014
rect 28264 27950 28316 27956
rect 27356 27334 27384 27950
rect 27344 27328 27396 27334
rect 27344 27270 27396 27276
rect 27252 25492 27304 25498
rect 27252 25434 27304 25440
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26608 23860 26660 23866
rect 26608 23802 26660 23808
rect 26056 23656 26108 23662
rect 26056 23598 26108 23604
rect 25872 22772 25924 22778
rect 25872 22714 25924 22720
rect 26068 21554 26096 23598
rect 26620 23118 26648 23802
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 26608 23112 26660 23118
rect 26608 23054 26660 23060
rect 26240 23044 26292 23050
rect 26240 22986 26292 22992
rect 26252 21690 26280 22986
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 26344 22030 26372 22374
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 26436 21894 26464 23054
rect 26424 21888 26476 21894
rect 26424 21830 26476 21836
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 26712 21554 26740 25230
rect 27356 24206 27384 27270
rect 27540 27130 27568 27950
rect 28368 27674 28396 28018
rect 28356 27668 28408 27674
rect 28356 27610 28408 27616
rect 28828 27470 28856 28426
rect 30208 28082 30236 28902
rect 30852 28762 30880 30194
rect 30840 28756 30892 28762
rect 30840 28698 30892 28704
rect 30932 28620 30984 28626
rect 30932 28562 30984 28568
rect 30196 28076 30248 28082
rect 30196 28018 30248 28024
rect 30944 28014 30972 28562
rect 29644 28008 29696 28014
rect 29644 27950 29696 27956
rect 30932 28008 30984 28014
rect 30932 27950 30984 27956
rect 31024 28008 31076 28014
rect 31024 27950 31076 27956
rect 29368 27532 29420 27538
rect 29368 27474 29420 27480
rect 28816 27464 28868 27470
rect 28816 27406 28868 27412
rect 29000 27328 29052 27334
rect 29000 27270 29052 27276
rect 27528 27124 27580 27130
rect 27528 27066 27580 27072
rect 27436 26988 27488 26994
rect 27436 26930 27488 26936
rect 27448 26586 27476 26930
rect 27436 26580 27488 26586
rect 27436 26522 27488 26528
rect 27344 24200 27396 24206
rect 27344 24142 27396 24148
rect 27252 24132 27304 24138
rect 27252 24074 27304 24080
rect 27068 24064 27120 24070
rect 27068 24006 27120 24012
rect 27080 23662 27108 24006
rect 27264 23798 27292 24074
rect 27252 23792 27304 23798
rect 27252 23734 27304 23740
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 27068 23656 27120 23662
rect 27068 23598 27120 23604
rect 26792 22772 26844 22778
rect 26792 22714 26844 22720
rect 26804 22574 26832 22714
rect 26792 22568 26844 22574
rect 26792 22510 26844 22516
rect 26056 21548 26108 21554
rect 26056 21490 26108 21496
rect 26700 21548 26752 21554
rect 26700 21490 26752 21496
rect 25780 21480 25832 21486
rect 25780 21422 25832 21428
rect 25596 21140 25648 21146
rect 25596 21082 25648 21088
rect 25792 20942 25820 21422
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 25792 20602 25820 20878
rect 25780 20596 25832 20602
rect 25780 20538 25832 20544
rect 25976 20398 26004 20878
rect 25964 20392 26016 20398
rect 25964 20334 26016 20340
rect 25780 20256 25832 20262
rect 25780 20198 25832 20204
rect 25792 19922 25820 20198
rect 26068 19990 26096 21490
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 26436 20534 26464 20742
rect 26424 20528 26476 20534
rect 26424 20470 26476 20476
rect 26056 19984 26108 19990
rect 26056 19926 26108 19932
rect 25780 19916 25832 19922
rect 25780 19858 25832 19864
rect 25228 19440 25280 19446
rect 25228 19382 25280 19388
rect 24400 19372 24452 19378
rect 24400 19314 24452 19320
rect 24676 19372 24728 19378
rect 24676 19314 24728 19320
rect 24308 19236 24360 19242
rect 24308 19178 24360 19184
rect 24688 18970 24716 19314
rect 25792 19174 25820 19858
rect 26240 19848 26292 19854
rect 26240 19790 26292 19796
rect 26252 19174 26280 19790
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 24676 18964 24728 18970
rect 24676 18906 24728 18912
rect 25792 18834 25820 19110
rect 25780 18828 25832 18834
rect 25780 18770 25832 18776
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23112 18148 23164 18154
rect 23112 18090 23164 18096
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 23124 17202 23152 18090
rect 23492 17898 23520 18090
rect 23308 17870 23520 17898
rect 23112 17196 23164 17202
rect 23112 17138 23164 17144
rect 22928 16992 22980 16998
rect 22928 16934 22980 16940
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22848 16182 22876 16390
rect 22836 16176 22888 16182
rect 22836 16118 22888 16124
rect 22652 16040 22704 16046
rect 22652 15982 22704 15988
rect 22284 15496 22336 15502
rect 22284 15438 22336 15444
rect 22468 15496 22520 15502
rect 22468 15438 22520 15444
rect 22296 15162 22324 15438
rect 22376 15360 22428 15366
rect 22376 15302 22428 15308
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 22388 15094 22416 15302
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 22008 15088 22060 15094
rect 22376 15088 22428 15094
rect 22060 15036 22140 15042
rect 22008 15030 22140 15036
rect 22376 15030 22428 15036
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21652 14346 21680 15030
rect 22020 15014 22140 15030
rect 21732 14816 21784 14822
rect 21732 14758 21784 14764
rect 21640 14340 21692 14346
rect 21640 14282 21692 14288
rect 21652 14006 21680 14282
rect 21744 14278 21772 14758
rect 22112 14414 22140 15014
rect 22480 14618 22508 15438
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21640 14000 21692 14006
rect 21640 13942 21692 13948
rect 21088 13728 21140 13734
rect 21088 13670 21140 13676
rect 20904 13524 20956 13530
rect 20956 13484 21036 13512
rect 20904 13466 20956 13472
rect 20904 13252 20956 13258
rect 20904 13194 20956 13200
rect 20916 12442 20944 13194
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 20364 10662 20668 10690
rect 20824 10674 20852 11698
rect 20812 10668 20864 10674
rect 20260 10532 20312 10538
rect 20260 10474 20312 10480
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20168 8492 20220 8498
rect 19996 8452 20168 8480
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19156 7948 19208 7954
rect 19156 7890 19208 7896
rect 19168 7410 19196 7890
rect 19260 7886 19288 8298
rect 19248 7880 19300 7886
rect 19248 7822 19300 7828
rect 19432 7812 19484 7818
rect 19432 7754 19484 7760
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19340 7404 19392 7410
rect 19444 7392 19472 7754
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19800 7404 19852 7410
rect 19444 7364 19800 7392
rect 19340 7346 19392 7352
rect 19800 7346 19852 7352
rect 19352 6730 19380 7346
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19444 6458 19472 6598
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6452 19484 6458
rect 19432 6394 19484 6400
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 19156 6316 19208 6322
rect 19156 6258 19208 6264
rect 19168 4010 19196 6258
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19352 4622 19380 6054
rect 19812 5778 19840 6326
rect 19996 5778 20024 8452
rect 20168 8434 20220 8440
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20180 7818 20208 8026
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 20364 7546 20392 10662
rect 20812 10610 20864 10616
rect 20536 10600 20588 10606
rect 20536 10542 20588 10548
rect 20548 10266 20576 10542
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20640 9722 20668 10406
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20916 9586 20944 12174
rect 21008 12102 21036 13484
rect 21272 12640 21324 12646
rect 21272 12582 21324 12588
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 21008 10538 21036 11698
rect 21100 11286 21128 12378
rect 21284 12238 21312 12582
rect 21744 12374 21772 14214
rect 22008 13932 22060 13938
rect 22008 13874 22060 13880
rect 21824 13728 21876 13734
rect 21824 13670 21876 13676
rect 21836 13326 21864 13670
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 22020 12986 22048 13874
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 21916 12844 21968 12850
rect 21916 12786 21968 12792
rect 21928 12442 21956 12786
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 21732 12368 21784 12374
rect 21732 12310 21784 12316
rect 21272 12232 21324 12238
rect 21272 12174 21324 12180
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21088 11280 21140 11286
rect 21088 11222 21140 11228
rect 21192 11082 21220 11290
rect 21916 11280 21968 11286
rect 21916 11222 21968 11228
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21376 10606 21404 10950
rect 21928 10810 21956 11222
rect 22112 11218 22140 14350
rect 22468 13184 22520 13190
rect 22468 13126 22520 13132
rect 22480 12986 22508 13126
rect 22468 12980 22520 12986
rect 22468 12922 22520 12928
rect 22664 12782 22692 15982
rect 22940 15366 22968 16934
rect 23124 16726 23152 17138
rect 23308 16998 23336 17870
rect 23676 17678 23704 18362
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 23664 17672 23716 17678
rect 23664 17614 23716 17620
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23400 17202 23428 17478
rect 23388 17196 23440 17202
rect 23388 17138 23440 17144
rect 23296 16992 23348 16998
rect 23296 16934 23348 16940
rect 23400 16794 23428 17138
rect 23756 17128 23808 17134
rect 23478 17096 23534 17105
rect 23756 17070 23808 17076
rect 23478 17031 23480 17040
rect 23532 17031 23534 17040
rect 23480 17002 23532 17008
rect 23388 16788 23440 16794
rect 23388 16730 23440 16736
rect 23112 16720 23164 16726
rect 23112 16662 23164 16668
rect 23572 16584 23624 16590
rect 23572 16526 23624 16532
rect 23584 16250 23612 16526
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23572 15632 23624 15638
rect 23572 15574 23624 15580
rect 23388 15428 23440 15434
rect 23388 15370 23440 15376
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22652 12776 22704 12782
rect 22652 12718 22704 12724
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22652 11212 22704 11218
rect 22652 11154 22704 11160
rect 21916 10804 21968 10810
rect 21916 10746 21968 10752
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 20996 10532 21048 10538
rect 20996 10474 21048 10480
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20444 8424 20496 8430
rect 20548 8412 20576 9386
rect 20640 8974 20668 9522
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20810 8936 20866 8945
rect 20810 8871 20866 8880
rect 20824 8838 20852 8871
rect 20812 8832 20864 8838
rect 20812 8774 20864 8780
rect 20628 8560 20680 8566
rect 20680 8520 20852 8548
rect 20628 8502 20680 8508
rect 20628 8424 20680 8430
rect 20548 8384 20628 8412
rect 20444 8366 20496 8372
rect 20628 8366 20680 8372
rect 20456 8242 20484 8366
rect 20456 8214 20576 8242
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20272 6798 20300 7278
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19432 5568 19484 5574
rect 19432 5510 19484 5516
rect 19444 5302 19472 5510
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19340 4616 19392 4622
rect 19340 4558 19392 4564
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19156 4004 19208 4010
rect 19156 3946 19208 3952
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 19260 800 19288 4490
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19996 4264 20024 5714
rect 20272 4826 20300 6734
rect 20456 5710 20484 7754
rect 20548 6746 20576 8214
rect 20640 6866 20668 8366
rect 20824 8090 20852 8520
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 20916 8022 20944 9522
rect 21192 9518 21220 9998
rect 21376 9926 21404 10542
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21560 10130 21588 10202
rect 21548 10124 21600 10130
rect 21548 10066 21600 10072
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 21560 9178 21588 10066
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21928 9178 21956 9522
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21836 8634 21864 8978
rect 21824 8628 21876 8634
rect 21824 8570 21876 8576
rect 21928 8378 21956 9114
rect 21836 8350 21956 8378
rect 21836 8090 21864 8350
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 20904 8016 20956 8022
rect 20904 7958 20956 7964
rect 21928 7886 21956 8230
rect 21916 7880 21968 7886
rect 21916 7822 21968 7828
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21836 7546 21864 7686
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 20996 7404 21048 7410
rect 20996 7346 21048 7352
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20548 6718 20668 6746
rect 20640 5846 20668 6718
rect 21008 6390 21036 7346
rect 21192 6798 21220 7482
rect 21180 6792 21232 6798
rect 21180 6734 21232 6740
rect 20996 6384 21048 6390
rect 20996 6326 21048 6332
rect 20536 5840 20588 5846
rect 20536 5782 20588 5788
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20456 5370 20484 5646
rect 20548 5370 20576 5782
rect 20640 5642 20668 5782
rect 20628 5636 20680 5642
rect 20628 5578 20680 5584
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20272 4282 20300 4762
rect 22020 4758 22048 10746
rect 22100 8832 22152 8838
rect 22100 8774 22152 8780
rect 22112 8498 22140 8774
rect 22664 8498 22692 11154
rect 22940 10810 22968 15302
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 23308 14074 23336 14282
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23400 13938 23428 15370
rect 23388 13932 23440 13938
rect 23388 13874 23440 13880
rect 23400 13462 23428 13874
rect 23388 13456 23440 13462
rect 23388 13398 23440 13404
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 22928 10804 22980 10810
rect 22928 10746 22980 10752
rect 22100 8492 22152 8498
rect 22652 8492 22704 8498
rect 22152 8452 22324 8480
rect 22100 8434 22152 8440
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22112 7342 22140 7754
rect 22204 7478 22232 7822
rect 22296 7478 22324 8452
rect 22652 8434 22704 8440
rect 22664 8090 22692 8434
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 22652 8084 22704 8090
rect 22652 8026 22704 8032
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22192 7472 22244 7478
rect 22192 7414 22244 7420
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 22204 7002 22232 7414
rect 22480 7342 22508 7890
rect 23032 7478 23060 8230
rect 23020 7472 23072 7478
rect 23020 7414 23072 7420
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 22192 6996 22244 7002
rect 22192 6938 22244 6944
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22204 6254 22232 6734
rect 22192 6248 22244 6254
rect 22192 6190 22244 6196
rect 22008 4752 22060 4758
rect 22008 4694 22060 4700
rect 22480 4690 22508 7278
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23032 6390 23060 6598
rect 23020 6384 23072 6390
rect 23020 6326 23072 6332
rect 23124 5778 23152 12718
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 23308 11354 23336 11630
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23492 10742 23520 12174
rect 23584 11286 23612 15574
rect 23768 15502 23796 17070
rect 24044 16998 24072 18022
rect 24492 17264 24544 17270
rect 24492 17206 24544 17212
rect 24032 16992 24084 16998
rect 24032 16934 24084 16940
rect 24044 15706 24072 16934
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23676 15094 23704 15302
rect 23664 15088 23716 15094
rect 23664 15030 23716 15036
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23676 14074 23704 14350
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23768 12238 23796 15438
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24228 14618 24256 14962
rect 24504 14822 24532 17206
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24596 16522 24624 17070
rect 24860 16584 24912 16590
rect 24860 16526 24912 16532
rect 24584 16516 24636 16522
rect 24584 16458 24636 16464
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24676 15972 24728 15978
rect 24676 15914 24728 15920
rect 24492 14816 24544 14822
rect 24492 14758 24544 14764
rect 24216 14612 24268 14618
rect 24216 14554 24268 14560
rect 24688 14550 24716 15914
rect 24676 14544 24728 14550
rect 24676 14486 24728 14492
rect 24780 14482 24808 16050
rect 24872 15434 24900 16526
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24768 14476 24820 14482
rect 24768 14418 24820 14424
rect 24964 13258 24992 18226
rect 25044 18216 25096 18222
rect 25044 18158 25096 18164
rect 25056 17202 25084 18158
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 25148 16658 25176 17614
rect 25424 17066 25452 18702
rect 26252 18698 26280 19110
rect 26436 18902 26464 20470
rect 26424 18896 26476 18902
rect 26424 18838 26476 18844
rect 26240 18692 26292 18698
rect 26240 18634 26292 18640
rect 25688 18624 25740 18630
rect 25688 18566 25740 18572
rect 25700 17678 25728 18566
rect 26252 18290 26280 18634
rect 26332 18420 26384 18426
rect 26332 18362 26384 18368
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 26344 18154 26372 18362
rect 26332 18148 26384 18154
rect 26332 18090 26384 18096
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 25884 17746 25912 18022
rect 25872 17740 25924 17746
rect 25872 17682 25924 17688
rect 25688 17672 25740 17678
rect 25688 17614 25740 17620
rect 26240 17604 26292 17610
rect 26240 17546 26292 17552
rect 25412 17060 25464 17066
rect 25412 17002 25464 17008
rect 25136 16652 25188 16658
rect 25136 16594 25188 16600
rect 25044 16516 25096 16522
rect 25044 16458 25096 16464
rect 24952 13252 25004 13258
rect 24952 13194 25004 13200
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24872 12782 24900 12922
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24412 11762 24440 12038
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 24492 11076 24544 11082
rect 24492 11018 24544 11024
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 24136 9382 24164 10066
rect 24504 9518 24532 11018
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24596 9654 24624 9998
rect 24584 9648 24636 9654
rect 24584 9590 24636 9596
rect 24492 9512 24544 9518
rect 24492 9454 24544 9460
rect 24124 9376 24176 9382
rect 24124 9318 24176 9324
rect 23480 8900 23532 8906
rect 23480 8842 23532 8848
rect 23492 8498 23520 8842
rect 23296 8492 23348 8498
rect 23480 8492 23532 8498
rect 23348 8452 23428 8480
rect 23296 8434 23348 8440
rect 23400 7886 23428 8452
rect 23480 8434 23532 8440
rect 23492 7886 23520 8434
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23204 6792 23256 6798
rect 23204 6734 23256 6740
rect 23216 6254 23244 6734
rect 23400 6662 23428 7822
rect 23848 6996 23900 7002
rect 23584 6956 23848 6984
rect 23584 6730 23612 6956
rect 23848 6938 23900 6944
rect 24032 6792 24084 6798
rect 23952 6740 24032 6746
rect 23952 6734 24084 6740
rect 23572 6724 23624 6730
rect 23572 6666 23624 6672
rect 23952 6718 24072 6734
rect 23388 6656 23440 6662
rect 23388 6598 23440 6604
rect 23584 6322 23612 6666
rect 23952 6662 23980 6718
rect 23940 6656 23992 6662
rect 23940 6598 23992 6604
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23204 6248 23256 6254
rect 23204 6190 23256 6196
rect 23112 5772 23164 5778
rect 23112 5714 23164 5720
rect 22560 5568 22612 5574
rect 22560 5510 22612 5516
rect 22572 5234 22600 5510
rect 22560 5228 22612 5234
rect 22560 5170 22612 5176
rect 23124 5166 23152 5714
rect 23952 5642 23980 6598
rect 24136 5710 24164 9318
rect 24400 8356 24452 8362
rect 24400 8298 24452 8304
rect 24412 7886 24440 8298
rect 24688 8090 24716 12174
rect 24872 11150 24900 12718
rect 24964 12646 24992 13194
rect 24952 12640 25004 12646
rect 24952 12582 25004 12588
rect 24964 11762 24992 12582
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 25056 11694 25084 16458
rect 25424 16250 25452 17002
rect 26148 16448 26200 16454
rect 26148 16390 26200 16396
rect 26160 16250 26188 16390
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26160 15570 26188 16186
rect 26148 15564 26200 15570
rect 26148 15506 26200 15512
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25320 13932 25372 13938
rect 25320 13874 25372 13880
rect 25332 12918 25360 13874
rect 25700 13870 25728 15302
rect 26252 15162 26280 17546
rect 26424 17128 26476 17134
rect 26424 17070 26476 17076
rect 26436 16794 26464 17070
rect 26424 16788 26476 16794
rect 26424 16730 26476 16736
rect 26240 15156 26292 15162
rect 26240 15098 26292 15104
rect 26804 15026 26832 22510
rect 27172 21690 27200 23666
rect 27448 23644 27476 26522
rect 29012 26382 29040 27270
rect 29380 26518 29408 27474
rect 29552 27056 29604 27062
rect 29552 26998 29604 27004
rect 29368 26512 29420 26518
rect 29368 26454 29420 26460
rect 29000 26376 29052 26382
rect 29000 26318 29052 26324
rect 27528 25764 27580 25770
rect 27528 25706 27580 25712
rect 27540 23798 27568 25706
rect 27712 25152 27764 25158
rect 27712 25094 27764 25100
rect 27724 24682 27752 25094
rect 29000 24948 29052 24954
rect 29000 24890 29052 24896
rect 28172 24744 28224 24750
rect 28172 24686 28224 24692
rect 28724 24744 28776 24750
rect 28724 24686 28776 24692
rect 27712 24676 27764 24682
rect 27712 24618 27764 24624
rect 27528 23792 27580 23798
rect 27528 23734 27580 23740
rect 27448 23616 27568 23644
rect 27344 22976 27396 22982
rect 27344 22918 27396 22924
rect 27356 22778 27384 22918
rect 27344 22772 27396 22778
rect 27344 22714 27396 22720
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27448 22234 27476 22714
rect 27436 22228 27488 22234
rect 27436 22170 27488 22176
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 27172 19922 27200 21490
rect 27344 20392 27396 20398
rect 27344 20334 27396 20340
rect 27356 20058 27384 20334
rect 27344 20052 27396 20058
rect 27344 19994 27396 20000
rect 27160 19916 27212 19922
rect 27160 19858 27212 19864
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 27252 18896 27304 18902
rect 27252 18838 27304 18844
rect 27068 18828 27120 18834
rect 27068 18770 27120 18776
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26988 17202 27016 18158
rect 26976 17196 27028 17202
rect 26976 17138 27028 17144
rect 27080 16046 27108 18770
rect 27264 18766 27292 18838
rect 27252 18760 27304 18766
rect 27252 18702 27304 18708
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27172 17610 27200 18226
rect 27264 17814 27292 18702
rect 27252 17808 27304 17814
rect 27252 17750 27304 17756
rect 27160 17604 27212 17610
rect 27160 17546 27212 17552
rect 27068 16040 27120 16046
rect 27068 15982 27120 15988
rect 27080 15162 27108 15982
rect 27356 15162 27384 19858
rect 27540 18154 27568 23616
rect 27724 23118 27752 24618
rect 28184 24138 28212 24686
rect 28736 24206 28764 24686
rect 29012 24614 29040 24890
rect 29184 24880 29236 24886
rect 29184 24822 29236 24828
rect 29092 24812 29144 24818
rect 29092 24754 29144 24760
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 29104 24410 29132 24754
rect 29196 24410 29224 24822
rect 29276 24812 29328 24818
rect 29276 24754 29328 24760
rect 29092 24404 29144 24410
rect 29092 24346 29144 24352
rect 29184 24404 29236 24410
rect 29184 24346 29236 24352
rect 28816 24268 28868 24274
rect 28816 24210 28868 24216
rect 28724 24200 28776 24206
rect 28724 24142 28776 24148
rect 28172 24132 28224 24138
rect 28172 24074 28224 24080
rect 28184 23322 28212 24074
rect 28828 23662 28856 24210
rect 29104 23730 29132 24346
rect 29288 23730 29316 24754
rect 29092 23724 29144 23730
rect 29092 23666 29144 23672
rect 29276 23724 29328 23730
rect 29276 23666 29328 23672
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 28264 23520 28316 23526
rect 28264 23462 28316 23468
rect 28172 23316 28224 23322
rect 28172 23258 28224 23264
rect 27712 23112 27764 23118
rect 27712 23054 27764 23060
rect 27804 22976 27856 22982
rect 27804 22918 27856 22924
rect 27816 22710 27844 22918
rect 27804 22704 27856 22710
rect 27804 22646 27856 22652
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 27816 21350 27844 21490
rect 27804 21344 27856 21350
rect 27804 21286 27856 21292
rect 27816 20262 27844 21286
rect 28276 20602 28304 23462
rect 29288 23322 29316 23666
rect 29276 23316 29328 23322
rect 29276 23258 29328 23264
rect 28356 23112 28408 23118
rect 28356 23054 28408 23060
rect 28264 20596 28316 20602
rect 28264 20538 28316 20544
rect 27804 20256 27856 20262
rect 27804 20198 27856 20204
rect 27816 18970 27844 20198
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 27528 18148 27580 18154
rect 27528 18090 27580 18096
rect 27724 17338 28028 17354
rect 27712 17332 28040 17338
rect 27764 17326 27988 17332
rect 27712 17274 27764 17280
rect 27988 17274 28040 17280
rect 28080 17196 28132 17202
rect 28080 17138 28132 17144
rect 27712 16584 27764 16590
rect 27712 16526 27764 16532
rect 27724 16250 27752 16526
rect 27712 16244 27764 16250
rect 27712 16186 27764 16192
rect 28092 15978 28120 17138
rect 28080 15972 28132 15978
rect 28080 15914 28132 15920
rect 28264 15904 28316 15910
rect 28264 15846 28316 15852
rect 28276 15706 28304 15846
rect 28080 15700 28132 15706
rect 28080 15642 28132 15648
rect 28264 15700 28316 15706
rect 28264 15642 28316 15648
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 27252 15156 27304 15162
rect 27252 15098 27304 15104
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 26792 15020 26844 15026
rect 26792 14962 26844 14968
rect 26516 14952 26568 14958
rect 26516 14894 26568 14900
rect 26528 14346 26556 14894
rect 26804 14618 26832 14962
rect 26792 14612 26844 14618
rect 26792 14554 26844 14560
rect 26516 14340 26568 14346
rect 26516 14282 26568 14288
rect 26424 14272 26476 14278
rect 26424 14214 26476 14220
rect 26436 14074 26464 14214
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26330 13968 26386 13977
rect 26330 13903 26386 13912
rect 26344 13870 26372 13903
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 25320 12912 25372 12918
rect 25320 12854 25372 12860
rect 25228 12232 25280 12238
rect 25228 12174 25280 12180
rect 25240 11830 25268 12174
rect 25332 11898 25360 12854
rect 25596 12776 25648 12782
rect 25596 12718 25648 12724
rect 25608 12238 25636 12718
rect 25700 12714 25728 13806
rect 26148 13184 26200 13190
rect 26148 13126 26200 13132
rect 26160 12918 26188 13126
rect 26344 12986 26372 13806
rect 26436 13462 26464 14010
rect 26528 13938 26556 14282
rect 26516 13932 26568 13938
rect 26516 13874 26568 13880
rect 26424 13456 26476 13462
rect 26424 13398 26476 13404
rect 26332 12980 26384 12986
rect 26332 12922 26384 12928
rect 26148 12912 26200 12918
rect 26148 12854 26200 12860
rect 26436 12850 26464 13398
rect 26528 12850 26556 13874
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 26424 12844 26476 12850
rect 26424 12786 26476 12792
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 25688 12708 25740 12714
rect 25688 12650 25740 12656
rect 25596 12232 25648 12238
rect 25596 12174 25648 12180
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25044 11688 25096 11694
rect 25044 11630 25096 11636
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 25056 10470 25084 11630
rect 25240 11218 25268 11766
rect 25228 11212 25280 11218
rect 25228 11154 25280 11160
rect 26160 10606 26188 12174
rect 26252 11762 26280 12786
rect 26804 12434 26832 14554
rect 27068 13796 27120 13802
rect 27068 13738 27120 13744
rect 27080 12782 27108 13738
rect 27068 12776 27120 12782
rect 27068 12718 27120 12724
rect 27080 12434 27108 12718
rect 26804 12406 26924 12434
rect 27080 12406 27200 12434
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 26240 11756 26292 11762
rect 26240 11698 26292 11704
rect 26252 11336 26280 11698
rect 26620 11626 26648 12174
rect 26608 11620 26660 11626
rect 26608 11562 26660 11568
rect 26252 11308 26372 11336
rect 26344 11218 26372 11308
rect 26804 11286 26832 12174
rect 26896 11898 26924 12406
rect 26884 11892 26936 11898
rect 26884 11834 26936 11840
rect 26976 11756 27028 11762
rect 26976 11698 27028 11704
rect 26792 11280 26844 11286
rect 26792 11222 26844 11228
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 25964 10600 26016 10606
rect 25964 10542 26016 10548
rect 26148 10600 26200 10606
rect 26148 10542 26200 10548
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24676 8084 24728 8090
rect 24676 8026 24728 8032
rect 24400 7880 24452 7886
rect 24400 7822 24452 7828
rect 24688 7410 24716 8026
rect 24676 7404 24728 7410
rect 24676 7346 24728 7352
rect 24780 7342 24808 9862
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 24768 7336 24820 7342
rect 24768 7278 24820 7284
rect 24964 6662 24992 8366
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 24964 5846 24992 6598
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 24124 5704 24176 5710
rect 24124 5646 24176 5652
rect 23940 5636 23992 5642
rect 23940 5578 23992 5584
rect 23112 5160 23164 5166
rect 23112 5102 23164 5108
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 22468 4684 22520 4690
rect 22468 4626 22520 4632
rect 22756 4622 22784 4966
rect 21088 4616 21140 4622
rect 21088 4558 21140 4564
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 19904 4236 20024 4264
rect 20260 4276 20312 4282
rect 19904 4078 19932 4236
rect 20260 4218 20312 4224
rect 21008 4146 21036 4422
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 19892 4072 19944 4078
rect 19892 4014 19944 4020
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 19352 1442 19380 3538
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19996 3194 20024 4082
rect 21100 4026 21128 4558
rect 23768 4146 23796 4966
rect 24136 4826 24164 5646
rect 24584 5024 24636 5030
rect 24584 4966 24636 4972
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24596 4622 24624 4966
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 24952 4480 25004 4486
rect 24952 4422 25004 4428
rect 24964 4146 24992 4422
rect 25056 4214 25084 10406
rect 25976 10266 26004 10542
rect 26252 10266 26280 11086
rect 26988 10674 27016 11698
rect 26424 10668 26476 10674
rect 26424 10610 26476 10616
rect 26976 10668 27028 10674
rect 26976 10610 27028 10616
rect 25964 10260 26016 10266
rect 25964 10202 26016 10208
rect 26240 10260 26292 10266
rect 26240 10202 26292 10208
rect 25976 9722 26004 10202
rect 26436 10062 26464 10610
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26332 9988 26384 9994
rect 26332 9930 26384 9936
rect 25964 9716 26016 9722
rect 25964 9658 26016 9664
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25320 9036 25372 9042
rect 25320 8978 25372 8984
rect 25332 8498 25360 8978
rect 25412 8968 25464 8974
rect 25412 8910 25464 8916
rect 25320 8492 25372 8498
rect 25320 8434 25372 8440
rect 25332 8090 25360 8434
rect 25424 8294 25452 8910
rect 25792 8634 25820 9522
rect 26240 9512 26292 9518
rect 26240 9454 26292 9460
rect 26252 9042 26280 9454
rect 26240 9036 26292 9042
rect 26240 8978 26292 8984
rect 26344 8634 26372 9930
rect 27068 9444 27120 9450
rect 27068 9386 27120 9392
rect 26424 9376 26476 9382
rect 26424 9318 26476 9324
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 26332 8628 26384 8634
rect 26332 8570 26384 8576
rect 26332 8492 26384 8498
rect 26332 8434 26384 8440
rect 25780 8424 25832 8430
rect 25780 8366 25832 8372
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25320 8084 25372 8090
rect 25320 8026 25372 8032
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 25240 6798 25268 7346
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 25228 6656 25280 6662
rect 25228 6598 25280 6604
rect 25240 6322 25268 6598
rect 25228 6316 25280 6322
rect 25228 6258 25280 6264
rect 25424 5234 25452 8230
rect 25792 8090 25820 8366
rect 25780 8084 25832 8090
rect 25780 8026 25832 8032
rect 25792 7818 25820 8026
rect 26344 8022 26372 8434
rect 26436 8362 26464 9318
rect 27080 9110 27108 9386
rect 27068 9104 27120 9110
rect 27068 9046 27120 9052
rect 26424 8356 26476 8362
rect 26424 8298 26476 8304
rect 26240 8016 26292 8022
rect 26240 7958 26292 7964
rect 26332 8016 26384 8022
rect 26332 7958 26384 7964
rect 25780 7812 25832 7818
rect 25780 7754 25832 7760
rect 26252 7274 26280 7958
rect 26240 7268 26292 7274
rect 26240 7210 26292 7216
rect 26056 6656 26108 6662
rect 26056 6598 26108 6604
rect 26068 5710 26096 6598
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 26252 5914 26280 6054
rect 26240 5908 26292 5914
rect 26240 5850 26292 5856
rect 26056 5704 26108 5710
rect 26056 5646 26108 5652
rect 26344 5302 26372 7958
rect 26436 7750 26464 8298
rect 27172 7834 27200 12406
rect 27264 8430 27292 15098
rect 27528 15088 27580 15094
rect 27528 15030 27580 15036
rect 27344 14816 27396 14822
rect 27344 14758 27396 14764
rect 27252 8424 27304 8430
rect 27252 8366 27304 8372
rect 27356 7954 27384 14758
rect 27436 14272 27488 14278
rect 27436 14214 27488 14220
rect 27448 13870 27476 14214
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27540 13394 27568 15030
rect 28092 15026 28120 15642
rect 28172 15564 28224 15570
rect 28172 15506 28224 15512
rect 28184 15366 28212 15506
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 28080 15020 28132 15026
rect 28080 14962 28132 14968
rect 28184 14550 28212 15302
rect 28368 15042 28396 23054
rect 29380 22098 29408 26454
rect 29564 26382 29592 26998
rect 29552 26376 29604 26382
rect 29552 26318 29604 26324
rect 29552 24608 29604 24614
rect 29552 24550 29604 24556
rect 29564 23118 29592 24550
rect 29552 23112 29604 23118
rect 29552 23054 29604 23060
rect 29368 22092 29420 22098
rect 29656 22094 29684 27950
rect 30288 27940 30340 27946
rect 30288 27882 30340 27888
rect 30300 27402 30328 27882
rect 30288 27396 30340 27402
rect 30288 27338 30340 27344
rect 30012 25356 30064 25362
rect 30012 25298 30064 25304
rect 29920 25288 29972 25294
rect 29920 25230 29972 25236
rect 29736 24812 29788 24818
rect 29736 24754 29788 24760
rect 29748 24614 29776 24754
rect 29932 24682 29960 25230
rect 29920 24676 29972 24682
rect 29920 24618 29972 24624
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29932 23730 29960 24618
rect 29920 23724 29972 23730
rect 29920 23666 29972 23672
rect 29828 23588 29880 23594
rect 29828 23530 29880 23536
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 29368 22034 29420 22040
rect 29564 22066 29684 22094
rect 28448 21412 28500 21418
rect 28448 21354 28500 21360
rect 28460 21146 28488 21354
rect 28540 21344 28592 21350
rect 28540 21286 28592 21292
rect 28448 21140 28500 21146
rect 28448 21082 28500 21088
rect 28448 20936 28500 20942
rect 28448 20878 28500 20884
rect 28460 20262 28488 20878
rect 28552 20874 28580 21286
rect 29564 21010 29592 22066
rect 29644 22024 29696 22030
rect 29644 21966 29696 21972
rect 29656 21554 29684 21966
rect 29644 21548 29696 21554
rect 29644 21490 29696 21496
rect 29552 21004 29604 21010
rect 29552 20946 29604 20952
rect 28540 20868 28592 20874
rect 28540 20810 28592 20816
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29380 20602 29408 20742
rect 29656 20618 29684 21490
rect 29748 21434 29776 23054
rect 29840 23050 29868 23530
rect 29920 23520 29972 23526
rect 29920 23462 29972 23468
rect 29932 23118 29960 23462
rect 29920 23112 29972 23118
rect 29920 23054 29972 23060
rect 29828 23044 29880 23050
rect 29828 22986 29880 22992
rect 29840 22030 29868 22986
rect 29920 22636 29972 22642
rect 30024 22624 30052 25298
rect 30300 24206 30328 27338
rect 30944 27062 30972 27950
rect 31036 27606 31064 27950
rect 31024 27600 31076 27606
rect 31024 27542 31076 27548
rect 30932 27056 30984 27062
rect 30932 26998 30984 27004
rect 31128 26450 31156 33322
rect 32416 32910 32444 33594
rect 34520 33516 34572 33522
rect 34520 33458 34572 33464
rect 35348 33516 35400 33522
rect 35348 33458 35400 33464
rect 34532 33318 34560 33458
rect 34520 33312 34572 33318
rect 34520 33254 34572 33260
rect 33140 32972 33192 32978
rect 33140 32914 33192 32920
rect 32404 32904 32456 32910
rect 32404 32846 32456 32852
rect 31484 31748 31536 31754
rect 31484 31690 31536 31696
rect 31496 31482 31524 31690
rect 32312 31680 32364 31686
rect 32312 31622 32364 31628
rect 31484 31476 31536 31482
rect 31484 31418 31536 31424
rect 32324 31278 32352 31622
rect 32312 31272 32364 31278
rect 32312 31214 32364 31220
rect 32680 31272 32732 31278
rect 32680 31214 32732 31220
rect 31944 31204 31996 31210
rect 31944 31146 31996 31152
rect 31300 30932 31352 30938
rect 31300 30874 31352 30880
rect 31312 28626 31340 30874
rect 31956 30734 31984 31146
rect 31944 30728 31996 30734
rect 31944 30670 31996 30676
rect 31392 29504 31444 29510
rect 31392 29446 31444 29452
rect 31300 28620 31352 28626
rect 31300 28562 31352 28568
rect 31404 28422 31432 29446
rect 31956 29238 31984 30670
rect 32036 30660 32088 30666
rect 32036 30602 32088 30608
rect 32048 30394 32076 30602
rect 32036 30388 32088 30394
rect 32036 30330 32088 30336
rect 31944 29232 31996 29238
rect 31944 29174 31996 29180
rect 31668 29096 31720 29102
rect 31668 29038 31720 29044
rect 31484 28620 31536 28626
rect 31484 28562 31536 28568
rect 31392 28416 31444 28422
rect 31392 28358 31444 28364
rect 31300 28212 31352 28218
rect 31300 28154 31352 28160
rect 31208 27940 31260 27946
rect 31208 27882 31260 27888
rect 31220 27538 31248 27882
rect 31312 27674 31340 28154
rect 31300 27668 31352 27674
rect 31300 27610 31352 27616
rect 31208 27532 31260 27538
rect 31208 27474 31260 27480
rect 31300 27464 31352 27470
rect 31300 27406 31352 27412
rect 31116 26444 31168 26450
rect 31116 26386 31168 26392
rect 30748 26308 30800 26314
rect 30748 26250 30800 26256
rect 30380 24336 30432 24342
rect 30380 24278 30432 24284
rect 30288 24200 30340 24206
rect 30288 24142 30340 24148
rect 30104 24064 30156 24070
rect 30104 24006 30156 24012
rect 30116 23118 30144 24006
rect 30288 23724 30340 23730
rect 30288 23666 30340 23672
rect 30104 23112 30156 23118
rect 30104 23054 30156 23060
rect 30116 22642 30144 23054
rect 30196 22976 30248 22982
rect 30196 22918 30248 22924
rect 29972 22596 30052 22624
rect 30104 22636 30156 22642
rect 29920 22578 29972 22584
rect 30104 22578 30156 22584
rect 30208 22098 30236 22918
rect 30300 22778 30328 23666
rect 30392 23662 30420 24278
rect 30760 23730 30788 26250
rect 31208 25152 31260 25158
rect 31208 25094 31260 25100
rect 30840 24404 30892 24410
rect 30840 24346 30892 24352
rect 30852 23730 30880 24346
rect 30748 23724 30800 23730
rect 30748 23666 30800 23672
rect 30840 23724 30892 23730
rect 30840 23666 30892 23672
rect 30380 23656 30432 23662
rect 30380 23598 30432 23604
rect 30392 23186 30420 23598
rect 30760 23526 30788 23666
rect 30748 23520 30800 23526
rect 30748 23462 30800 23468
rect 30852 23254 30880 23666
rect 30840 23248 30892 23254
rect 30840 23190 30892 23196
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 31220 23050 31248 25094
rect 31208 23044 31260 23050
rect 31208 22986 31260 22992
rect 30288 22772 30340 22778
rect 30288 22714 30340 22720
rect 30288 22568 30340 22574
rect 30288 22510 30340 22516
rect 29920 22092 29972 22098
rect 29920 22034 29972 22040
rect 30196 22092 30248 22098
rect 30196 22034 30248 22040
rect 29828 22024 29880 22030
rect 29828 21966 29880 21972
rect 29840 21622 29868 21966
rect 29932 21690 29960 22034
rect 30300 21690 30328 22510
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 30288 21684 30340 21690
rect 30288 21626 30340 21632
rect 30380 21684 30432 21690
rect 30380 21626 30432 21632
rect 29828 21616 29880 21622
rect 29828 21558 29880 21564
rect 29920 21548 29972 21554
rect 29920 21490 29972 21496
rect 29932 21434 29960 21490
rect 29748 21406 29960 21434
rect 29932 21146 29960 21406
rect 29920 21140 29972 21146
rect 29920 21082 29972 21088
rect 30104 20936 30156 20942
rect 30104 20878 30156 20884
rect 29368 20596 29420 20602
rect 29656 20590 29868 20618
rect 29368 20538 29420 20544
rect 28448 20256 28500 20262
rect 28448 20198 28500 20204
rect 29276 19916 29328 19922
rect 29276 19858 29328 19864
rect 29184 18692 29236 18698
rect 29184 18634 29236 18640
rect 29196 18426 29224 18634
rect 29184 18420 29236 18426
rect 29184 18362 29236 18368
rect 28908 15904 28960 15910
rect 28908 15846 28960 15852
rect 28920 15706 28948 15846
rect 28908 15700 28960 15706
rect 28908 15642 28960 15648
rect 28540 15360 28592 15366
rect 28540 15302 28592 15308
rect 28276 15026 28396 15042
rect 28552 15026 28580 15302
rect 28264 15020 28396 15026
rect 28316 15014 28396 15020
rect 28264 14962 28316 14968
rect 28368 14618 28396 15014
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 28356 14612 28408 14618
rect 28356 14554 28408 14560
rect 28172 14544 28224 14550
rect 28172 14486 28224 14492
rect 27528 13388 27580 13394
rect 27528 13330 27580 13336
rect 28080 13388 28132 13394
rect 28080 13330 28132 13336
rect 27712 13320 27764 13326
rect 27712 13262 27764 13268
rect 27724 12986 27752 13262
rect 27712 12980 27764 12986
rect 27712 12922 27764 12928
rect 27436 12708 27488 12714
rect 27436 12650 27488 12656
rect 27448 11762 27476 12650
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 28092 11218 28120 13330
rect 28816 12708 28868 12714
rect 28816 12650 28868 12656
rect 28828 11694 28856 12650
rect 29288 12442 29316 19858
rect 29380 18970 29408 20538
rect 29644 20460 29696 20466
rect 29644 20402 29696 20408
rect 29656 18970 29684 20402
rect 29840 20398 29868 20590
rect 30116 20466 30144 20878
rect 30288 20868 30340 20874
rect 30288 20810 30340 20816
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 29828 20392 29880 20398
rect 29828 20334 29880 20340
rect 29840 19922 29868 20334
rect 29828 19916 29880 19922
rect 29828 19858 29880 19864
rect 30116 19854 30144 20402
rect 30104 19848 30156 19854
rect 30104 19790 30156 19796
rect 29368 18964 29420 18970
rect 29368 18906 29420 18912
rect 29644 18964 29696 18970
rect 29644 18906 29696 18912
rect 30116 18902 30144 19790
rect 30104 18896 30156 18902
rect 30104 18838 30156 18844
rect 30196 18624 30248 18630
rect 30196 18566 30248 18572
rect 29460 16584 29512 16590
rect 29460 16526 29512 16532
rect 29472 16250 29500 16526
rect 29920 16448 29972 16454
rect 29920 16390 29972 16396
rect 29932 16250 29960 16390
rect 29460 16244 29512 16250
rect 29460 16186 29512 16192
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 29828 16108 29880 16114
rect 29828 16050 29880 16056
rect 29368 15496 29420 15502
rect 29368 15438 29420 15444
rect 29380 14414 29408 15438
rect 29552 15360 29604 15366
rect 29552 15302 29604 15308
rect 29460 15020 29512 15026
rect 29460 14962 29512 14968
rect 29472 14618 29500 14962
rect 29564 14958 29592 15302
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29460 14612 29512 14618
rect 29460 14554 29512 14560
rect 29368 14408 29420 14414
rect 29368 14350 29420 14356
rect 29276 12436 29328 12442
rect 29380 12434 29408 14350
rect 29736 14272 29788 14278
rect 29736 14214 29788 14220
rect 29380 12406 29500 12434
rect 29276 12378 29328 12384
rect 28908 11756 28960 11762
rect 28908 11698 28960 11704
rect 28816 11688 28868 11694
rect 28816 11630 28868 11636
rect 28920 11354 28948 11698
rect 29000 11620 29052 11626
rect 29000 11562 29052 11568
rect 29012 11354 29040 11562
rect 28908 11348 28960 11354
rect 28908 11290 28960 11296
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 29472 11286 29500 12406
rect 28264 11280 28316 11286
rect 28264 11222 28316 11228
rect 29460 11280 29512 11286
rect 29460 11222 29512 11228
rect 28080 11212 28132 11218
rect 28080 11154 28132 11160
rect 27988 9512 28040 9518
rect 27988 9454 28040 9460
rect 28000 8906 28028 9454
rect 28092 9178 28120 11154
rect 28172 9988 28224 9994
rect 28172 9930 28224 9936
rect 28080 9172 28132 9178
rect 28080 9114 28132 9120
rect 27988 8900 28040 8906
rect 27988 8842 28040 8848
rect 28000 8786 28028 8842
rect 27908 8758 28028 8786
rect 27344 7948 27396 7954
rect 27344 7890 27396 7896
rect 27436 7880 27488 7886
rect 27172 7806 27384 7834
rect 27436 7822 27488 7828
rect 26424 7744 26476 7750
rect 26424 7686 26476 7692
rect 26424 6996 26476 7002
rect 26424 6938 26476 6944
rect 27160 6996 27212 7002
rect 27160 6938 27212 6944
rect 27252 6996 27304 7002
rect 27252 6938 27304 6944
rect 26436 6798 26464 6938
rect 26424 6792 26476 6798
rect 26424 6734 26476 6740
rect 27172 6730 27200 6938
rect 27160 6724 27212 6730
rect 27160 6666 27212 6672
rect 27264 6662 27292 6938
rect 27356 6866 27384 7806
rect 27448 7002 27476 7822
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 27436 6996 27488 7002
rect 27436 6938 27488 6944
rect 27344 6860 27396 6866
rect 27344 6802 27396 6808
rect 27252 6656 27304 6662
rect 27252 6598 27304 6604
rect 27264 6225 27292 6598
rect 27356 6390 27384 6802
rect 27344 6384 27396 6390
rect 27344 6326 27396 6332
rect 27528 6384 27580 6390
rect 27528 6326 27580 6332
rect 27356 6254 27384 6326
rect 27344 6248 27396 6254
rect 27250 6216 27306 6225
rect 26424 6180 26476 6186
rect 27344 6190 27396 6196
rect 27250 6151 27306 6160
rect 26424 6122 26476 6128
rect 26436 5710 26464 6122
rect 27540 5710 27568 6326
rect 27724 6322 27752 7346
rect 27908 6914 27936 8758
rect 27988 8628 28040 8634
rect 28092 8616 28120 9114
rect 28040 8588 28120 8616
rect 27988 8570 28040 8576
rect 28184 8362 28212 9930
rect 28276 9586 28304 11222
rect 29092 11212 29144 11218
rect 29092 11154 29144 11160
rect 28632 9920 28684 9926
rect 28632 9862 28684 9868
rect 28264 9580 28316 9586
rect 28264 9522 28316 9528
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 28264 8492 28316 8498
rect 28264 8434 28316 8440
rect 28172 8356 28224 8362
rect 28172 8298 28224 8304
rect 28276 8090 28304 8434
rect 28264 8084 28316 8090
rect 28264 8026 28316 8032
rect 28276 7546 28304 8026
rect 28356 7812 28408 7818
rect 28356 7754 28408 7760
rect 28368 7546 28396 7754
rect 28264 7540 28316 7546
rect 28264 7482 28316 7488
rect 28356 7540 28408 7546
rect 28356 7482 28408 7488
rect 27908 6886 28028 6914
rect 28000 6458 28028 6886
rect 27988 6452 28040 6458
rect 27988 6394 28040 6400
rect 28460 6390 28488 8910
rect 28644 8090 28672 9862
rect 29104 9382 29132 11154
rect 29184 11076 29236 11082
rect 29184 11018 29236 11024
rect 29196 10606 29224 11018
rect 29184 10600 29236 10606
rect 29184 10542 29236 10548
rect 29196 10266 29224 10542
rect 29552 10464 29604 10470
rect 29552 10406 29604 10412
rect 29184 10260 29236 10266
rect 29184 10202 29236 10208
rect 29564 10198 29592 10406
rect 29552 10192 29604 10198
rect 29552 10134 29604 10140
rect 29184 10124 29236 10130
rect 29184 10066 29236 10072
rect 29092 9376 29144 9382
rect 29092 9318 29144 9324
rect 29000 8968 29052 8974
rect 29000 8910 29052 8916
rect 29012 8634 29040 8910
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 29104 8498 29132 9318
rect 29092 8492 29144 8498
rect 29092 8434 29144 8440
rect 28632 8084 28684 8090
rect 28632 8026 28684 8032
rect 28816 7540 28868 7546
rect 28816 7482 28868 7488
rect 28632 7336 28684 7342
rect 28632 7278 28684 7284
rect 28644 6866 28672 7278
rect 28632 6860 28684 6866
rect 28632 6802 28684 6808
rect 28448 6384 28500 6390
rect 28448 6326 28500 6332
rect 27712 6316 27764 6322
rect 27712 6258 27764 6264
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 27632 6118 27660 6190
rect 27620 6112 27672 6118
rect 27620 6054 27672 6060
rect 27724 5914 27752 6258
rect 27988 6112 28040 6118
rect 27988 6054 28040 6060
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 26424 5704 26476 5710
rect 26424 5646 26476 5652
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 26332 5296 26384 5302
rect 26332 5238 26384 5244
rect 25412 5228 25464 5234
rect 25412 5170 25464 5176
rect 25780 5228 25832 5234
rect 25780 5170 25832 5176
rect 25044 4208 25096 4214
rect 25044 4150 25096 4156
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 24952 4140 25004 4146
rect 24952 4082 25004 4088
rect 21008 3998 21128 4026
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19812 2922 19840 2994
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19800 2916 19852 2922
rect 19800 2858 19852 2864
rect 19444 1578 19472 2858
rect 19812 2650 19840 2858
rect 19800 2644 19852 2650
rect 19800 2586 19852 2592
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19444 1550 19840 1578
rect 19352 1414 19564 1442
rect 19536 800 19564 1414
rect 19812 800 19840 1550
rect 20088 800 20116 3470
rect 20272 2650 20300 3674
rect 20548 3602 20576 3878
rect 20628 3664 20680 3670
rect 20628 3606 20680 3612
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 20352 2848 20404 2854
rect 20352 2790 20404 2796
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 20364 800 20392 2790
rect 20640 800 20668 3606
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20916 800 20944 2926
rect 21008 800 21036 3998
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 24400 3936 24452 3942
rect 24400 3878 24452 3884
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21100 3194 21128 3470
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 21272 2916 21324 2922
rect 21272 2858 21324 2864
rect 21180 2576 21232 2582
rect 21180 2518 21232 2524
rect 21192 800 21220 2518
rect 21284 800 21312 2858
rect 21456 2848 21508 2854
rect 21456 2790 21508 2796
rect 21468 800 21496 2790
rect 21640 2372 21692 2378
rect 21640 2314 21692 2320
rect 21548 2304 21600 2310
rect 21548 2246 21600 2252
rect 21560 800 21588 2246
rect 21652 2106 21680 2314
rect 21640 2100 21692 2106
rect 21640 2042 21692 2048
rect 21744 800 21772 3878
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 21836 800 21864 2994
rect 22020 800 22048 3470
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22204 800 22232 2450
rect 22480 800 22508 3470
rect 22744 2440 22796 2446
rect 22744 2382 22796 2388
rect 22756 800 22784 2382
rect 23032 800 23060 3878
rect 23952 3534 23980 3878
rect 24412 3602 24440 3878
rect 25792 3738 25820 5170
rect 26344 4282 26372 5238
rect 26332 4276 26384 4282
rect 26332 4218 26384 4224
rect 26436 4010 26464 5646
rect 27540 5234 27568 5646
rect 27528 5228 27580 5234
rect 27528 5170 27580 5176
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 27816 4826 27844 5170
rect 27804 4820 27856 4826
rect 27804 4762 27856 4768
rect 28000 4622 28028 6054
rect 28644 5370 28672 6802
rect 28724 6724 28776 6730
rect 28724 6666 28776 6672
rect 28736 6361 28764 6666
rect 28722 6352 28778 6361
rect 28722 6287 28724 6296
rect 28776 6287 28778 6296
rect 28724 6258 28776 6264
rect 28736 5914 28764 6258
rect 28828 6254 28856 7482
rect 29196 7478 29224 10066
rect 29644 9512 29696 9518
rect 29644 9454 29696 9460
rect 29656 9178 29684 9454
rect 29748 9178 29776 14214
rect 29840 13802 29868 16050
rect 29932 15502 29960 16186
rect 29920 15496 29972 15502
rect 29920 15438 29972 15444
rect 30104 15020 30156 15026
rect 30104 14962 30156 14968
rect 30116 14482 30144 14962
rect 30104 14476 30156 14482
rect 30104 14418 30156 14424
rect 29828 13796 29880 13802
rect 29828 13738 29880 13744
rect 30116 13530 30144 14418
rect 30104 13524 30156 13530
rect 30104 13466 30156 13472
rect 30208 11354 30236 18566
rect 30300 17882 30328 20810
rect 30392 19514 30420 21626
rect 30748 21548 30800 21554
rect 30748 21490 30800 21496
rect 30472 21344 30524 21350
rect 30472 21286 30524 21292
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30288 17876 30340 17882
rect 30288 17818 30340 17824
rect 30196 11348 30248 11354
rect 30196 11290 30248 11296
rect 30484 11150 30512 21286
rect 30760 21146 30788 21490
rect 30748 21140 30800 21146
rect 30748 21082 30800 21088
rect 31312 20602 31340 27406
rect 31404 25242 31432 28358
rect 31496 25430 31524 28562
rect 31680 28218 31708 29038
rect 31668 28212 31720 28218
rect 31668 28154 31720 28160
rect 32324 28082 32352 31214
rect 32692 30938 32720 31214
rect 32680 30932 32732 30938
rect 32680 30874 32732 30880
rect 32588 30592 32640 30598
rect 32588 30534 32640 30540
rect 32600 30326 32628 30534
rect 32588 30320 32640 30326
rect 32588 30262 32640 30268
rect 32496 30252 32548 30258
rect 32496 30194 32548 30200
rect 32508 29850 32536 30194
rect 32496 29844 32548 29850
rect 32496 29786 32548 29792
rect 32600 28558 32628 30262
rect 32692 30190 32720 30874
rect 32680 30184 32732 30190
rect 32680 30126 32732 30132
rect 32588 28552 32640 28558
rect 32588 28494 32640 28500
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 32404 27872 32456 27878
rect 32404 27814 32456 27820
rect 32416 27606 32444 27814
rect 32404 27600 32456 27606
rect 32404 27542 32456 27548
rect 32128 26988 32180 26994
rect 32128 26930 32180 26936
rect 31852 26580 31904 26586
rect 31852 26522 31904 26528
rect 31484 25424 31536 25430
rect 31484 25366 31536 25372
rect 31864 25362 31892 26522
rect 31944 26308 31996 26314
rect 31944 26250 31996 26256
rect 31852 25356 31904 25362
rect 31852 25298 31904 25304
rect 31404 25214 31524 25242
rect 31496 23118 31524 25214
rect 31956 24750 31984 26250
rect 32036 25832 32088 25838
rect 32036 25774 32088 25780
rect 32048 24818 32076 25774
rect 32140 25498 32168 26930
rect 32312 26376 32364 26382
rect 32312 26318 32364 26324
rect 32324 26042 32352 26318
rect 32588 26308 32640 26314
rect 32588 26250 32640 26256
rect 32312 26036 32364 26042
rect 32312 25978 32364 25984
rect 32128 25492 32180 25498
rect 32128 25434 32180 25440
rect 32324 25362 32352 25978
rect 32312 25356 32364 25362
rect 32312 25298 32364 25304
rect 32600 24818 32628 26250
rect 32680 26240 32732 26246
rect 32680 26182 32732 26188
rect 32692 25294 32720 26182
rect 32772 25900 32824 25906
rect 32772 25842 32824 25848
rect 32680 25288 32732 25294
rect 32680 25230 32732 25236
rect 32036 24812 32088 24818
rect 32036 24754 32088 24760
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32588 24812 32640 24818
rect 32588 24754 32640 24760
rect 31944 24744 31996 24750
rect 31944 24686 31996 24692
rect 31956 23798 31984 24686
rect 32036 24268 32088 24274
rect 32036 24210 32088 24216
rect 31944 23792 31996 23798
rect 31944 23734 31996 23740
rect 31944 23656 31996 23662
rect 31944 23598 31996 23604
rect 31576 23588 31628 23594
rect 31576 23530 31628 23536
rect 31588 23186 31616 23530
rect 31576 23180 31628 23186
rect 31576 23122 31628 23128
rect 31484 23112 31536 23118
rect 31484 23054 31536 23060
rect 31956 22778 31984 23598
rect 31944 22772 31996 22778
rect 31944 22714 31996 22720
rect 31760 22636 31812 22642
rect 31760 22578 31812 22584
rect 31484 22500 31536 22506
rect 31484 22442 31536 22448
rect 31496 22098 31524 22442
rect 31484 22092 31536 22098
rect 31484 22034 31536 22040
rect 31772 21978 31800 22578
rect 31944 22024 31996 22030
rect 31772 21962 31892 21978
rect 31944 21966 31996 21972
rect 31772 21956 31904 21962
rect 31772 21950 31852 21956
rect 31852 21898 31904 21904
rect 31864 21418 31892 21898
rect 31956 21418 31984 21966
rect 31852 21412 31904 21418
rect 31852 21354 31904 21360
rect 31944 21412 31996 21418
rect 31944 21354 31996 21360
rect 31864 21078 31892 21354
rect 31852 21072 31904 21078
rect 31852 21014 31904 21020
rect 32048 20890 32076 24210
rect 32220 23724 32272 23730
rect 32220 23666 32272 23672
rect 32232 22778 32260 23666
rect 32324 23662 32352 24754
rect 32312 23656 32364 23662
rect 32312 23598 32364 23604
rect 32784 23118 32812 25842
rect 32956 25492 33008 25498
rect 32956 25434 33008 25440
rect 32864 24064 32916 24070
rect 32864 24006 32916 24012
rect 32772 23112 32824 23118
rect 32772 23054 32824 23060
rect 32404 22976 32456 22982
rect 32404 22918 32456 22924
rect 32220 22772 32272 22778
rect 32220 22714 32272 22720
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 32140 22094 32168 22374
rect 32140 22066 32352 22094
rect 32232 22030 32260 22066
rect 32220 22024 32272 22030
rect 32220 21966 32272 21972
rect 32128 21956 32180 21962
rect 32128 21898 32180 21904
rect 31864 20862 32076 20890
rect 31300 20596 31352 20602
rect 31300 20538 31352 20544
rect 31668 20052 31720 20058
rect 31668 19994 31720 20000
rect 31116 19712 31168 19718
rect 31116 19654 31168 19660
rect 31128 18698 31156 19654
rect 31116 18692 31168 18698
rect 31116 18634 31168 18640
rect 31680 18290 31708 19994
rect 31760 19508 31812 19514
rect 31760 19450 31812 19456
rect 31772 18698 31800 19450
rect 31760 18692 31812 18698
rect 31760 18634 31812 18640
rect 31668 18284 31720 18290
rect 31668 18226 31720 18232
rect 31680 17746 31708 18226
rect 31668 17740 31720 17746
rect 31668 17682 31720 17688
rect 30748 17604 30800 17610
rect 30748 17546 30800 17552
rect 31760 17604 31812 17610
rect 31760 17546 31812 17552
rect 30760 17066 30788 17546
rect 31024 17536 31076 17542
rect 31024 17478 31076 17484
rect 31036 17134 31064 17478
rect 31024 17128 31076 17134
rect 31024 17070 31076 17076
rect 30748 17060 30800 17066
rect 30748 17002 30800 17008
rect 31208 16992 31260 16998
rect 31208 16934 31260 16940
rect 30564 14952 30616 14958
rect 30564 14894 30616 14900
rect 30576 14414 30604 14894
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 30656 11756 30708 11762
rect 30656 11698 30708 11704
rect 30932 11756 30984 11762
rect 30932 11698 30984 11704
rect 31116 11756 31168 11762
rect 31116 11698 31168 11704
rect 30472 11144 30524 11150
rect 30472 11086 30524 11092
rect 30668 10810 30696 11698
rect 30748 11076 30800 11082
rect 30748 11018 30800 11024
rect 30656 10804 30708 10810
rect 30656 10746 30708 10752
rect 30760 10674 30788 11018
rect 30840 10736 30892 10742
rect 30840 10678 30892 10684
rect 30748 10668 30800 10674
rect 30748 10610 30800 10616
rect 30852 10470 30880 10678
rect 30380 10464 30432 10470
rect 30380 10406 30432 10412
rect 30840 10464 30892 10470
rect 30840 10406 30892 10412
rect 30392 10062 30420 10406
rect 30944 10266 30972 11698
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 31128 10062 31156 11698
rect 31220 11150 31248 16934
rect 31772 16726 31800 17546
rect 31760 16720 31812 16726
rect 31760 16662 31812 16668
rect 31864 14958 31892 20862
rect 32036 19372 32088 19378
rect 32036 19314 32088 19320
rect 32048 18426 32076 19314
rect 32036 18420 32088 18426
rect 32036 18362 32088 18368
rect 32036 17672 32088 17678
rect 32036 17614 32088 17620
rect 31944 17536 31996 17542
rect 31944 17478 31996 17484
rect 31956 17202 31984 17478
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 31484 14952 31536 14958
rect 31484 14894 31536 14900
rect 31852 14952 31904 14958
rect 31852 14894 31904 14900
rect 31300 12232 31352 12238
rect 31300 12174 31352 12180
rect 31312 11354 31340 12174
rect 31392 11756 31444 11762
rect 31392 11698 31444 11704
rect 31404 11558 31432 11698
rect 31392 11552 31444 11558
rect 31392 11494 31444 11500
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31208 11144 31260 11150
rect 31208 11086 31260 11092
rect 31220 10266 31248 11086
rect 31208 10260 31260 10266
rect 31208 10202 31260 10208
rect 30380 10056 30432 10062
rect 30380 9998 30432 10004
rect 30656 10056 30708 10062
rect 30656 9998 30708 10004
rect 31116 10056 31168 10062
rect 31116 9998 31168 10004
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 29644 9172 29696 9178
rect 29644 9114 29696 9120
rect 29736 9172 29788 9178
rect 29736 9114 29788 9120
rect 29840 8634 29868 9522
rect 30380 9376 30432 9382
rect 30380 9318 30432 9324
rect 29828 8628 29880 8634
rect 29828 8570 29880 8576
rect 29644 8492 29696 8498
rect 29644 8434 29696 8440
rect 29552 8288 29604 8294
rect 29552 8230 29604 8236
rect 29564 7478 29592 8230
rect 29656 8090 29684 8434
rect 29644 8084 29696 8090
rect 29644 8026 29696 8032
rect 29184 7472 29236 7478
rect 29184 7414 29236 7420
rect 29552 7472 29604 7478
rect 29552 7414 29604 7420
rect 29656 6934 29684 8026
rect 30392 7886 30420 9318
rect 30564 8900 30616 8906
rect 30564 8842 30616 8848
rect 30576 8090 30604 8842
rect 30668 8362 30696 9998
rect 30932 9512 30984 9518
rect 30932 9454 30984 9460
rect 30944 8430 30972 9454
rect 31220 8634 31248 10202
rect 31404 9994 31432 11494
rect 31496 10674 31524 14894
rect 31944 14816 31996 14822
rect 31944 14758 31996 14764
rect 31956 14482 31984 14758
rect 31944 14476 31996 14482
rect 31944 14418 31996 14424
rect 31944 13320 31996 13326
rect 31944 13262 31996 13268
rect 31668 12096 31720 12102
rect 31668 12038 31720 12044
rect 31680 11150 31708 12038
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 31956 10810 31984 13262
rect 32048 12170 32076 17614
rect 32036 12164 32088 12170
rect 32036 12106 32088 12112
rect 32140 11830 32168 21898
rect 32324 21554 32352 22066
rect 32416 22030 32444 22918
rect 32784 22681 32812 23054
rect 32770 22672 32826 22681
rect 32770 22607 32826 22616
rect 32404 22024 32456 22030
rect 32404 21966 32456 21972
rect 32416 21554 32444 21966
rect 32312 21548 32364 21554
rect 32312 21490 32364 21496
rect 32404 21548 32456 21554
rect 32404 21490 32456 21496
rect 32680 21480 32732 21486
rect 32680 21422 32732 21428
rect 32772 21480 32824 21486
rect 32772 21422 32824 21428
rect 32692 21146 32720 21422
rect 32680 21140 32732 21146
rect 32680 21082 32732 21088
rect 32496 21004 32548 21010
rect 32496 20946 32548 20952
rect 32220 20936 32272 20942
rect 32220 20878 32272 20884
rect 32232 20534 32260 20878
rect 32220 20528 32272 20534
rect 32220 20470 32272 20476
rect 32508 20466 32536 20946
rect 32784 20602 32812 21422
rect 32876 21418 32904 24006
rect 32968 23866 32996 25434
rect 33152 25362 33180 32914
rect 33324 32768 33376 32774
rect 33324 32710 33376 32716
rect 33232 26784 33284 26790
rect 33232 26726 33284 26732
rect 33244 25974 33272 26726
rect 33232 25968 33284 25974
rect 33232 25910 33284 25916
rect 33232 25696 33284 25702
rect 33232 25638 33284 25644
rect 33140 25356 33192 25362
rect 33140 25298 33192 25304
rect 33244 25294 33272 25638
rect 33232 25288 33284 25294
rect 33232 25230 33284 25236
rect 33336 24834 33364 32710
rect 34532 32570 34560 33254
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35360 32910 35388 33458
rect 37740 33448 37792 33454
rect 37740 33390 37792 33396
rect 35900 33380 35952 33386
rect 35900 33322 35952 33328
rect 35912 32910 35940 33322
rect 37188 33312 37240 33318
rect 37188 33254 37240 33260
rect 36544 32972 36596 32978
rect 36544 32914 36596 32920
rect 35348 32904 35400 32910
rect 35348 32846 35400 32852
rect 35900 32904 35952 32910
rect 35900 32846 35952 32852
rect 34520 32564 34572 32570
rect 34520 32506 34572 32512
rect 35360 32502 35388 32846
rect 35348 32496 35400 32502
rect 35348 32438 35400 32444
rect 34520 32428 34572 32434
rect 34520 32370 34572 32376
rect 33968 32224 34020 32230
rect 33968 32166 34020 32172
rect 33980 31346 34008 32166
rect 34532 31686 34560 32370
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34520 31680 34572 31686
rect 34520 31622 34572 31628
rect 34532 31482 34560 31622
rect 34520 31476 34572 31482
rect 34520 31418 34572 31424
rect 34716 31414 34744 31758
rect 35360 31482 35388 32438
rect 36556 32434 36584 32914
rect 37200 32910 37228 33254
rect 37188 32904 37240 32910
rect 37188 32846 37240 32852
rect 37200 32434 37228 32846
rect 37752 32434 37780 33390
rect 38660 32972 38712 32978
rect 38660 32914 38712 32920
rect 38292 32904 38344 32910
rect 38292 32846 38344 32852
rect 35808 32428 35860 32434
rect 35808 32370 35860 32376
rect 36544 32428 36596 32434
rect 36544 32370 36596 32376
rect 37188 32428 37240 32434
rect 37188 32370 37240 32376
rect 37740 32428 37792 32434
rect 37740 32370 37792 32376
rect 35532 32360 35584 32366
rect 35532 32302 35584 32308
rect 35348 31476 35400 31482
rect 35348 31418 35400 31424
rect 34704 31408 34756 31414
rect 34704 31350 34756 31356
rect 33968 31340 34020 31346
rect 33968 31282 34020 31288
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35348 29232 35400 29238
rect 35348 29174 35400 29180
rect 34704 29096 34756 29102
rect 34704 29038 34756 29044
rect 33416 28416 33468 28422
rect 33416 28358 33468 28364
rect 33428 28082 33456 28358
rect 33416 28076 33468 28082
rect 33416 28018 33468 28024
rect 33600 27872 33652 27878
rect 33600 27814 33652 27820
rect 33508 25832 33560 25838
rect 33508 25774 33560 25780
rect 33416 25152 33468 25158
rect 33416 25094 33468 25100
rect 33428 24954 33456 25094
rect 33416 24948 33468 24954
rect 33416 24890 33468 24896
rect 33336 24806 33456 24834
rect 32956 23860 33008 23866
rect 32956 23802 33008 23808
rect 33048 23724 33100 23730
rect 33048 23666 33100 23672
rect 33324 23724 33376 23730
rect 33324 23666 33376 23672
rect 32864 21412 32916 21418
rect 32864 21354 32916 21360
rect 32876 20942 32904 21354
rect 32864 20936 32916 20942
rect 32864 20878 32916 20884
rect 32772 20596 32824 20602
rect 32772 20538 32824 20544
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 32508 19990 32536 20402
rect 32496 19984 32548 19990
rect 32496 19926 32548 19932
rect 32496 19712 32548 19718
rect 32496 19654 32548 19660
rect 32508 19378 32536 19654
rect 32220 19372 32272 19378
rect 32220 19314 32272 19320
rect 32496 19372 32548 19378
rect 32496 19314 32548 19320
rect 32232 18766 32260 19314
rect 32588 18964 32640 18970
rect 32588 18906 32640 18912
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32232 17610 32260 18702
rect 32496 18692 32548 18698
rect 32496 18634 32548 18640
rect 32508 18290 32536 18634
rect 32600 18426 32628 18906
rect 32588 18420 32640 18426
rect 32588 18362 32640 18368
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 32508 17610 32536 18226
rect 32680 18216 32732 18222
rect 32680 18158 32732 18164
rect 32588 18080 32640 18086
rect 32588 18022 32640 18028
rect 32220 17604 32272 17610
rect 32220 17546 32272 17552
rect 32496 17604 32548 17610
rect 32496 17546 32548 17552
rect 32508 17134 32536 17546
rect 32600 17270 32628 18022
rect 32588 17264 32640 17270
rect 32588 17206 32640 17212
rect 32496 17128 32548 17134
rect 32496 17070 32548 17076
rect 32404 17060 32456 17066
rect 32404 17002 32456 17008
rect 32416 16794 32444 17002
rect 32692 16998 32720 18158
rect 32680 16992 32732 16998
rect 32680 16934 32732 16940
rect 32404 16788 32456 16794
rect 32404 16730 32456 16736
rect 32692 16658 32720 16934
rect 32680 16652 32732 16658
rect 32680 16594 32732 16600
rect 32312 16584 32364 16590
rect 32312 16526 32364 16532
rect 32324 16250 32352 16526
rect 32496 16448 32548 16454
rect 32496 16390 32548 16396
rect 32312 16244 32364 16250
rect 32312 16186 32364 16192
rect 32508 15434 32536 16390
rect 32692 15978 32720 16594
rect 32772 16040 32824 16046
rect 32772 15982 32824 15988
rect 32680 15972 32732 15978
rect 32680 15914 32732 15920
rect 32496 15428 32548 15434
rect 32496 15370 32548 15376
rect 32784 15366 32812 15982
rect 32864 15496 32916 15502
rect 32864 15438 32916 15444
rect 32772 15360 32824 15366
rect 32772 15302 32824 15308
rect 32312 15020 32364 15026
rect 32312 14962 32364 14968
rect 32324 14618 32352 14962
rect 32312 14612 32364 14618
rect 32312 14554 32364 14560
rect 32784 14414 32812 15302
rect 32876 15094 32904 15438
rect 32864 15088 32916 15094
rect 32864 15030 32916 15036
rect 32772 14408 32824 14414
rect 32772 14350 32824 14356
rect 32876 13870 32904 15030
rect 32864 13864 32916 13870
rect 32864 13806 32916 13812
rect 32496 13796 32548 13802
rect 32496 13738 32548 13744
rect 32588 13796 32640 13802
rect 32588 13738 32640 13744
rect 32508 13190 32536 13738
rect 32600 13394 32628 13738
rect 32588 13388 32640 13394
rect 32588 13330 32640 13336
rect 32496 13184 32548 13190
rect 32496 13126 32548 13132
rect 32128 11824 32180 11830
rect 32128 11766 32180 11772
rect 31944 10804 31996 10810
rect 31944 10746 31996 10752
rect 31484 10668 31536 10674
rect 31484 10610 31536 10616
rect 31852 10464 31904 10470
rect 31852 10406 31904 10412
rect 31392 9988 31444 9994
rect 31392 9930 31444 9936
rect 31208 8628 31260 8634
rect 31208 8570 31260 8576
rect 30932 8424 30984 8430
rect 30932 8366 30984 8372
rect 30656 8356 30708 8362
rect 30656 8298 30708 8304
rect 30564 8084 30616 8090
rect 30564 8026 30616 8032
rect 30380 7880 30432 7886
rect 30380 7822 30432 7828
rect 31220 7546 31248 8570
rect 31300 8424 31352 8430
rect 31300 8366 31352 8372
rect 31312 8022 31340 8366
rect 31300 8016 31352 8022
rect 31300 7958 31352 7964
rect 31208 7540 31260 7546
rect 31208 7482 31260 7488
rect 30656 7404 30708 7410
rect 30656 7346 30708 7352
rect 29644 6928 29696 6934
rect 29644 6870 29696 6876
rect 29276 6792 29328 6798
rect 29276 6734 29328 6740
rect 29644 6792 29696 6798
rect 29644 6734 29696 6740
rect 29288 6322 29316 6734
rect 29656 6458 29684 6734
rect 30668 6730 30696 7346
rect 30656 6724 30708 6730
rect 30656 6666 30708 6672
rect 30288 6656 30340 6662
rect 30288 6598 30340 6604
rect 31116 6656 31168 6662
rect 31116 6598 31168 6604
rect 29644 6452 29696 6458
rect 29644 6394 29696 6400
rect 30300 6322 30328 6598
rect 29276 6316 29328 6322
rect 29276 6258 29328 6264
rect 30288 6316 30340 6322
rect 30288 6258 30340 6264
rect 28816 6248 28868 6254
rect 28816 6190 28868 6196
rect 30380 6112 30432 6118
rect 30380 6054 30432 6060
rect 28724 5908 28776 5914
rect 28724 5850 28776 5856
rect 30392 5846 30420 6054
rect 31128 5914 31156 6598
rect 31760 6316 31812 6322
rect 31760 6258 31812 6264
rect 31116 5908 31168 5914
rect 31116 5850 31168 5856
rect 30380 5840 30432 5846
rect 30380 5782 30432 5788
rect 30656 5568 30708 5574
rect 30656 5510 30708 5516
rect 28632 5364 28684 5370
rect 28632 5306 28684 5312
rect 30668 5030 30696 5510
rect 31128 5370 31156 5850
rect 31772 5778 31800 6258
rect 31760 5772 31812 5778
rect 31760 5714 31812 5720
rect 31116 5364 31168 5370
rect 31116 5306 31168 5312
rect 30656 5024 30708 5030
rect 30656 4966 30708 4972
rect 27988 4616 28040 4622
rect 27988 4558 28040 4564
rect 29920 4616 29972 4622
rect 29920 4558 29972 4564
rect 26424 4004 26476 4010
rect 26424 3946 26476 3952
rect 25780 3732 25832 3738
rect 25780 3674 25832 3680
rect 26436 3602 26464 3946
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 29552 3936 29604 3942
rect 29552 3878 29604 3884
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 24400 3596 24452 3602
rect 24400 3538 24452 3544
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23940 3528 23992 3534
rect 23940 3470 23992 3476
rect 26056 3528 26108 3534
rect 26056 3470 26108 3476
rect 27436 3528 27488 3534
rect 27436 3470 27488 3476
rect 23296 2848 23348 2854
rect 23296 2790 23348 2796
rect 23308 800 23336 2790
rect 23584 800 23612 3470
rect 24400 3460 24452 3466
rect 24400 3402 24452 3408
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23860 800 23888 2926
rect 24124 2576 24176 2582
rect 24124 2518 24176 2524
rect 24136 800 24164 2518
rect 24412 800 24440 3402
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 24952 2916 25004 2922
rect 24952 2858 25004 2864
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 24688 800 24716 2450
rect 24964 800 24992 2858
rect 25504 2848 25556 2854
rect 25504 2790 25556 2796
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25240 800 25268 2382
rect 25516 800 25544 2790
rect 25792 800 25820 2926
rect 26068 800 26096 3470
rect 26332 2848 26384 2854
rect 26332 2790 26384 2796
rect 26884 2848 26936 2854
rect 26884 2790 26936 2796
rect 26344 800 26372 2790
rect 26608 2372 26660 2378
rect 26608 2314 26660 2320
rect 26620 800 26648 2314
rect 26896 800 26924 2790
rect 27160 2576 27212 2582
rect 27160 2518 27212 2524
rect 27172 800 27200 2518
rect 27448 800 27476 3470
rect 27724 800 27752 3878
rect 28264 3528 28316 3534
rect 28264 3470 28316 3476
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 27988 2508 28040 2514
rect 27988 2450 28040 2456
rect 28000 800 28028 2450
rect 28276 800 28304 3470
rect 28540 2916 28592 2922
rect 28540 2858 28592 2864
rect 28552 800 28580 2858
rect 28828 800 28856 3470
rect 29012 1986 29040 3878
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 29104 3058 29132 3538
rect 29460 3528 29512 3534
rect 29460 3470 29512 3476
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 29368 2984 29420 2990
rect 29368 2926 29420 2932
rect 29012 1958 29132 1986
rect 29104 800 29132 1958
rect 29380 800 29408 2926
rect 29472 1850 29500 3470
rect 29564 3194 29592 3878
rect 29552 3188 29604 3194
rect 29552 3130 29604 3136
rect 29656 3126 29684 3878
rect 29644 3120 29696 3126
rect 29644 3062 29696 3068
rect 29472 1822 29684 1850
rect 29656 800 29684 1822
rect 29932 800 29960 4558
rect 30472 2848 30524 2854
rect 30472 2790 30524 2796
rect 30196 2576 30248 2582
rect 30196 2518 30248 2524
rect 30208 800 30236 2518
rect 30484 800 30512 2790
rect 30668 2378 30696 4966
rect 31864 4808 31892 10406
rect 31956 8634 31984 10746
rect 32600 10674 32628 13330
rect 32876 12170 32904 13806
rect 33060 13802 33088 23666
rect 33232 23520 33284 23526
rect 33232 23462 33284 23468
rect 33244 22574 33272 23462
rect 33336 23254 33364 23666
rect 33324 23248 33376 23254
rect 33324 23190 33376 23196
rect 33428 22642 33456 24806
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33232 22568 33284 22574
rect 33232 22510 33284 22516
rect 33520 21010 33548 25774
rect 33612 23798 33640 27814
rect 34612 27668 34664 27674
rect 34612 27610 34664 27616
rect 34520 26988 34572 26994
rect 34520 26930 34572 26936
rect 34428 26920 34480 26926
rect 34428 26862 34480 26868
rect 34440 25922 34468 26862
rect 34532 26042 34560 26930
rect 34520 26036 34572 26042
rect 34520 25978 34572 25984
rect 34624 25974 34652 27610
rect 34716 26382 34744 29038
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28416 34848 28422
rect 34796 28358 34848 28364
rect 34808 27674 34836 28358
rect 35360 28218 35388 29174
rect 35544 29170 35572 32302
rect 35716 31748 35768 31754
rect 35716 31690 35768 31696
rect 35728 31482 35756 31690
rect 35820 31686 35848 32370
rect 35900 32224 35952 32230
rect 35900 32166 35952 32172
rect 35808 31680 35860 31686
rect 35808 31622 35860 31628
rect 35716 31476 35768 31482
rect 35716 31418 35768 31424
rect 35820 30666 35848 31622
rect 35912 31346 35940 32166
rect 36556 32026 36584 32370
rect 37648 32292 37700 32298
rect 37648 32234 37700 32240
rect 37280 32224 37332 32230
rect 37280 32166 37332 32172
rect 37464 32224 37516 32230
rect 37464 32166 37516 32172
rect 36544 32020 36596 32026
rect 36544 31962 36596 31968
rect 36452 31952 36504 31958
rect 36452 31894 36504 31900
rect 36464 31754 36492 31894
rect 37292 31822 37320 32166
rect 37476 31822 37504 32166
rect 37660 31890 37688 32234
rect 38200 31952 38252 31958
rect 38200 31894 38252 31900
rect 37648 31884 37700 31890
rect 37648 31826 37700 31832
rect 37280 31816 37332 31822
rect 37280 31758 37332 31764
rect 37464 31816 37516 31822
rect 37464 31758 37516 31764
rect 38212 31754 38240 31894
rect 38304 31890 38332 32846
rect 38672 32570 38700 32914
rect 38752 32768 38804 32774
rect 38752 32710 38804 32716
rect 38660 32564 38712 32570
rect 38660 32506 38712 32512
rect 38764 32450 38792 32710
rect 38672 32422 38792 32450
rect 38672 32026 38700 32422
rect 40500 32360 40552 32366
rect 40500 32302 40552 32308
rect 40040 32224 40092 32230
rect 40040 32166 40092 32172
rect 38660 32020 38712 32026
rect 38660 31962 38712 31968
rect 38292 31884 38344 31890
rect 38292 31826 38344 31832
rect 38568 31816 38620 31822
rect 38568 31758 38620 31764
rect 36452 31748 36504 31754
rect 38212 31726 38332 31754
rect 36452 31690 36504 31696
rect 35900 31340 35952 31346
rect 35900 31282 35952 31288
rect 35992 31272 36044 31278
rect 35992 31214 36044 31220
rect 35808 30660 35860 30666
rect 35808 30602 35860 30608
rect 36004 29714 36032 31214
rect 36464 30938 36492 31690
rect 37004 31340 37056 31346
rect 37004 31282 37056 31288
rect 37016 30938 37044 31282
rect 37464 31136 37516 31142
rect 37464 31078 37516 31084
rect 36452 30932 36504 30938
rect 36452 30874 36504 30880
rect 37004 30932 37056 30938
rect 37004 30874 37056 30880
rect 37476 30802 37504 31078
rect 37464 30796 37516 30802
rect 37464 30738 37516 30744
rect 37280 30728 37332 30734
rect 37200 30676 37280 30682
rect 37200 30670 37332 30676
rect 37200 30654 37320 30670
rect 36360 30048 36412 30054
rect 36360 29990 36412 29996
rect 35992 29708 36044 29714
rect 35992 29650 36044 29656
rect 35900 29640 35952 29646
rect 35900 29582 35952 29588
rect 35532 29164 35584 29170
rect 35532 29106 35584 29112
rect 35348 28212 35400 28218
rect 35348 28154 35400 28160
rect 35544 28014 35572 29106
rect 35624 28416 35676 28422
rect 35624 28358 35676 28364
rect 35636 28082 35664 28358
rect 35912 28218 35940 29582
rect 36004 28626 36032 29650
rect 36176 29028 36228 29034
rect 36176 28970 36228 28976
rect 35992 28620 36044 28626
rect 35992 28562 36044 28568
rect 35900 28212 35952 28218
rect 35900 28154 35952 28160
rect 35624 28076 35676 28082
rect 35624 28018 35676 28024
rect 35532 28008 35584 28014
rect 35532 27950 35584 27956
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34796 27668 34848 27674
rect 34796 27610 34848 27616
rect 35544 27418 35572 27950
rect 35452 27390 35572 27418
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 34808 26382 34836 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34704 26376 34756 26382
rect 34704 26318 34756 26324
rect 34796 26376 34848 26382
rect 34796 26318 34848 26324
rect 34612 25968 34664 25974
rect 34440 25894 34560 25922
rect 34612 25910 34664 25916
rect 34532 25378 34560 25894
rect 34532 25350 34652 25378
rect 34520 25220 34572 25226
rect 34520 25162 34572 25168
rect 34532 24818 34560 25162
rect 34520 24812 34572 24818
rect 34520 24754 34572 24760
rect 34624 24750 34652 25350
rect 34612 24744 34664 24750
rect 34612 24686 34664 24692
rect 34624 24342 34652 24686
rect 34520 24336 34572 24342
rect 34520 24278 34572 24284
rect 34612 24336 34664 24342
rect 34612 24278 34664 24284
rect 34532 24070 34560 24278
rect 34520 24064 34572 24070
rect 34520 24006 34572 24012
rect 33600 23792 33652 23798
rect 33600 23734 33652 23740
rect 33692 23520 33744 23526
rect 33692 23462 33744 23468
rect 33704 22234 33732 23462
rect 34520 23112 34572 23118
rect 34520 23054 34572 23060
rect 33692 22228 33744 22234
rect 33692 22170 33744 22176
rect 33508 21004 33560 21010
rect 33508 20946 33560 20952
rect 33520 20398 33548 20946
rect 33600 20528 33652 20534
rect 33600 20470 33652 20476
rect 33508 20392 33560 20398
rect 33508 20334 33560 20340
rect 33324 19848 33376 19854
rect 33324 19790 33376 19796
rect 33336 18970 33364 19790
rect 33520 19446 33548 20334
rect 33612 19514 33640 20470
rect 33784 20460 33836 20466
rect 33784 20402 33836 20408
rect 33796 20058 33824 20402
rect 33784 20052 33836 20058
rect 33784 19994 33836 20000
rect 33600 19508 33652 19514
rect 33600 19450 33652 19456
rect 33508 19440 33560 19446
rect 33508 19382 33560 19388
rect 33324 18964 33376 18970
rect 33324 18906 33376 18912
rect 33612 18834 33640 19450
rect 33600 18828 33652 18834
rect 33600 18770 33652 18776
rect 33876 18828 33928 18834
rect 33876 18770 33928 18776
rect 33888 18426 33916 18770
rect 34532 18630 34560 23054
rect 34624 22094 34652 24278
rect 34716 24274 34744 26318
rect 35452 25838 35480 27390
rect 35532 27328 35584 27334
rect 35532 27270 35584 27276
rect 35440 25832 35492 25838
rect 35360 25780 35440 25786
rect 35360 25774 35492 25780
rect 35360 25758 35480 25774
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34704 24268 34756 24274
rect 34704 24210 34756 24216
rect 35360 23866 35388 25758
rect 35440 24744 35492 24750
rect 35440 24686 35492 24692
rect 35452 24410 35480 24686
rect 35440 24404 35492 24410
rect 35440 24346 35492 24352
rect 35348 23860 35400 23866
rect 35348 23802 35400 23808
rect 35348 23724 35400 23730
rect 35348 23666 35400 23672
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34704 22500 34756 22506
rect 34704 22442 34756 22448
rect 34716 22234 34744 22442
rect 34796 22432 34848 22438
rect 34796 22374 34848 22380
rect 34704 22228 34756 22234
rect 34704 22170 34756 22176
rect 34624 22066 34744 22094
rect 34612 21344 34664 21350
rect 34612 21286 34664 21292
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 33876 18420 33928 18426
rect 33876 18362 33928 18368
rect 33508 18216 33560 18222
rect 33508 18158 33560 18164
rect 33520 17882 33548 18158
rect 33508 17876 33560 17882
rect 33508 17818 33560 17824
rect 33520 17105 33548 17818
rect 33784 17604 33836 17610
rect 33784 17546 33836 17552
rect 33506 17096 33562 17105
rect 33506 17031 33562 17040
rect 33796 16590 33824 17546
rect 33784 16584 33836 16590
rect 33784 16526 33836 16532
rect 33508 16176 33560 16182
rect 33508 16118 33560 16124
rect 33232 15020 33284 15026
rect 33232 14962 33284 14968
rect 33140 14408 33192 14414
rect 33140 14350 33192 14356
rect 33048 13796 33100 13802
rect 33048 13738 33100 13744
rect 33152 13530 33180 14350
rect 33140 13524 33192 13530
rect 33140 13466 33192 13472
rect 33244 13462 33272 14962
rect 33416 14272 33468 14278
rect 33416 14214 33468 14220
rect 33428 13938 33456 14214
rect 33416 13932 33468 13938
rect 33416 13874 33468 13880
rect 33232 13456 33284 13462
rect 33232 13398 33284 13404
rect 33416 13320 33468 13326
rect 33416 13262 33468 13268
rect 33324 12912 33376 12918
rect 33324 12854 33376 12860
rect 33140 12640 33192 12646
rect 33140 12582 33192 12588
rect 32864 12164 32916 12170
rect 32864 12106 32916 12112
rect 33048 12164 33100 12170
rect 33048 12106 33100 12112
rect 33060 11694 33088 12106
rect 33152 11762 33180 12582
rect 33140 11756 33192 11762
rect 33140 11698 33192 11704
rect 33048 11688 33100 11694
rect 33048 11630 33100 11636
rect 33060 11150 33088 11630
rect 33140 11620 33192 11626
rect 33140 11562 33192 11568
rect 33152 11286 33180 11562
rect 33140 11280 33192 11286
rect 33140 11222 33192 11228
rect 33048 11144 33100 11150
rect 33048 11086 33100 11092
rect 32312 10668 32364 10674
rect 32312 10610 32364 10616
rect 32588 10668 32640 10674
rect 32588 10610 32640 10616
rect 32128 10124 32180 10130
rect 32128 10066 32180 10072
rect 32140 9654 32168 10066
rect 32324 9722 32352 10610
rect 32600 10130 32628 10610
rect 32588 10124 32640 10130
rect 32588 10066 32640 10072
rect 32312 9716 32364 9722
rect 32312 9658 32364 9664
rect 32128 9648 32180 9654
rect 32128 9590 32180 9596
rect 32140 9178 32168 9590
rect 32588 9512 32640 9518
rect 32588 9454 32640 9460
rect 32128 9172 32180 9178
rect 32128 9114 32180 9120
rect 32312 8900 32364 8906
rect 32312 8842 32364 8848
rect 31944 8628 31996 8634
rect 31944 8570 31996 8576
rect 32324 8498 32352 8842
rect 32312 8492 32364 8498
rect 32312 8434 32364 8440
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 32508 7834 32536 8434
rect 32600 7954 32628 9454
rect 33060 8974 33088 11086
rect 33336 9586 33364 12854
rect 33428 12850 33456 13262
rect 33416 12844 33468 12850
rect 33416 12786 33468 12792
rect 33520 10810 33548 16118
rect 33796 12918 33824 16526
rect 33888 13394 33916 18362
rect 34520 18284 34572 18290
rect 34520 18226 34572 18232
rect 34532 17338 34560 18226
rect 34520 17332 34572 17338
rect 34520 17274 34572 17280
rect 34520 16720 34572 16726
rect 34520 16662 34572 16668
rect 33968 16516 34020 16522
rect 33968 16458 34020 16464
rect 33980 16250 34008 16458
rect 34152 16448 34204 16454
rect 34152 16390 34204 16396
rect 34428 16448 34480 16454
rect 34428 16390 34480 16396
rect 33968 16244 34020 16250
rect 33968 16186 34020 16192
rect 34164 16114 34192 16390
rect 34440 16182 34468 16390
rect 34428 16176 34480 16182
rect 34428 16118 34480 16124
rect 34152 16108 34204 16114
rect 34152 16050 34204 16056
rect 34428 15904 34480 15910
rect 34428 15846 34480 15852
rect 34440 15094 34468 15846
rect 34532 15162 34560 16662
rect 34624 16046 34652 21286
rect 34716 18222 34744 22066
rect 34808 22030 34836 22374
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34888 22228 34940 22234
rect 34888 22170 34940 22176
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34900 21350 34928 22170
rect 35256 21480 35308 21486
rect 35256 21422 35308 21428
rect 34888 21344 34940 21350
rect 34888 21286 34940 21292
rect 35268 21298 35296 21422
rect 35360 21298 35388 23666
rect 35440 23316 35492 23322
rect 35440 23258 35492 23264
rect 35452 22778 35480 23258
rect 35544 23118 35572 27270
rect 35624 26988 35676 26994
rect 35624 26930 35676 26936
rect 35636 26790 35664 26930
rect 35624 26784 35676 26790
rect 35624 26726 35676 26732
rect 35532 23112 35584 23118
rect 35532 23054 35584 23060
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35440 22772 35492 22778
rect 35440 22714 35492 22720
rect 35440 21956 35492 21962
rect 35440 21898 35492 21904
rect 35452 21486 35480 21898
rect 35544 21622 35572 22918
rect 35532 21616 35584 21622
rect 35532 21558 35584 21564
rect 35440 21480 35492 21486
rect 35440 21422 35492 21428
rect 35268 21270 35388 21298
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34704 18216 34756 18222
rect 34704 18158 34756 18164
rect 34704 18080 34756 18086
rect 34704 18022 34756 18028
rect 34716 17678 34744 18022
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35072 17740 35124 17746
rect 35072 17682 35124 17688
rect 34704 17672 34756 17678
rect 34704 17614 34756 17620
rect 34796 17536 34848 17542
rect 34796 17478 34848 17484
rect 34808 17134 34836 17478
rect 35084 17338 35112 17682
rect 35072 17332 35124 17338
rect 35072 17274 35124 17280
rect 35360 17270 35388 21270
rect 35452 21078 35480 21422
rect 35440 21072 35492 21078
rect 35440 21014 35492 21020
rect 35440 19916 35492 19922
rect 35440 19858 35492 19864
rect 35452 19174 35480 19858
rect 35544 19786 35572 21558
rect 35636 20806 35664 26726
rect 35900 25152 35952 25158
rect 35900 25094 35952 25100
rect 35716 24812 35768 24818
rect 35716 24754 35768 24760
rect 35728 22982 35756 24754
rect 35808 24336 35860 24342
rect 35808 24278 35860 24284
rect 35820 23730 35848 24278
rect 35912 24206 35940 25094
rect 36004 24274 36032 28562
rect 36188 28558 36216 28970
rect 36372 28558 36400 29990
rect 37200 28762 37228 30654
rect 37280 30252 37332 30258
rect 37280 30194 37332 30200
rect 37292 29306 37320 30194
rect 37648 29844 37700 29850
rect 37648 29786 37700 29792
rect 37372 29504 37424 29510
rect 37372 29446 37424 29452
rect 37280 29300 37332 29306
rect 37280 29242 37332 29248
rect 36452 28756 36504 28762
rect 36452 28698 36504 28704
rect 37188 28756 37240 28762
rect 37188 28698 37240 28704
rect 36176 28552 36228 28558
rect 36176 28494 36228 28500
rect 36360 28552 36412 28558
rect 36360 28494 36412 28500
rect 36084 28484 36136 28490
rect 36084 28426 36136 28432
rect 36096 28082 36124 28426
rect 36084 28076 36136 28082
rect 36084 28018 36136 28024
rect 36096 27674 36124 28018
rect 36084 27668 36136 27674
rect 36084 27610 36136 27616
rect 36464 27606 36492 28698
rect 37384 28218 37412 29446
rect 37660 29306 37688 29786
rect 37648 29300 37700 29306
rect 37648 29242 37700 29248
rect 37464 29096 37516 29102
rect 37464 29038 37516 29044
rect 37476 28626 37504 29038
rect 37830 28656 37886 28665
rect 37464 28620 37516 28626
rect 37830 28591 37886 28600
rect 37464 28562 37516 28568
rect 37476 28422 37504 28562
rect 37464 28416 37516 28422
rect 37464 28358 37516 28364
rect 37372 28212 37424 28218
rect 37372 28154 37424 28160
rect 37384 28014 37412 28154
rect 37372 28008 37424 28014
rect 37372 27950 37424 27956
rect 36452 27600 36504 27606
rect 36452 27542 36504 27548
rect 36084 26920 36136 26926
rect 36084 26862 36136 26868
rect 36096 26246 36124 26862
rect 36464 26586 36492 27542
rect 37476 27470 37504 28358
rect 37844 28218 37872 28591
rect 38108 28552 38160 28558
rect 38108 28494 38160 28500
rect 37832 28212 37884 28218
rect 37832 28154 37884 28160
rect 37924 27940 37976 27946
rect 37924 27882 37976 27888
rect 37936 27674 37964 27882
rect 37924 27668 37976 27674
rect 37844 27628 37924 27656
rect 37464 27464 37516 27470
rect 37464 27406 37516 27412
rect 36728 27328 36780 27334
rect 36728 27270 36780 27276
rect 36740 26858 36768 27270
rect 36728 26852 36780 26858
rect 36728 26794 36780 26800
rect 36452 26580 36504 26586
rect 36452 26522 36504 26528
rect 36452 26308 36504 26314
rect 36452 26250 36504 26256
rect 36084 26240 36136 26246
rect 36084 26182 36136 26188
rect 36096 25770 36124 26182
rect 36084 25764 36136 25770
rect 36084 25706 36136 25712
rect 36464 25702 36492 26250
rect 37464 26240 37516 26246
rect 37464 26182 37516 26188
rect 37476 25838 37504 26182
rect 37464 25832 37516 25838
rect 37464 25774 37516 25780
rect 36452 25696 36504 25702
rect 36452 25638 36504 25644
rect 36360 24608 36412 24614
rect 36360 24550 36412 24556
rect 35992 24268 36044 24274
rect 35992 24210 36044 24216
rect 35900 24200 35952 24206
rect 35900 24142 35952 24148
rect 36372 24138 36400 24550
rect 36360 24132 36412 24138
rect 36360 24074 36412 24080
rect 35808 23724 35860 23730
rect 35808 23666 35860 23672
rect 35716 22976 35768 22982
rect 35716 22918 35768 22924
rect 35820 22438 35848 23666
rect 35808 22432 35860 22438
rect 35808 22374 35860 22380
rect 35716 21548 35768 21554
rect 35716 21490 35768 21496
rect 35728 21146 35756 21490
rect 36268 21344 36320 21350
rect 36268 21286 36320 21292
rect 35716 21140 35768 21146
rect 35716 21082 35768 21088
rect 35624 20800 35676 20806
rect 35624 20742 35676 20748
rect 36280 20466 36308 21286
rect 36268 20460 36320 20466
rect 36268 20402 36320 20408
rect 35808 20256 35860 20262
rect 35808 20198 35860 20204
rect 35820 19854 35848 20198
rect 35808 19848 35860 19854
rect 35808 19790 35860 19796
rect 35532 19780 35584 19786
rect 35532 19722 35584 19728
rect 36464 19174 36492 25638
rect 37476 25294 37504 25774
rect 37740 25764 37792 25770
rect 37740 25706 37792 25712
rect 37752 25498 37780 25706
rect 37740 25492 37792 25498
rect 37740 25434 37792 25440
rect 37464 25288 37516 25294
rect 37464 25230 37516 25236
rect 37648 24404 37700 24410
rect 37648 24346 37700 24352
rect 37660 23730 37688 24346
rect 37648 23724 37700 23730
rect 37648 23666 37700 23672
rect 37844 23322 37872 27628
rect 37924 27610 37976 27616
rect 37924 26376 37976 26382
rect 37924 26318 37976 26324
rect 37936 25498 37964 26318
rect 38016 26308 38068 26314
rect 38016 26250 38068 26256
rect 37924 25492 37976 25498
rect 37924 25434 37976 25440
rect 37832 23316 37884 23322
rect 37832 23258 37884 23264
rect 37844 23186 37872 23258
rect 37832 23180 37884 23186
rect 37832 23122 37884 23128
rect 37556 22976 37608 22982
rect 37556 22918 37608 22924
rect 36728 22024 36780 22030
rect 36728 21966 36780 21972
rect 36740 21554 36768 21966
rect 37372 21888 37424 21894
rect 37372 21830 37424 21836
rect 36728 21548 36780 21554
rect 36728 21490 36780 21496
rect 37384 21486 37412 21830
rect 37372 21480 37424 21486
rect 37372 21422 37424 21428
rect 37568 21418 37596 22918
rect 38028 22094 38056 26250
rect 38120 24070 38148 28494
rect 38200 26920 38252 26926
rect 38200 26862 38252 26868
rect 38212 26586 38240 26862
rect 38200 26580 38252 26586
rect 38200 26522 38252 26528
rect 38200 26308 38252 26314
rect 38200 26250 38252 26256
rect 38212 26042 38240 26250
rect 38200 26036 38252 26042
rect 38200 25978 38252 25984
rect 38108 24064 38160 24070
rect 38108 24006 38160 24012
rect 38108 23316 38160 23322
rect 38108 23258 38160 23264
rect 37936 22066 38056 22094
rect 37832 22024 37884 22030
rect 37832 21966 37884 21972
rect 37740 21888 37792 21894
rect 37740 21830 37792 21836
rect 37556 21412 37608 21418
rect 37556 21354 37608 21360
rect 37280 20868 37332 20874
rect 37280 20810 37332 20816
rect 37292 20602 37320 20810
rect 37280 20596 37332 20602
rect 37280 20538 37332 20544
rect 37568 20534 37596 21354
rect 37752 21350 37780 21830
rect 37740 21344 37792 21350
rect 37740 21286 37792 21292
rect 37752 20942 37780 21286
rect 37844 21010 37872 21966
rect 37832 21004 37884 21010
rect 37832 20946 37884 20952
rect 37740 20936 37792 20942
rect 37740 20878 37792 20884
rect 37556 20528 37608 20534
rect 37556 20470 37608 20476
rect 37936 20058 37964 22066
rect 38120 21554 38148 23258
rect 38304 22030 38332 31726
rect 38580 31142 38608 31758
rect 38568 31136 38620 31142
rect 38568 31078 38620 31084
rect 38672 29510 38700 31962
rect 40052 31822 40080 32166
rect 40040 31816 40092 31822
rect 40040 31758 40092 31764
rect 40408 31680 40460 31686
rect 40408 31622 40460 31628
rect 40420 30258 40448 31622
rect 40408 30252 40460 30258
rect 40408 30194 40460 30200
rect 40132 30048 40184 30054
rect 40132 29990 40184 29996
rect 38660 29504 38712 29510
rect 38660 29446 38712 29452
rect 39672 29164 39724 29170
rect 39672 29106 39724 29112
rect 38752 29096 38804 29102
rect 38752 29038 38804 29044
rect 38660 27328 38712 27334
rect 38660 27270 38712 27276
rect 38672 25684 38700 27270
rect 38764 27062 38792 29038
rect 39304 28008 39356 28014
rect 39304 27950 39356 27956
rect 39212 27532 39264 27538
rect 39212 27474 39264 27480
rect 38752 27056 38804 27062
rect 38752 26998 38804 27004
rect 38844 26988 38896 26994
rect 38844 26930 38896 26936
rect 38856 26382 38884 26930
rect 39224 26790 39252 27474
rect 39316 27470 39344 27950
rect 39304 27464 39356 27470
rect 39304 27406 39356 27412
rect 39212 26784 39264 26790
rect 39212 26726 39264 26732
rect 39224 26382 39252 26726
rect 38844 26376 38896 26382
rect 38844 26318 38896 26324
rect 39212 26376 39264 26382
rect 39212 26318 39264 26324
rect 38752 25696 38804 25702
rect 38672 25656 38752 25684
rect 38752 25638 38804 25644
rect 38764 24682 38792 25638
rect 38752 24676 38804 24682
rect 38752 24618 38804 24624
rect 38568 24200 38620 24206
rect 38568 24142 38620 24148
rect 38580 23186 38608 24142
rect 38660 23656 38712 23662
rect 38660 23598 38712 23604
rect 38672 23322 38700 23598
rect 38660 23316 38712 23322
rect 38660 23258 38712 23264
rect 38568 23180 38620 23186
rect 38568 23122 38620 23128
rect 38292 22024 38344 22030
rect 38292 21966 38344 21972
rect 38108 21548 38160 21554
rect 38108 21490 38160 21496
rect 38016 20800 38068 20806
rect 38016 20742 38068 20748
rect 37924 20052 37976 20058
rect 37924 19994 37976 20000
rect 38028 19922 38056 20742
rect 38016 19916 38068 19922
rect 38016 19858 38068 19864
rect 38856 19378 38884 26318
rect 39028 23180 39080 23186
rect 39028 23122 39080 23128
rect 39040 22642 39068 23122
rect 39028 22636 39080 22642
rect 39028 22578 39080 22584
rect 38844 19372 38896 19378
rect 38844 19314 38896 19320
rect 39224 19310 39252 26318
rect 39316 25906 39344 27406
rect 39580 27328 39632 27334
rect 39580 27270 39632 27276
rect 39592 26994 39620 27270
rect 39580 26988 39632 26994
rect 39580 26930 39632 26936
rect 39684 26586 39712 29106
rect 39764 27396 39816 27402
rect 39764 27338 39816 27344
rect 39776 26994 39804 27338
rect 39764 26988 39816 26994
rect 39764 26930 39816 26936
rect 39856 26920 39908 26926
rect 39856 26862 39908 26868
rect 39672 26580 39724 26586
rect 39672 26522 39724 26528
rect 39868 26042 39896 26862
rect 40040 26852 40092 26858
rect 40040 26794 40092 26800
rect 40052 26382 40080 26794
rect 40040 26376 40092 26382
rect 40040 26318 40092 26324
rect 39856 26036 39908 26042
rect 39856 25978 39908 25984
rect 39304 25900 39356 25906
rect 39304 25842 39356 25848
rect 39316 24818 39344 25842
rect 39304 24812 39356 24818
rect 39304 24754 39356 24760
rect 39764 24268 39816 24274
rect 39764 24210 39816 24216
rect 39776 23662 39804 24210
rect 39764 23656 39816 23662
rect 39764 23598 39816 23604
rect 39776 22574 39804 23598
rect 39856 22976 39908 22982
rect 39856 22918 39908 22924
rect 39948 22976 40000 22982
rect 39948 22918 40000 22924
rect 39764 22568 39816 22574
rect 39764 22510 39816 22516
rect 39868 22030 39896 22918
rect 39960 22642 39988 22918
rect 39948 22636 40000 22642
rect 39948 22578 40000 22584
rect 40040 22636 40092 22642
rect 40040 22578 40092 22584
rect 40052 22234 40080 22578
rect 40040 22228 40092 22234
rect 40040 22170 40092 22176
rect 39856 22024 39908 22030
rect 39856 21966 39908 21972
rect 39856 21344 39908 21350
rect 39856 21286 39908 21292
rect 39868 20942 39896 21286
rect 40144 21146 40172 29990
rect 40316 29096 40368 29102
rect 40316 29038 40368 29044
rect 40328 27606 40356 29038
rect 40316 27600 40368 27606
rect 40316 27542 40368 27548
rect 40224 27328 40276 27334
rect 40224 27270 40276 27276
rect 40236 27130 40264 27270
rect 40224 27124 40276 27130
rect 40224 27066 40276 27072
rect 40236 25906 40264 27066
rect 40328 26382 40356 27542
rect 40512 27130 40540 32302
rect 41144 32224 41196 32230
rect 41144 32166 41196 32172
rect 41156 31890 41184 32166
rect 41144 31884 41196 31890
rect 41144 31826 41196 31832
rect 41236 31816 41288 31822
rect 41236 31758 41288 31764
rect 41880 31816 41932 31822
rect 41880 31758 41932 31764
rect 40868 31680 40920 31686
rect 40868 31622 40920 31628
rect 40684 30252 40736 30258
rect 40684 30194 40736 30200
rect 40776 30252 40828 30258
rect 40776 30194 40828 30200
rect 40592 30184 40644 30190
rect 40592 30126 40644 30132
rect 40604 29850 40632 30126
rect 40592 29844 40644 29850
rect 40592 29786 40644 29792
rect 40696 29306 40724 30194
rect 40788 29782 40816 30194
rect 40880 30054 40908 31622
rect 41248 31482 41276 31758
rect 41892 31482 41920 31758
rect 42064 31680 42116 31686
rect 42064 31622 42116 31628
rect 41236 31476 41288 31482
rect 41236 31418 41288 31424
rect 41880 31476 41932 31482
rect 41880 31418 41932 31424
rect 41248 30938 41276 31418
rect 41512 31204 41564 31210
rect 41512 31146 41564 31152
rect 41236 30932 41288 30938
rect 41236 30874 41288 30880
rect 41524 30054 41552 31146
rect 42076 30734 42104 31622
rect 42432 31340 42484 31346
rect 42432 31282 42484 31288
rect 42064 30728 42116 30734
rect 42064 30670 42116 30676
rect 42444 30394 42472 31282
rect 43536 31136 43588 31142
rect 43536 31078 43588 31084
rect 42432 30388 42484 30394
rect 42432 30330 42484 30336
rect 43548 30326 43576 31078
rect 43812 30728 43864 30734
rect 43812 30670 43864 30676
rect 43536 30320 43588 30326
rect 43536 30262 43588 30268
rect 43824 30258 43852 30670
rect 43812 30252 43864 30258
rect 43812 30194 43864 30200
rect 41604 30116 41656 30122
rect 41604 30058 41656 30064
rect 40868 30048 40920 30054
rect 40868 29990 40920 29996
rect 41512 30048 41564 30054
rect 41512 29990 41564 29996
rect 40776 29776 40828 29782
rect 40776 29718 40828 29724
rect 41052 29708 41104 29714
rect 41052 29650 41104 29656
rect 40960 29504 41012 29510
rect 40960 29446 41012 29452
rect 40684 29300 40736 29306
rect 40684 29242 40736 29248
rect 40684 29164 40736 29170
rect 40684 29106 40736 29112
rect 40696 28694 40724 29106
rect 40684 28688 40736 28694
rect 40684 28630 40736 28636
rect 40500 27124 40552 27130
rect 40500 27066 40552 27072
rect 40408 26512 40460 26518
rect 40408 26454 40460 26460
rect 40592 26512 40644 26518
rect 40592 26454 40644 26460
rect 40316 26376 40368 26382
rect 40316 26318 40368 26324
rect 40224 25900 40276 25906
rect 40224 25842 40276 25848
rect 40420 24698 40448 26454
rect 40604 24818 40632 26454
rect 40696 26382 40724 28630
rect 40776 27056 40828 27062
rect 40776 26998 40828 27004
rect 40788 26586 40816 26998
rect 40776 26580 40828 26586
rect 40776 26522 40828 26528
rect 40684 26376 40736 26382
rect 40684 26318 40736 26324
rect 40788 25906 40816 26522
rect 40776 25900 40828 25906
rect 40776 25842 40828 25848
rect 40592 24812 40644 24818
rect 40592 24754 40644 24760
rect 40328 24670 40448 24698
rect 40132 21140 40184 21146
rect 40132 21082 40184 21088
rect 39948 21004 40000 21010
rect 39948 20946 40000 20952
rect 39856 20936 39908 20942
rect 39856 20878 39908 20884
rect 39304 20868 39356 20874
rect 39304 20810 39356 20816
rect 39316 20398 39344 20810
rect 39304 20392 39356 20398
rect 39304 20334 39356 20340
rect 39316 19446 39344 20334
rect 39960 19990 39988 20946
rect 40132 20936 40184 20942
rect 40132 20878 40184 20884
rect 40144 20602 40172 20878
rect 40132 20596 40184 20602
rect 40132 20538 40184 20544
rect 40328 20466 40356 24670
rect 40408 24608 40460 24614
rect 40408 24550 40460 24556
rect 40420 20466 40448 24550
rect 40500 24404 40552 24410
rect 40500 24346 40552 24352
rect 40512 24206 40540 24346
rect 40500 24200 40552 24206
rect 40500 24142 40552 24148
rect 40512 22098 40540 24142
rect 40776 24132 40828 24138
rect 40776 24074 40828 24080
rect 40788 23866 40816 24074
rect 40776 23860 40828 23866
rect 40776 23802 40828 23808
rect 40868 23860 40920 23866
rect 40868 23802 40920 23808
rect 40880 23186 40908 23802
rect 40868 23180 40920 23186
rect 40868 23122 40920 23128
rect 40776 23044 40828 23050
rect 40776 22986 40828 22992
rect 40788 22710 40816 22986
rect 40776 22704 40828 22710
rect 40776 22646 40828 22652
rect 40500 22092 40552 22098
rect 40972 22094 41000 29446
rect 41064 29306 41092 29650
rect 41052 29300 41104 29306
rect 41052 29242 41104 29248
rect 41420 27872 41472 27878
rect 41420 27814 41472 27820
rect 41432 27470 41460 27814
rect 41524 27538 41552 29990
rect 41616 29646 41644 30058
rect 41604 29640 41656 29646
rect 41604 29582 41656 29588
rect 42800 29504 42852 29510
rect 42800 29446 42852 29452
rect 42812 29102 42840 29446
rect 43352 29164 43404 29170
rect 43352 29106 43404 29112
rect 42800 29096 42852 29102
rect 42800 29038 42852 29044
rect 42812 28558 42840 29038
rect 43364 28626 43392 29106
rect 43628 29028 43680 29034
rect 43628 28970 43680 28976
rect 43444 28960 43496 28966
rect 43444 28902 43496 28908
rect 43352 28620 43404 28626
rect 43352 28562 43404 28568
rect 43456 28558 43484 28902
rect 42248 28552 42300 28558
rect 42246 28520 42248 28529
rect 42800 28552 42852 28558
rect 42300 28520 42302 28529
rect 42800 28494 42852 28500
rect 43444 28552 43496 28558
rect 43444 28494 43496 28500
rect 42246 28455 42302 28464
rect 43456 27538 43484 28494
rect 41512 27532 41564 27538
rect 41512 27474 41564 27480
rect 43444 27532 43496 27538
rect 43444 27474 43496 27480
rect 43640 27470 43668 28970
rect 43720 28076 43772 28082
rect 43824 28064 43852 30194
rect 43996 28416 44048 28422
rect 43996 28358 44048 28364
rect 44008 28150 44036 28358
rect 43996 28144 44048 28150
rect 43996 28086 44048 28092
rect 43772 28036 43852 28064
rect 43720 28018 43772 28024
rect 41420 27464 41472 27470
rect 41420 27406 41472 27412
rect 43628 27464 43680 27470
rect 43628 27406 43680 27412
rect 41328 27328 41380 27334
rect 41328 27270 41380 27276
rect 42432 27328 42484 27334
rect 42432 27270 42484 27276
rect 41052 26988 41104 26994
rect 41052 26930 41104 26936
rect 41064 26042 41092 26930
rect 41340 26518 41368 27270
rect 41328 26512 41380 26518
rect 41328 26454 41380 26460
rect 42444 26382 42472 27270
rect 43628 26988 43680 26994
rect 43732 26976 43760 28018
rect 43904 27328 43956 27334
rect 43904 27270 43956 27276
rect 43916 27062 43944 27270
rect 43904 27056 43956 27062
rect 43904 26998 43956 27004
rect 43680 26948 43760 26976
rect 43628 26930 43680 26936
rect 43640 26450 43668 26930
rect 43628 26444 43680 26450
rect 43628 26386 43680 26392
rect 41144 26376 41196 26382
rect 41144 26318 41196 26324
rect 42432 26376 42484 26382
rect 42432 26318 42484 26324
rect 41052 26036 41104 26042
rect 41052 25978 41104 25984
rect 41064 25702 41092 25978
rect 41052 25696 41104 25702
rect 41052 25638 41104 25644
rect 41156 24750 41184 26318
rect 41512 25696 41564 25702
rect 41512 25638 41564 25644
rect 41144 24744 41196 24750
rect 41144 24686 41196 24692
rect 41236 23724 41288 23730
rect 41236 23666 41288 23672
rect 41248 23322 41276 23666
rect 41236 23316 41288 23322
rect 41236 23258 41288 23264
rect 41236 22432 41288 22438
rect 41236 22374 41288 22380
rect 41248 22234 41276 22374
rect 41236 22228 41288 22234
rect 41236 22170 41288 22176
rect 40972 22066 41184 22094
rect 40500 22034 40552 22040
rect 40040 20460 40092 20466
rect 40040 20402 40092 20408
rect 40316 20460 40368 20466
rect 40316 20402 40368 20408
rect 40408 20460 40460 20466
rect 40408 20402 40460 20408
rect 40052 20058 40080 20402
rect 40040 20052 40092 20058
rect 40040 19994 40092 20000
rect 40328 19990 40356 20402
rect 39948 19984 40000 19990
rect 39948 19926 40000 19932
rect 40316 19984 40368 19990
rect 40316 19926 40368 19932
rect 40420 19854 40448 20402
rect 40408 19848 40460 19854
rect 40408 19790 40460 19796
rect 41156 19786 41184 22066
rect 41236 20868 41288 20874
rect 41236 20810 41288 20816
rect 41248 20602 41276 20810
rect 41236 20596 41288 20602
rect 41236 20538 41288 20544
rect 41420 20256 41472 20262
rect 41420 20198 41472 20204
rect 41432 20058 41460 20198
rect 41420 20052 41472 20058
rect 41420 19994 41472 20000
rect 40592 19780 40644 19786
rect 40592 19722 40644 19728
rect 40684 19780 40736 19786
rect 40684 19722 40736 19728
rect 41144 19780 41196 19786
rect 41144 19722 41196 19728
rect 39304 19440 39356 19446
rect 39304 19382 39356 19388
rect 39212 19304 39264 19310
rect 39212 19246 39264 19252
rect 35440 19168 35492 19174
rect 35440 19110 35492 19116
rect 36452 19168 36504 19174
rect 36452 19110 36504 19116
rect 36084 17672 36136 17678
rect 36084 17614 36136 17620
rect 35348 17264 35400 17270
rect 35348 17206 35400 17212
rect 34796 17128 34848 17134
rect 34796 17070 34848 17076
rect 34808 16114 34836 17070
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 36096 16658 36124 17614
rect 36464 17610 36492 19110
rect 39316 18834 39344 19382
rect 39672 19372 39724 19378
rect 39672 19314 39724 19320
rect 40132 19372 40184 19378
rect 40132 19314 40184 19320
rect 39304 18828 39356 18834
rect 39304 18770 39356 18776
rect 38016 18692 38068 18698
rect 38016 18634 38068 18640
rect 38844 18692 38896 18698
rect 38844 18634 38896 18640
rect 37924 18624 37976 18630
rect 37924 18566 37976 18572
rect 37936 18426 37964 18566
rect 38028 18426 38056 18634
rect 38856 18426 38884 18634
rect 37924 18420 37976 18426
rect 37924 18362 37976 18368
rect 38016 18420 38068 18426
rect 38016 18362 38068 18368
rect 38844 18420 38896 18426
rect 38844 18362 38896 18368
rect 37832 18216 37884 18222
rect 37832 18158 37884 18164
rect 37844 17882 37872 18158
rect 37832 17876 37884 17882
rect 37832 17818 37884 17824
rect 36452 17604 36504 17610
rect 36452 17546 36504 17552
rect 37464 17604 37516 17610
rect 37464 17546 37516 17552
rect 36464 16998 36492 17546
rect 37476 17338 37504 17546
rect 37188 17332 37240 17338
rect 37188 17274 37240 17280
rect 37464 17332 37516 17338
rect 37464 17274 37516 17280
rect 36452 16992 36504 16998
rect 36452 16934 36504 16940
rect 36464 16794 36492 16934
rect 36452 16788 36504 16794
rect 36452 16730 36504 16736
rect 36084 16652 36136 16658
rect 36084 16594 36136 16600
rect 34796 16108 34848 16114
rect 34796 16050 34848 16056
rect 34612 16040 34664 16046
rect 34612 15982 34664 15988
rect 34520 15156 34572 15162
rect 34520 15098 34572 15104
rect 34428 15088 34480 15094
rect 34428 15030 34480 15036
rect 34520 13728 34572 13734
rect 34520 13670 34572 13676
rect 33876 13388 33928 13394
rect 33876 13330 33928 13336
rect 33784 12912 33836 12918
rect 33784 12854 33836 12860
rect 33888 12782 33916 13330
rect 34532 13326 34560 13670
rect 34520 13320 34572 13326
rect 34520 13262 34572 13268
rect 33600 12776 33652 12782
rect 33600 12718 33652 12724
rect 33692 12776 33744 12782
rect 33692 12718 33744 12724
rect 33876 12776 33928 12782
rect 33876 12718 33928 12724
rect 33612 11558 33640 12718
rect 33600 11552 33652 11558
rect 33600 11494 33652 11500
rect 33600 11144 33652 11150
rect 33600 11086 33652 11092
rect 33612 10810 33640 11086
rect 33704 11082 33732 12718
rect 33968 12096 34020 12102
rect 33968 12038 34020 12044
rect 33784 11756 33836 11762
rect 33784 11698 33836 11704
rect 33796 11354 33824 11698
rect 33784 11348 33836 11354
rect 33784 11290 33836 11296
rect 33692 11076 33744 11082
rect 33692 11018 33744 11024
rect 33508 10804 33560 10810
rect 33508 10746 33560 10752
rect 33600 10804 33652 10810
rect 33600 10746 33652 10752
rect 33520 10266 33548 10746
rect 33704 10606 33732 11018
rect 33692 10600 33744 10606
rect 33692 10542 33744 10548
rect 33508 10260 33560 10266
rect 33508 10202 33560 10208
rect 33520 9926 33548 10202
rect 33980 9926 34008 12038
rect 34428 10192 34480 10198
rect 34428 10134 34480 10140
rect 33508 9920 33560 9926
rect 33508 9862 33560 9868
rect 33968 9920 34020 9926
rect 33968 9862 34020 9868
rect 33980 9722 34008 9862
rect 33968 9716 34020 9722
rect 33968 9658 34020 9664
rect 33324 9580 33376 9586
rect 33324 9522 33376 9528
rect 34440 9450 34468 10134
rect 34428 9444 34480 9450
rect 34428 9386 34480 9392
rect 34624 9178 34652 15982
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 37200 15026 37228 17274
rect 37280 17196 37332 17202
rect 37280 17138 37332 17144
rect 37292 16794 37320 17138
rect 37280 16788 37332 16794
rect 37280 16730 37332 16736
rect 37844 16658 37872 17818
rect 39316 17678 39344 18770
rect 39684 18154 39712 19314
rect 39764 19304 39816 19310
rect 39764 19246 39816 19252
rect 39672 18148 39724 18154
rect 39672 18090 39724 18096
rect 38660 17672 38712 17678
rect 38660 17614 38712 17620
rect 39304 17672 39356 17678
rect 39304 17614 39356 17620
rect 38672 17270 38700 17614
rect 38936 17536 38988 17542
rect 38936 17478 38988 17484
rect 38948 17270 38976 17478
rect 38660 17264 38712 17270
rect 38660 17206 38712 17212
rect 38936 17264 38988 17270
rect 38936 17206 38988 17212
rect 38568 16788 38620 16794
rect 38568 16730 38620 16736
rect 38580 16658 38608 16730
rect 38948 16726 38976 17206
rect 38936 16720 38988 16726
rect 38936 16662 38988 16668
rect 37832 16652 37884 16658
rect 37832 16594 37884 16600
rect 38568 16652 38620 16658
rect 38568 16594 38620 16600
rect 38108 16448 38160 16454
rect 38108 16390 38160 16396
rect 38844 16448 38896 16454
rect 38844 16390 38896 16396
rect 37188 15020 37240 15026
rect 37188 14962 37240 14968
rect 36452 14816 36504 14822
rect 36452 14758 36504 14764
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35532 14544 35584 14550
rect 35532 14486 35584 14492
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35544 12918 35572 14486
rect 36176 14340 36228 14346
rect 36176 14282 36228 14288
rect 36188 14074 36216 14282
rect 35992 14068 36044 14074
rect 35992 14010 36044 14016
rect 36176 14068 36228 14074
rect 36176 14010 36228 14016
rect 35624 14000 35676 14006
rect 35624 13942 35676 13948
rect 35532 12912 35584 12918
rect 35532 12854 35584 12860
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34704 11552 34756 11558
rect 34704 11494 34756 11500
rect 34716 10742 34744 11494
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34704 10736 34756 10742
rect 34704 10678 34756 10684
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35348 9580 35400 9586
rect 35348 9522 35400 9528
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34612 9172 34664 9178
rect 34612 9114 34664 9120
rect 33048 8968 33100 8974
rect 33048 8910 33100 8916
rect 33140 8968 33192 8974
rect 33140 8910 33192 8916
rect 33598 8936 33654 8945
rect 32680 8900 32732 8906
rect 32680 8842 32732 8848
rect 32692 8566 32720 8842
rect 33152 8820 33180 8910
rect 33598 8871 33654 8880
rect 33060 8792 33180 8820
rect 33060 8634 33088 8792
rect 33048 8628 33100 8634
rect 33048 8570 33100 8576
rect 32680 8560 32732 8566
rect 32680 8502 32732 8508
rect 33612 8430 33640 8871
rect 33600 8424 33652 8430
rect 33600 8366 33652 8372
rect 32956 8288 33008 8294
rect 32956 8230 33008 8236
rect 32588 7948 32640 7954
rect 32588 7890 32640 7896
rect 32416 7806 32536 7834
rect 32416 7750 32444 7806
rect 32404 7744 32456 7750
rect 32404 7686 32456 7692
rect 32416 7410 32444 7686
rect 32404 7404 32456 7410
rect 32404 7346 32456 7352
rect 32128 7336 32180 7342
rect 32128 7278 32180 7284
rect 32140 6934 32168 7278
rect 32128 6928 32180 6934
rect 32128 6870 32180 6876
rect 32140 6458 32168 6870
rect 32128 6452 32180 6458
rect 32128 6394 32180 6400
rect 32600 6322 32628 7890
rect 32968 7886 32996 8230
rect 33612 7886 33640 8366
rect 34244 8288 34296 8294
rect 34244 8230 34296 8236
rect 34704 8288 34756 8294
rect 34704 8230 34756 8236
rect 34256 8090 34284 8230
rect 34244 8084 34296 8090
rect 34244 8026 34296 8032
rect 32956 7880 33008 7886
rect 32956 7822 33008 7828
rect 33600 7880 33652 7886
rect 33600 7822 33652 7828
rect 34428 7744 34480 7750
rect 34428 7686 34480 7692
rect 34440 7410 34468 7686
rect 34716 7410 34744 8230
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35360 8090 35388 9522
rect 35440 8832 35492 8838
rect 35440 8774 35492 8780
rect 35452 8566 35480 8774
rect 35440 8560 35492 8566
rect 35440 8502 35492 8508
rect 34796 8084 34848 8090
rect 34796 8026 34848 8032
rect 35348 8084 35400 8090
rect 35348 8026 35400 8032
rect 34808 7818 34836 8026
rect 35452 7954 35480 8502
rect 35440 7948 35492 7954
rect 35440 7890 35492 7896
rect 34796 7812 34848 7818
rect 34796 7754 34848 7760
rect 34428 7404 34480 7410
rect 34428 7346 34480 7352
rect 34704 7404 34756 7410
rect 34704 7346 34756 7352
rect 33324 7200 33376 7206
rect 33324 7142 33376 7148
rect 32772 6928 32824 6934
rect 32772 6870 32824 6876
rect 32588 6316 32640 6322
rect 32588 6258 32640 6264
rect 32784 5914 32812 6870
rect 33336 6390 33364 7142
rect 34808 7002 34836 7754
rect 35348 7404 35400 7410
rect 35348 7346 35400 7352
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34796 6996 34848 7002
rect 34796 6938 34848 6944
rect 35360 6798 35388 7346
rect 35452 7342 35480 7890
rect 35532 7880 35584 7886
rect 35532 7822 35584 7828
rect 35544 7546 35572 7822
rect 35532 7540 35584 7546
rect 35532 7482 35584 7488
rect 35440 7336 35492 7342
rect 35440 7278 35492 7284
rect 35636 6866 35664 13942
rect 36004 13530 36032 14010
rect 35992 13524 36044 13530
rect 35992 13466 36044 13472
rect 36464 13258 36492 14758
rect 37200 14482 37228 14962
rect 37280 14952 37332 14958
rect 37280 14894 37332 14900
rect 37292 14618 37320 14894
rect 37280 14612 37332 14618
rect 37280 14554 37332 14560
rect 37188 14476 37240 14482
rect 37188 14418 37240 14424
rect 37292 14346 37320 14554
rect 37280 14340 37332 14346
rect 37280 14282 37332 14288
rect 37292 13870 37320 14282
rect 38120 14278 38148 16390
rect 38384 15700 38436 15706
rect 38384 15642 38436 15648
rect 37372 14272 37424 14278
rect 37372 14214 37424 14220
rect 38108 14272 38160 14278
rect 38108 14214 38160 14220
rect 37384 13938 37412 14214
rect 37372 13932 37424 13938
rect 37372 13874 37424 13880
rect 37280 13864 37332 13870
rect 37280 13806 37332 13812
rect 38120 13530 38148 14214
rect 38396 13530 38424 15642
rect 38856 15162 38884 16390
rect 39672 15428 39724 15434
rect 39672 15370 39724 15376
rect 38844 15156 38896 15162
rect 38844 15098 38896 15104
rect 38752 14952 38804 14958
rect 38752 14894 38804 14900
rect 38764 14414 38792 14894
rect 38476 14408 38528 14414
rect 38476 14350 38528 14356
rect 38752 14408 38804 14414
rect 38752 14350 38804 14356
rect 38488 13938 38516 14350
rect 38476 13932 38528 13938
rect 38476 13874 38528 13880
rect 38752 13932 38804 13938
rect 38752 13874 38804 13880
rect 38108 13524 38160 13530
rect 38108 13466 38160 13472
rect 38384 13524 38436 13530
rect 38384 13466 38436 13472
rect 36452 13252 36504 13258
rect 36452 13194 36504 13200
rect 36544 13252 36596 13258
rect 36544 13194 36596 13200
rect 36556 12986 36584 13194
rect 36544 12980 36596 12986
rect 36544 12922 36596 12928
rect 38488 12918 38516 13874
rect 38764 13530 38792 13874
rect 38752 13524 38804 13530
rect 38752 13466 38804 13472
rect 38856 13258 38884 15098
rect 39212 15020 39264 15026
rect 39212 14962 39264 14968
rect 39120 14816 39172 14822
rect 39120 14758 39172 14764
rect 39132 13326 39160 14758
rect 39224 14618 39252 14962
rect 39212 14612 39264 14618
rect 39212 14554 39264 14560
rect 39684 14006 39712 15370
rect 39776 15162 39804 19246
rect 40144 18766 40172 19314
rect 40604 18970 40632 19722
rect 40696 19514 40724 19722
rect 40684 19508 40736 19514
rect 40684 19450 40736 19456
rect 40684 19372 40736 19378
rect 40684 19314 40736 19320
rect 40592 18964 40644 18970
rect 40592 18906 40644 18912
rect 40696 18766 40724 19314
rect 40132 18760 40184 18766
rect 40132 18702 40184 18708
rect 40684 18760 40736 18766
rect 40684 18702 40736 18708
rect 40132 17672 40184 17678
rect 40132 17614 40184 17620
rect 39856 17536 39908 17542
rect 39856 17478 39908 17484
rect 39868 17202 39896 17478
rect 39856 17196 39908 17202
rect 39856 17138 39908 17144
rect 40040 16992 40092 16998
rect 40040 16934 40092 16940
rect 40052 16590 40080 16934
rect 40040 16584 40092 16590
rect 40040 16526 40092 16532
rect 40144 16454 40172 17614
rect 41524 16726 41552 25638
rect 43640 24410 43668 26386
rect 43628 24404 43680 24410
rect 43628 24346 43680 24352
rect 42524 24132 42576 24138
rect 42524 24074 42576 24080
rect 42248 24064 42300 24070
rect 42248 24006 42300 24012
rect 42340 24064 42392 24070
rect 42340 24006 42392 24012
rect 42260 23254 42288 24006
rect 42352 23866 42380 24006
rect 42536 23866 42564 24074
rect 42340 23860 42392 23866
rect 42340 23802 42392 23808
rect 42524 23860 42576 23866
rect 42524 23802 42576 23808
rect 43640 23730 43668 24346
rect 44100 24138 44128 35866
rect 65654 35388 65962 35397
rect 65654 35386 65660 35388
rect 65716 35386 65740 35388
rect 65796 35386 65820 35388
rect 65876 35386 65900 35388
rect 65956 35386 65962 35388
rect 65716 35334 65718 35386
rect 65898 35334 65900 35386
rect 65654 35332 65660 35334
rect 65716 35332 65740 35334
rect 65796 35332 65820 35334
rect 65876 35332 65900 35334
rect 65956 35332 65962 35334
rect 65654 35323 65962 35332
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 65654 34300 65962 34309
rect 65654 34298 65660 34300
rect 65716 34298 65740 34300
rect 65796 34298 65820 34300
rect 65876 34298 65900 34300
rect 65956 34298 65962 34300
rect 65716 34246 65718 34298
rect 65898 34246 65900 34298
rect 65654 34244 65660 34246
rect 65716 34244 65740 34246
rect 65796 34244 65820 34246
rect 65876 34244 65900 34246
rect 65956 34244 65962 34246
rect 65654 34235 65962 34244
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 65654 33212 65962 33221
rect 65654 33210 65660 33212
rect 65716 33210 65740 33212
rect 65796 33210 65820 33212
rect 65876 33210 65900 33212
rect 65956 33210 65962 33212
rect 65716 33158 65718 33210
rect 65898 33158 65900 33210
rect 65654 33156 65660 33158
rect 65716 33156 65740 33158
rect 65796 33156 65820 33158
rect 65876 33156 65900 33158
rect 65956 33156 65962 33158
rect 65654 33147 65962 33156
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 65654 32124 65962 32133
rect 65654 32122 65660 32124
rect 65716 32122 65740 32124
rect 65796 32122 65820 32124
rect 65876 32122 65900 32124
rect 65956 32122 65962 32124
rect 65716 32070 65718 32122
rect 65898 32070 65900 32122
rect 65654 32068 65660 32070
rect 65716 32068 65740 32070
rect 65796 32068 65820 32070
rect 65876 32068 65900 32070
rect 65956 32068 65962 32070
rect 65654 32059 65962 32068
rect 57704 31816 57756 31822
rect 57704 31758 57756 31764
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 45284 29300 45336 29306
rect 45284 29242 45336 29248
rect 45008 29164 45060 29170
rect 45008 29106 45060 29112
rect 44272 28960 44324 28966
rect 44272 28902 44324 28908
rect 44284 28626 44312 28902
rect 44272 28620 44324 28626
rect 44272 28562 44324 28568
rect 45020 27606 45048 29106
rect 45296 28558 45324 29242
rect 45928 29096 45980 29102
rect 45928 29038 45980 29044
rect 45284 28552 45336 28558
rect 45284 28494 45336 28500
rect 45940 28218 45968 29038
rect 54576 28552 54628 28558
rect 54576 28494 54628 28500
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 45468 28212 45520 28218
rect 45468 28154 45520 28160
rect 45928 28212 45980 28218
rect 45928 28154 45980 28160
rect 45480 28082 45508 28154
rect 45836 28144 45888 28150
rect 45836 28086 45888 28092
rect 45468 28076 45520 28082
rect 45468 28018 45520 28024
rect 45192 28008 45244 28014
rect 45192 27950 45244 27956
rect 45204 27606 45232 27950
rect 45008 27600 45060 27606
rect 45008 27542 45060 27548
rect 45192 27600 45244 27606
rect 45192 27542 45244 27548
rect 45204 27130 45232 27542
rect 45480 27538 45508 28018
rect 45468 27532 45520 27538
rect 45468 27474 45520 27480
rect 45848 27130 45876 28086
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 45192 27124 45244 27130
rect 45192 27066 45244 27072
rect 45836 27124 45888 27130
rect 45836 27066 45888 27072
rect 45008 26988 45060 26994
rect 45008 26930 45060 26936
rect 45284 26988 45336 26994
rect 45284 26930 45336 26936
rect 45020 26586 45048 26930
rect 45008 26580 45060 26586
rect 45008 26522 45060 26528
rect 45296 26382 45324 26930
rect 45284 26376 45336 26382
rect 45284 26318 45336 26324
rect 45192 24948 45244 24954
rect 45192 24890 45244 24896
rect 45008 24812 45060 24818
rect 45008 24754 45060 24760
rect 44180 24608 44232 24614
rect 44180 24550 44232 24556
rect 44088 24132 44140 24138
rect 44088 24074 44140 24080
rect 44192 23798 44220 24550
rect 45020 24410 45048 24754
rect 45008 24404 45060 24410
rect 45008 24346 45060 24352
rect 45204 24274 45232 24890
rect 45296 24818 45324 26318
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 45284 24812 45336 24818
rect 45284 24754 45336 24760
rect 45296 24342 45324 24754
rect 45836 24744 45888 24750
rect 45836 24686 45888 24692
rect 45468 24608 45520 24614
rect 45468 24550 45520 24556
rect 45284 24336 45336 24342
rect 45284 24278 45336 24284
rect 45192 24268 45244 24274
rect 45192 24210 45244 24216
rect 44272 24200 44324 24206
rect 44272 24142 44324 24148
rect 45284 24200 45336 24206
rect 45284 24142 45336 24148
rect 44180 23792 44232 23798
rect 44180 23734 44232 23740
rect 43260 23724 43312 23730
rect 43260 23666 43312 23672
rect 43628 23724 43680 23730
rect 43628 23666 43680 23672
rect 42800 23656 42852 23662
rect 42800 23598 42852 23604
rect 42812 23254 42840 23598
rect 43272 23322 43300 23666
rect 43260 23316 43312 23322
rect 43260 23258 43312 23264
rect 42248 23248 42300 23254
rect 42248 23190 42300 23196
rect 42800 23248 42852 23254
rect 42800 23190 42852 23196
rect 41880 23112 41932 23118
rect 41880 23054 41932 23060
rect 41892 22234 41920 23054
rect 42616 23044 42668 23050
rect 42616 22986 42668 22992
rect 42628 22545 42656 22986
rect 43640 22642 43668 23666
rect 44284 23662 44312 24142
rect 44732 24132 44784 24138
rect 44732 24074 44784 24080
rect 44640 24064 44692 24070
rect 44640 24006 44692 24012
rect 44652 23798 44680 24006
rect 44640 23792 44692 23798
rect 44640 23734 44692 23740
rect 44272 23656 44324 23662
rect 44272 23598 44324 23604
rect 44548 23520 44600 23526
rect 44548 23462 44600 23468
rect 43720 23248 43772 23254
rect 43720 23190 43772 23196
rect 43732 22710 43760 23190
rect 44560 23118 44588 23462
rect 44548 23112 44600 23118
rect 44548 23054 44600 23060
rect 44180 22976 44232 22982
rect 44180 22918 44232 22924
rect 44192 22710 44220 22918
rect 43720 22704 43772 22710
rect 43720 22646 43772 22652
rect 44180 22704 44232 22710
rect 44180 22646 44232 22652
rect 43628 22636 43680 22642
rect 43628 22578 43680 22584
rect 41970 22536 42026 22545
rect 41970 22471 42026 22480
rect 42614 22536 42670 22545
rect 42614 22471 42670 22480
rect 41880 22228 41932 22234
rect 41880 22170 41932 22176
rect 41880 21956 41932 21962
rect 41880 21898 41932 21904
rect 41892 21146 41920 21898
rect 41880 21140 41932 21146
rect 41880 21082 41932 21088
rect 41604 20800 41656 20806
rect 41604 20742 41656 20748
rect 41616 20330 41644 20742
rect 41604 20324 41656 20330
rect 41604 20266 41656 20272
rect 41616 18222 41644 20266
rect 41880 18760 41932 18766
rect 41880 18702 41932 18708
rect 41604 18216 41656 18222
rect 41604 18158 41656 18164
rect 41604 17536 41656 17542
rect 41604 17478 41656 17484
rect 41616 17202 41644 17478
rect 41604 17196 41656 17202
rect 41604 17138 41656 17144
rect 41788 17128 41840 17134
rect 41788 17070 41840 17076
rect 41512 16720 41564 16726
rect 41512 16662 41564 16668
rect 40316 16652 40368 16658
rect 40316 16594 40368 16600
rect 40132 16448 40184 16454
rect 40132 16390 40184 16396
rect 40040 15700 40092 15706
rect 40040 15642 40092 15648
rect 39764 15156 39816 15162
rect 39764 15098 39816 15104
rect 40052 15094 40080 15642
rect 40328 15638 40356 16594
rect 41052 16584 41104 16590
rect 41052 16526 41104 16532
rect 40408 16448 40460 16454
rect 40408 16390 40460 16396
rect 40316 15632 40368 15638
rect 40316 15574 40368 15580
rect 40040 15088 40092 15094
rect 40040 15030 40092 15036
rect 40328 14618 40356 15574
rect 40420 15366 40448 16390
rect 40408 15360 40460 15366
rect 40408 15302 40460 15308
rect 40420 15162 40448 15302
rect 41064 15162 41092 16526
rect 41328 15700 41380 15706
rect 41328 15642 41380 15648
rect 40408 15156 40460 15162
rect 40408 15098 40460 15104
rect 41052 15156 41104 15162
rect 41052 15098 41104 15104
rect 41340 15026 41368 15642
rect 41800 15638 41828 17070
rect 41892 16998 41920 18702
rect 41984 17542 42012 22471
rect 44272 21548 44324 21554
rect 44272 21490 44324 21496
rect 43812 21480 43864 21486
rect 43812 21422 43864 21428
rect 42340 21344 42392 21350
rect 42340 21286 42392 21292
rect 42352 20942 42380 21286
rect 42432 21072 42484 21078
rect 42432 21014 42484 21020
rect 42340 20936 42392 20942
rect 42340 20878 42392 20884
rect 42444 20466 42472 21014
rect 42616 21004 42668 21010
rect 42616 20946 42668 20952
rect 42628 20602 42656 20946
rect 42800 20936 42852 20942
rect 42800 20878 42852 20884
rect 42812 20806 42840 20878
rect 42708 20800 42760 20806
rect 42708 20742 42760 20748
rect 42800 20800 42852 20806
rect 42800 20742 42852 20748
rect 42616 20596 42668 20602
rect 42616 20538 42668 20544
rect 42720 20466 42748 20742
rect 42432 20460 42484 20466
rect 42432 20402 42484 20408
rect 42708 20460 42760 20466
rect 42708 20402 42760 20408
rect 42720 20058 42748 20402
rect 42708 20052 42760 20058
rect 42708 19994 42760 20000
rect 42812 19922 42840 20742
rect 43824 20534 43852 21422
rect 43904 21344 43956 21350
rect 43904 21286 43956 21292
rect 43812 20528 43864 20534
rect 43812 20470 43864 20476
rect 43352 20392 43404 20398
rect 43352 20334 43404 20340
rect 43076 20256 43128 20262
rect 43076 20198 43128 20204
rect 42800 19916 42852 19922
rect 42800 19858 42852 19864
rect 43088 19854 43116 20198
rect 43076 19848 43128 19854
rect 43076 19790 43128 19796
rect 42432 19780 42484 19786
rect 42432 19722 42484 19728
rect 41972 17536 42024 17542
rect 41972 17478 42024 17484
rect 42156 17060 42208 17066
rect 42156 17002 42208 17008
rect 41880 16992 41932 16998
rect 41880 16934 41932 16940
rect 41788 15632 41840 15638
rect 41788 15574 41840 15580
rect 41604 15564 41656 15570
rect 41604 15506 41656 15512
rect 41512 15360 41564 15366
rect 41512 15302 41564 15308
rect 41524 15026 41552 15302
rect 41616 15094 41644 15506
rect 41604 15088 41656 15094
rect 41604 15030 41656 15036
rect 40408 15020 40460 15026
rect 40408 14962 40460 14968
rect 41328 15020 41380 15026
rect 41328 14962 41380 14968
rect 41512 15020 41564 15026
rect 41512 14962 41564 14968
rect 40420 14618 40448 14962
rect 41144 14884 41196 14890
rect 41144 14826 41196 14832
rect 40316 14612 40368 14618
rect 40316 14554 40368 14560
rect 40408 14612 40460 14618
rect 40408 14554 40460 14560
rect 41156 14414 41184 14826
rect 39856 14408 39908 14414
rect 39856 14350 39908 14356
rect 40040 14408 40092 14414
rect 40040 14350 40092 14356
rect 40868 14408 40920 14414
rect 40868 14350 40920 14356
rect 41144 14408 41196 14414
rect 41144 14350 41196 14356
rect 39868 14074 39896 14350
rect 39856 14068 39908 14074
rect 39856 14010 39908 14016
rect 39672 14000 39724 14006
rect 39672 13942 39724 13948
rect 39856 13864 39908 13870
rect 39856 13806 39908 13812
rect 39868 13394 39896 13806
rect 39856 13388 39908 13394
rect 39856 13330 39908 13336
rect 39120 13320 39172 13326
rect 39120 13262 39172 13268
rect 38844 13252 38896 13258
rect 38844 13194 38896 13200
rect 40052 12986 40080 14350
rect 40880 13870 40908 14350
rect 41696 14272 41748 14278
rect 41696 14214 41748 14220
rect 41708 13938 41736 14214
rect 41696 13932 41748 13938
rect 41696 13874 41748 13880
rect 40868 13864 40920 13870
rect 40868 13806 40920 13812
rect 41604 13864 41656 13870
rect 41604 13806 41656 13812
rect 41420 13184 41472 13190
rect 41420 13126 41472 13132
rect 40040 12980 40092 12986
rect 40040 12922 40092 12928
rect 36360 12912 36412 12918
rect 36360 12854 36412 12860
rect 38476 12912 38528 12918
rect 38476 12854 38528 12860
rect 41236 12912 41288 12918
rect 41236 12854 41288 12860
rect 36372 12306 36400 12854
rect 37740 12640 37792 12646
rect 37740 12582 37792 12588
rect 38200 12640 38252 12646
rect 38200 12582 38252 12588
rect 37752 12442 37780 12582
rect 37740 12436 37792 12442
rect 37740 12378 37792 12384
rect 36084 12300 36136 12306
rect 36084 12242 36136 12248
rect 36360 12300 36412 12306
rect 36360 12242 36412 12248
rect 36096 11558 36124 12242
rect 36912 12232 36964 12238
rect 36912 12174 36964 12180
rect 37188 12232 37240 12238
rect 37372 12232 37424 12238
rect 37240 12192 37372 12220
rect 37188 12174 37240 12180
rect 37372 12174 37424 12180
rect 36924 12102 36952 12174
rect 36912 12096 36964 12102
rect 36912 12038 36964 12044
rect 36924 11694 36952 12038
rect 37752 11898 37780 12378
rect 38212 12238 38240 12582
rect 38200 12232 38252 12238
rect 38200 12174 38252 12180
rect 37280 11892 37332 11898
rect 37280 11834 37332 11840
rect 37740 11892 37792 11898
rect 37740 11834 37792 11840
rect 36912 11688 36964 11694
rect 36912 11630 36964 11636
rect 36084 11552 36136 11558
rect 36084 11494 36136 11500
rect 36096 11354 36124 11494
rect 36084 11348 36136 11354
rect 36084 11290 36136 11296
rect 36924 11218 36952 11630
rect 36912 11212 36964 11218
rect 36912 11154 36964 11160
rect 37292 11150 37320 11834
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 37280 11144 37332 11150
rect 36174 11112 36230 11121
rect 37280 11086 37332 11092
rect 36174 11047 36176 11056
rect 36228 11047 36230 11056
rect 36176 11018 36228 11024
rect 37844 10674 37872 11494
rect 38212 11218 38240 12174
rect 38292 12096 38344 12102
rect 38292 12038 38344 12044
rect 38304 11830 38332 12038
rect 38488 11898 38516 12854
rect 38568 12844 38620 12850
rect 38568 12786 38620 12792
rect 38752 12844 38804 12850
rect 38752 12786 38804 12792
rect 40316 12844 40368 12850
rect 40316 12786 40368 12792
rect 38580 12238 38608 12786
rect 38764 12442 38792 12786
rect 38752 12436 38804 12442
rect 38752 12378 38804 12384
rect 38568 12232 38620 12238
rect 38568 12174 38620 12180
rect 38476 11892 38528 11898
rect 38476 11834 38528 11840
rect 38292 11824 38344 11830
rect 38292 11766 38344 11772
rect 38580 11354 38608 12174
rect 38568 11348 38620 11354
rect 38568 11290 38620 11296
rect 38200 11212 38252 11218
rect 38200 11154 38252 11160
rect 38212 10742 38240 11154
rect 38384 11144 38436 11150
rect 38384 11086 38436 11092
rect 38396 10742 38424 11086
rect 38200 10736 38252 10742
rect 38200 10678 38252 10684
rect 38384 10736 38436 10742
rect 38384 10678 38436 10684
rect 37832 10668 37884 10674
rect 37832 10610 37884 10616
rect 38764 10062 38792 12378
rect 40328 12374 40356 12786
rect 40316 12368 40368 12374
rect 40316 12310 40368 12316
rect 40132 12232 40184 12238
rect 40132 12174 40184 12180
rect 38936 11212 38988 11218
rect 38936 11154 38988 11160
rect 38948 10810 38976 11154
rect 39856 11144 39908 11150
rect 39856 11086 39908 11092
rect 38936 10804 38988 10810
rect 38936 10746 38988 10752
rect 39028 10464 39080 10470
rect 39028 10406 39080 10412
rect 38108 10056 38160 10062
rect 38108 9998 38160 10004
rect 38752 10056 38804 10062
rect 38752 9998 38804 10004
rect 36452 9920 36504 9926
rect 36452 9862 36504 9868
rect 35716 9512 35768 9518
rect 35716 9454 35768 9460
rect 35728 8294 35756 9454
rect 35808 9104 35860 9110
rect 35808 9046 35860 9052
rect 35716 8288 35768 8294
rect 35716 8230 35768 8236
rect 35728 8090 35756 8230
rect 35716 8084 35768 8090
rect 35716 8026 35768 8032
rect 35624 6860 35676 6866
rect 35624 6802 35676 6808
rect 34796 6792 34848 6798
rect 34796 6734 34848 6740
rect 35348 6792 35400 6798
rect 35348 6734 35400 6740
rect 34808 6458 34836 6734
rect 34796 6452 34848 6458
rect 34796 6394 34848 6400
rect 33324 6384 33376 6390
rect 33324 6326 33376 6332
rect 33876 6384 33928 6390
rect 33876 6326 33928 6332
rect 33888 5914 33916 6326
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 32772 5908 32824 5914
rect 32772 5850 32824 5856
rect 33876 5908 33928 5914
rect 33876 5850 33928 5856
rect 35820 5778 35848 9046
rect 36464 8906 36492 9862
rect 38120 9722 38148 9998
rect 38108 9716 38160 9722
rect 38108 9658 38160 9664
rect 36728 9376 36780 9382
rect 36728 9318 36780 9324
rect 36740 9178 36768 9318
rect 36728 9172 36780 9178
rect 36728 9114 36780 9120
rect 36452 8900 36504 8906
rect 36452 8842 36504 8848
rect 36912 8900 36964 8906
rect 36912 8842 36964 8848
rect 36924 8634 36952 8842
rect 36912 8628 36964 8634
rect 36912 8570 36964 8576
rect 38014 7576 38070 7585
rect 38014 7511 38070 7520
rect 38028 7410 38056 7511
rect 38016 7404 38068 7410
rect 38016 7346 38068 7352
rect 37464 7200 37516 7206
rect 37464 7142 37516 7148
rect 37476 7002 37504 7142
rect 37464 6996 37516 7002
rect 37464 6938 37516 6944
rect 37372 6112 37424 6118
rect 37372 6054 37424 6060
rect 35808 5772 35860 5778
rect 35808 5714 35860 5720
rect 33784 5704 33836 5710
rect 33784 5646 33836 5652
rect 32680 5636 32732 5642
rect 32680 5578 32732 5584
rect 32692 5370 32720 5578
rect 32680 5364 32732 5370
rect 32680 5306 32732 5312
rect 33796 5234 33824 5646
rect 33784 5228 33836 5234
rect 33784 5170 33836 5176
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 31772 4780 31892 4808
rect 31116 4616 31168 4622
rect 31116 4558 31168 4564
rect 31024 3460 31076 3466
rect 31024 3402 31076 3408
rect 31036 3194 31064 3402
rect 31024 3188 31076 3194
rect 31024 3130 31076 3136
rect 30748 2508 30800 2514
rect 30748 2450 30800 2456
rect 30656 2372 30708 2378
rect 30656 2314 30708 2320
rect 30760 800 30788 2450
rect 31128 1442 31156 4558
rect 31772 4146 31800 4780
rect 35820 4622 35848 5714
rect 37384 5710 37412 6054
rect 37476 5914 37504 6938
rect 38660 6316 38712 6322
rect 38660 6258 38712 6264
rect 37464 5908 37516 5914
rect 37464 5850 37516 5856
rect 37372 5704 37424 5710
rect 37372 5646 37424 5652
rect 35900 5636 35952 5642
rect 35900 5578 35952 5584
rect 35912 5370 35940 5578
rect 37280 5568 37332 5574
rect 37280 5510 37332 5516
rect 37372 5568 37424 5574
rect 37372 5510 37424 5516
rect 37292 5370 37320 5510
rect 35900 5364 35952 5370
rect 35900 5306 35952 5312
rect 37280 5364 37332 5370
rect 37280 5306 37332 5312
rect 37188 5024 37240 5030
rect 37188 4966 37240 4972
rect 37200 4622 37228 4966
rect 31852 4616 31904 4622
rect 35808 4616 35860 4622
rect 31852 4558 31904 4564
rect 33046 4584 33102 4593
rect 31760 4140 31812 4146
rect 31760 4082 31812 4088
rect 31484 3936 31536 3942
rect 31484 3878 31536 3884
rect 31496 3466 31524 3878
rect 31576 3732 31628 3738
rect 31576 3674 31628 3680
rect 31484 3460 31536 3466
rect 31484 3402 31536 3408
rect 31300 2440 31352 2446
rect 31300 2382 31352 2388
rect 31036 1414 31156 1442
rect 31036 800 31064 1414
rect 31312 800 31340 2382
rect 31588 800 31616 3674
rect 31864 800 31892 4558
rect 35808 4558 35860 4564
rect 37188 4616 37240 4622
rect 37188 4558 37240 4564
rect 33046 4519 33102 4528
rect 32956 4480 33008 4486
rect 32956 4422 33008 4428
rect 32968 4078 32996 4422
rect 33060 4282 33088 4519
rect 33048 4276 33100 4282
rect 33048 4218 33100 4224
rect 32128 4072 32180 4078
rect 32128 4014 32180 4020
rect 32956 4072 33008 4078
rect 32956 4014 33008 4020
rect 32140 3194 32168 4014
rect 32220 3936 32272 3942
rect 32220 3878 32272 3884
rect 32128 3188 32180 3194
rect 32128 3130 32180 3136
rect 32232 3058 32260 3878
rect 32588 3732 32640 3738
rect 32588 3674 32640 3680
rect 32312 3596 32364 3602
rect 32312 3538 32364 3544
rect 32220 3052 32272 3058
rect 32220 2994 32272 3000
rect 32324 1850 32352 3538
rect 32600 3194 32628 3674
rect 32588 3188 32640 3194
rect 32588 3130 32640 3136
rect 32968 2990 32996 4014
rect 33060 3738 33088 4218
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 33048 3732 33100 3738
rect 33048 3674 33100 3680
rect 35820 3602 35848 4558
rect 36084 4548 36136 4554
rect 36084 4490 36136 4496
rect 36096 4282 36124 4490
rect 36084 4276 36136 4282
rect 36084 4218 36136 4224
rect 37384 4146 37412 5510
rect 37476 4146 37504 5850
rect 38384 5772 38436 5778
rect 38384 5714 38436 5720
rect 38108 5568 38160 5574
rect 38108 5510 38160 5516
rect 38120 5234 38148 5510
rect 38108 5228 38160 5234
rect 38108 5170 38160 5176
rect 38120 4758 38148 5170
rect 38396 5166 38424 5714
rect 38672 5273 38700 6258
rect 38844 5568 38896 5574
rect 38844 5510 38896 5516
rect 38658 5264 38714 5273
rect 38856 5234 38884 5510
rect 38658 5199 38660 5208
rect 38712 5199 38714 5208
rect 38844 5228 38896 5234
rect 38660 5170 38712 5176
rect 38844 5170 38896 5176
rect 38384 5160 38436 5166
rect 38384 5102 38436 5108
rect 38108 4752 38160 4758
rect 38108 4694 38160 4700
rect 38752 4616 38804 4622
rect 38752 4558 38804 4564
rect 38658 4312 38714 4321
rect 38658 4247 38714 4256
rect 37372 4140 37424 4146
rect 37372 4082 37424 4088
rect 37464 4140 37516 4146
rect 37464 4082 37516 4088
rect 37924 4072 37976 4078
rect 37924 4014 37976 4020
rect 37372 3936 37424 3942
rect 37372 3878 37424 3884
rect 37648 3936 37700 3942
rect 37648 3878 37700 3884
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 37384 3534 37412 3878
rect 33232 3528 33284 3534
rect 33232 3470 33284 3476
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 32772 2984 32824 2990
rect 32772 2926 32824 2932
rect 32956 2984 33008 2990
rect 32956 2926 33008 2932
rect 32784 2650 32812 2926
rect 32772 2644 32824 2650
rect 32772 2586 32824 2592
rect 32404 2576 32456 2582
rect 32404 2518 32456 2524
rect 32140 1822 32352 1850
rect 32140 800 32168 1822
rect 32416 800 32444 2518
rect 32680 2508 32732 2514
rect 32680 2450 32732 2456
rect 32692 800 32720 2450
rect 32956 2440 33008 2446
rect 32956 2382 33008 2388
rect 32968 800 32996 2382
rect 33244 800 33272 3470
rect 33784 2848 33836 2854
rect 33784 2790 33836 2796
rect 34336 2848 34388 2854
rect 34336 2790 34388 2796
rect 34796 2848 34848 2854
rect 34796 2790 34848 2796
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 36268 2848 36320 2854
rect 36268 2790 36320 2796
rect 36820 2848 36872 2854
rect 36820 2790 36872 2796
rect 33508 2576 33560 2582
rect 33508 2518 33560 2524
rect 33520 800 33548 2518
rect 33796 800 33824 2790
rect 34060 2440 34112 2446
rect 34060 2382 34112 2388
rect 34072 800 34100 2382
rect 34348 800 34376 2790
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 34624 800 34652 2382
rect 34808 1442 34836 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35164 2440 35216 2446
rect 35164 2382 35216 2388
rect 34808 1414 34928 1442
rect 34900 800 34928 1414
rect 35176 800 35204 2382
rect 35452 800 35480 2790
rect 35716 2440 35768 2446
rect 35716 2382 35768 2388
rect 35992 2440 36044 2446
rect 35992 2382 36044 2388
rect 35728 800 35756 2382
rect 36004 800 36032 2382
rect 36280 800 36308 2790
rect 36544 2440 36596 2446
rect 36544 2382 36596 2388
rect 36556 800 36584 2382
rect 36832 800 36860 2790
rect 37096 2508 37148 2514
rect 37096 2450 37148 2456
rect 37108 800 37136 2450
rect 37372 2440 37424 2446
rect 37372 2382 37424 2388
rect 37384 800 37412 2382
rect 37660 800 37688 3878
rect 37936 800 37964 4014
rect 38476 3936 38528 3942
rect 38476 3878 38528 3884
rect 38200 2916 38252 2922
rect 38200 2858 38252 2864
rect 38212 800 38240 2858
rect 38488 800 38516 3878
rect 38568 3528 38620 3534
rect 38568 3470 38620 3476
rect 38580 2990 38608 3470
rect 38568 2984 38620 2990
rect 38568 2926 38620 2932
rect 38672 2922 38700 4247
rect 38660 2916 38712 2922
rect 38660 2858 38712 2864
rect 38764 800 38792 4558
rect 38856 4214 38884 5170
rect 38936 4684 38988 4690
rect 38936 4626 38988 4632
rect 38844 4208 38896 4214
rect 38844 4150 38896 4156
rect 38856 3194 38884 4150
rect 38844 3188 38896 3194
rect 38844 3130 38896 3136
rect 38948 2292 38976 4626
rect 39040 4010 39068 10406
rect 39212 9376 39264 9382
rect 39212 9318 39264 9324
rect 39224 7886 39252 9318
rect 39580 8288 39632 8294
rect 39580 8230 39632 8236
rect 39212 7880 39264 7886
rect 39212 7822 39264 7828
rect 39592 7478 39620 8230
rect 39580 7472 39632 7478
rect 39580 7414 39632 7420
rect 39304 5704 39356 5710
rect 39304 5646 39356 5652
rect 39028 4004 39080 4010
rect 39028 3946 39080 3952
rect 39040 3534 39068 3946
rect 39028 3528 39080 3534
rect 39028 3470 39080 3476
rect 39028 3392 39080 3398
rect 39028 3334 39080 3340
rect 39040 3126 39068 3334
rect 39028 3120 39080 3126
rect 39028 3062 39080 3068
rect 38948 2264 39068 2292
rect 39040 800 39068 2264
rect 39316 800 39344 5646
rect 39868 5642 39896 11086
rect 40040 10056 40092 10062
rect 40040 9998 40092 10004
rect 39948 9920 40000 9926
rect 39948 9862 40000 9868
rect 39960 9654 39988 9862
rect 40052 9722 40080 9998
rect 40040 9716 40092 9722
rect 40040 9658 40092 9664
rect 39948 9648 40000 9654
rect 39948 9590 40000 9596
rect 40052 8498 40080 9658
rect 40040 8492 40092 8498
rect 40040 8434 40092 8440
rect 40144 7970 40172 12174
rect 40684 12096 40736 12102
rect 40684 12038 40736 12044
rect 40500 10668 40552 10674
rect 40500 10610 40552 10616
rect 40512 10266 40540 10610
rect 40592 10532 40644 10538
rect 40592 10474 40644 10480
rect 40500 10260 40552 10266
rect 40500 10202 40552 10208
rect 40316 9988 40368 9994
rect 40316 9930 40368 9936
rect 40328 9654 40356 9930
rect 40316 9648 40368 9654
rect 40316 9590 40368 9596
rect 40224 9512 40276 9518
rect 40224 9454 40276 9460
rect 40236 8634 40264 9454
rect 40328 9042 40356 9590
rect 40316 9036 40368 9042
rect 40316 8978 40368 8984
rect 40224 8628 40276 8634
rect 40224 8570 40276 8576
rect 40224 8356 40276 8362
rect 40224 8298 40276 8304
rect 40236 8090 40264 8298
rect 40224 8084 40276 8090
rect 40224 8026 40276 8032
rect 39960 7942 40172 7970
rect 39960 6934 39988 7942
rect 40040 7812 40092 7818
rect 40040 7754 40092 7760
rect 40052 6934 40080 7754
rect 40328 7478 40356 8978
rect 40500 8900 40552 8906
rect 40500 8842 40552 8848
rect 40512 8634 40540 8842
rect 40500 8628 40552 8634
rect 40500 8570 40552 8576
rect 40408 7812 40460 7818
rect 40460 7772 40540 7800
rect 40408 7754 40460 7760
rect 40316 7472 40368 7478
rect 40316 7414 40368 7420
rect 40224 7336 40276 7342
rect 40224 7278 40276 7284
rect 40132 7200 40184 7206
rect 40132 7142 40184 7148
rect 39948 6928 40000 6934
rect 39948 6870 40000 6876
rect 40040 6928 40092 6934
rect 40040 6870 40092 6876
rect 40040 6248 40092 6254
rect 40040 6190 40092 6196
rect 39856 5636 39908 5642
rect 39856 5578 39908 5584
rect 39764 5568 39816 5574
rect 39764 5510 39816 5516
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 39592 800 39620 3674
rect 39776 3126 39804 5510
rect 40052 5370 40080 6190
rect 40144 5778 40172 7142
rect 40236 7002 40264 7278
rect 40512 7002 40540 7772
rect 40224 6996 40276 7002
rect 40224 6938 40276 6944
rect 40500 6996 40552 7002
rect 40500 6938 40552 6944
rect 40512 6798 40540 6938
rect 40500 6792 40552 6798
rect 40500 6734 40552 6740
rect 40224 6248 40276 6254
rect 40224 6190 40276 6196
rect 40316 6248 40368 6254
rect 40316 6190 40368 6196
rect 40132 5772 40184 5778
rect 40132 5714 40184 5720
rect 40040 5364 40092 5370
rect 40040 5306 40092 5312
rect 39948 5228 40000 5234
rect 39948 5170 40000 5176
rect 39856 4480 39908 4486
rect 39856 4422 39908 4428
rect 39868 4146 39896 4422
rect 39960 4321 39988 5170
rect 40144 5098 40172 5714
rect 40132 5092 40184 5098
rect 40132 5034 40184 5040
rect 40236 4826 40264 6190
rect 40328 5098 40356 6190
rect 40408 5704 40460 5710
rect 40408 5646 40460 5652
rect 40316 5092 40368 5098
rect 40316 5034 40368 5040
rect 40224 4820 40276 4826
rect 40224 4762 40276 4768
rect 39946 4312 40002 4321
rect 39946 4247 40002 4256
rect 39856 4140 39908 4146
rect 39908 4100 39988 4128
rect 39856 4082 39908 4088
rect 39856 4004 39908 4010
rect 39856 3946 39908 3952
rect 39868 3913 39896 3946
rect 39854 3904 39910 3913
rect 39854 3839 39910 3848
rect 39856 3528 39908 3534
rect 39856 3470 39908 3476
rect 39868 3194 39896 3470
rect 39856 3188 39908 3194
rect 39856 3130 39908 3136
rect 39764 3120 39816 3126
rect 39764 3062 39816 3068
rect 39960 2514 39988 4100
rect 40420 4010 40448 5646
rect 40604 5273 40632 10474
rect 40696 6730 40724 12038
rect 40776 11076 40828 11082
rect 40776 11018 40828 11024
rect 40788 10810 40816 11018
rect 40776 10804 40828 10810
rect 40776 10746 40828 10752
rect 41248 10198 41276 12854
rect 41432 12322 41460 13126
rect 41340 12294 41460 12322
rect 41340 12102 41368 12294
rect 41328 12096 41380 12102
rect 41328 12038 41380 12044
rect 41616 11898 41644 13806
rect 41604 11892 41656 11898
rect 41604 11834 41656 11840
rect 41420 11756 41472 11762
rect 41420 11698 41472 11704
rect 41432 10674 41460 11698
rect 41616 11218 41644 11834
rect 41892 11762 41920 16934
rect 42168 16590 42196 17002
rect 42444 16794 42472 19722
rect 43364 19378 43392 20334
rect 43824 19990 43852 20470
rect 43812 19984 43864 19990
rect 43812 19926 43864 19932
rect 43628 19712 43680 19718
rect 43628 19654 43680 19660
rect 43640 19446 43668 19654
rect 43628 19440 43680 19446
rect 43628 19382 43680 19388
rect 43352 19372 43404 19378
rect 43352 19314 43404 19320
rect 43076 17672 43128 17678
rect 43076 17614 43128 17620
rect 42708 17536 42760 17542
rect 42708 17478 42760 17484
rect 42616 17332 42668 17338
rect 42616 17274 42668 17280
rect 42432 16788 42484 16794
rect 42432 16730 42484 16736
rect 42156 16584 42208 16590
rect 42208 16544 42288 16572
rect 42156 16526 42208 16532
rect 42260 13530 42288 16544
rect 42628 16522 42656 17274
rect 42616 16516 42668 16522
rect 42616 16458 42668 16464
rect 42628 16250 42656 16458
rect 42616 16244 42668 16250
rect 42616 16186 42668 16192
rect 42432 16040 42484 16046
rect 42432 15982 42484 15988
rect 42444 14958 42472 15982
rect 42628 15706 42656 16186
rect 42616 15700 42668 15706
rect 42616 15642 42668 15648
rect 42432 14952 42484 14958
rect 42432 14894 42484 14900
rect 42444 13870 42472 14894
rect 42628 14414 42656 15642
rect 42616 14408 42668 14414
rect 42616 14350 42668 14356
rect 42432 13864 42484 13870
rect 42432 13806 42484 13812
rect 42248 13524 42300 13530
rect 42248 13466 42300 13472
rect 42720 12434 42748 17478
rect 43088 16794 43116 17614
rect 43260 17536 43312 17542
rect 43260 17478 43312 17484
rect 43272 17270 43300 17478
rect 43260 17264 43312 17270
rect 43260 17206 43312 17212
rect 43364 17202 43392 19314
rect 43536 18080 43588 18086
rect 43536 18022 43588 18028
rect 43548 17610 43576 18022
rect 43812 17740 43864 17746
rect 43812 17682 43864 17688
rect 43536 17604 43588 17610
rect 43536 17546 43588 17552
rect 43352 17196 43404 17202
rect 43352 17138 43404 17144
rect 43076 16788 43128 16794
rect 43076 16730 43128 16736
rect 43260 16448 43312 16454
rect 43260 16390 43312 16396
rect 43272 15502 43300 16390
rect 43168 15496 43220 15502
rect 43168 15438 43220 15444
rect 43260 15496 43312 15502
rect 43260 15438 43312 15444
rect 43548 15450 43576 17546
rect 43720 17536 43772 17542
rect 43720 17478 43772 17484
rect 43732 16114 43760 17478
rect 43824 16794 43852 17682
rect 43812 16788 43864 16794
rect 43812 16730 43864 16736
rect 43824 16658 43852 16730
rect 43812 16652 43864 16658
rect 43812 16594 43864 16600
rect 43720 16108 43772 16114
rect 43720 16050 43772 16056
rect 43180 15026 43208 15438
rect 43272 15144 43300 15438
rect 43548 15422 43668 15450
rect 43536 15360 43588 15366
rect 43536 15302 43588 15308
rect 43272 15116 43392 15144
rect 43364 15026 43392 15116
rect 43548 15094 43576 15302
rect 43536 15088 43588 15094
rect 43536 15030 43588 15036
rect 43168 15020 43220 15026
rect 43168 14962 43220 14968
rect 43352 15020 43404 15026
rect 43352 14962 43404 14968
rect 43076 14272 43128 14278
rect 43076 14214 43128 14220
rect 43088 13734 43116 14214
rect 43180 14074 43208 14962
rect 43364 14346 43392 14962
rect 43352 14340 43404 14346
rect 43352 14282 43404 14288
rect 43168 14068 43220 14074
rect 43168 14010 43220 14016
rect 43076 13728 43128 13734
rect 43076 13670 43128 13676
rect 43088 13326 43116 13670
rect 43548 13530 43576 15030
rect 43640 14278 43668 15422
rect 43628 14272 43680 14278
rect 43628 14214 43680 14220
rect 43352 13524 43404 13530
rect 43352 13466 43404 13472
rect 43536 13524 43588 13530
rect 43536 13466 43588 13472
rect 43076 13320 43128 13326
rect 43076 13262 43128 13268
rect 43364 12986 43392 13466
rect 43352 12980 43404 12986
rect 43352 12922 43404 12928
rect 43640 12850 43668 14214
rect 43720 12980 43772 12986
rect 43720 12922 43772 12928
rect 43628 12844 43680 12850
rect 43628 12786 43680 12792
rect 42628 12406 42748 12434
rect 42156 11892 42208 11898
rect 42156 11834 42208 11840
rect 41880 11756 41932 11762
rect 41880 11698 41932 11704
rect 41604 11212 41656 11218
rect 41604 11154 41656 11160
rect 42168 11150 42196 11834
rect 42156 11144 42208 11150
rect 42156 11086 42208 11092
rect 41420 10668 41472 10674
rect 41420 10610 41472 10616
rect 41236 10192 41288 10198
rect 41236 10134 41288 10140
rect 41432 10130 41460 10610
rect 42628 10470 42656 12406
rect 43732 12238 43760 12922
rect 43916 12434 43944 21286
rect 44180 20800 44232 20806
rect 44180 20742 44232 20748
rect 44192 20534 44220 20742
rect 44180 20528 44232 20534
rect 44180 20470 44232 20476
rect 44284 20398 44312 21490
rect 44272 20392 44324 20398
rect 44272 20334 44324 20340
rect 44272 19440 44324 19446
rect 44272 19382 44324 19388
rect 44284 18970 44312 19382
rect 44272 18964 44324 18970
rect 44272 18906 44324 18912
rect 44744 17270 44772 24074
rect 45296 23186 45324 24142
rect 45284 23180 45336 23186
rect 45284 23122 45336 23128
rect 45296 22556 45324 23122
rect 45480 22710 45508 24550
rect 45848 24342 45876 24686
rect 45836 24336 45888 24342
rect 45836 24278 45888 24284
rect 46848 24336 46900 24342
rect 46848 24278 46900 24284
rect 45652 24064 45704 24070
rect 45652 24006 45704 24012
rect 45664 23322 45692 24006
rect 45652 23316 45704 23322
rect 45652 23258 45704 23264
rect 45848 23118 45876 24278
rect 46020 24268 46072 24274
rect 46020 24210 46072 24216
rect 46032 23662 46060 24210
rect 46860 23662 46888 24278
rect 46940 24064 46992 24070
rect 46940 24006 46992 24012
rect 46020 23656 46072 23662
rect 46020 23598 46072 23604
rect 46848 23656 46900 23662
rect 46848 23598 46900 23604
rect 46032 23254 46060 23598
rect 46952 23594 46980 24006
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 47584 23792 47636 23798
rect 47584 23734 47636 23740
rect 46940 23588 46992 23594
rect 46940 23530 46992 23536
rect 46020 23248 46072 23254
rect 46020 23190 46072 23196
rect 45836 23112 45888 23118
rect 45836 23054 45888 23060
rect 45468 22704 45520 22710
rect 45468 22646 45520 22652
rect 45376 22568 45428 22574
rect 45296 22528 45376 22556
rect 45376 22510 45428 22516
rect 45848 21622 45876 23054
rect 46032 22778 46060 23190
rect 46952 23186 46980 23530
rect 47400 23520 47452 23526
rect 47400 23462 47452 23468
rect 46940 23180 46992 23186
rect 46940 23122 46992 23128
rect 47412 23118 47440 23462
rect 47400 23112 47452 23118
rect 47400 23054 47452 23060
rect 47596 22982 47624 23734
rect 48688 23724 48740 23730
rect 48688 23666 48740 23672
rect 46112 22976 46164 22982
rect 46112 22918 46164 22924
rect 47584 22976 47636 22982
rect 47584 22918 47636 22924
rect 46020 22772 46072 22778
rect 46020 22714 46072 22720
rect 46124 22642 46152 22918
rect 47596 22642 47624 22918
rect 46112 22636 46164 22642
rect 46112 22578 46164 22584
rect 47584 22636 47636 22642
rect 47584 22578 47636 22584
rect 46020 22432 46072 22438
rect 46020 22374 46072 22380
rect 45836 21616 45888 21622
rect 45836 21558 45888 21564
rect 46032 21554 46060 22374
rect 46124 22098 46152 22578
rect 46112 22092 46164 22098
rect 46112 22034 46164 22040
rect 46020 21548 46072 21554
rect 46020 21490 46072 21496
rect 46848 21548 46900 21554
rect 46848 21490 46900 21496
rect 45008 21344 45060 21350
rect 45008 21286 45060 21292
rect 45020 20942 45048 21286
rect 46112 21140 46164 21146
rect 46112 21082 46164 21088
rect 45008 20936 45060 20942
rect 45008 20878 45060 20884
rect 45652 20936 45704 20942
rect 45652 20878 45704 20884
rect 45192 20800 45244 20806
rect 45192 20742 45244 20748
rect 45204 20466 45232 20742
rect 45008 20460 45060 20466
rect 45008 20402 45060 20408
rect 45192 20460 45244 20466
rect 45192 20402 45244 20408
rect 44916 20392 44968 20398
rect 44916 20334 44968 20340
rect 44928 19922 44956 20334
rect 44916 19916 44968 19922
rect 44916 19858 44968 19864
rect 45020 18970 45048 20402
rect 45192 20256 45244 20262
rect 45192 20198 45244 20204
rect 45100 19984 45152 19990
rect 45100 19926 45152 19932
rect 45112 19514 45140 19926
rect 45100 19508 45152 19514
rect 45100 19450 45152 19456
rect 45008 18964 45060 18970
rect 45008 18906 45060 18912
rect 44732 17264 44784 17270
rect 44732 17206 44784 17212
rect 44916 16992 44968 16998
rect 44916 16934 44968 16940
rect 45008 16992 45060 16998
rect 45008 16934 45060 16940
rect 44928 16522 44956 16934
rect 45020 16658 45048 16934
rect 45204 16726 45232 20198
rect 45664 20058 45692 20878
rect 46124 20806 46152 21082
rect 46112 20800 46164 20806
rect 46112 20742 46164 20748
rect 46124 20466 46152 20742
rect 46112 20460 46164 20466
rect 46112 20402 46164 20408
rect 45652 20052 45704 20058
rect 45652 19994 45704 20000
rect 45560 17536 45612 17542
rect 45560 17478 45612 17484
rect 45192 16720 45244 16726
rect 45192 16662 45244 16668
rect 45572 16658 45600 17478
rect 46020 17060 46072 17066
rect 46020 17002 46072 17008
rect 45008 16652 45060 16658
rect 45008 16594 45060 16600
rect 45560 16652 45612 16658
rect 45560 16594 45612 16600
rect 45376 16584 45428 16590
rect 45376 16526 45428 16532
rect 44916 16516 44968 16522
rect 44916 16458 44968 16464
rect 45388 15638 45416 16526
rect 45572 16250 45600 16594
rect 46032 16590 46060 17002
rect 46020 16584 46072 16590
rect 46020 16526 46072 16532
rect 45560 16244 45612 16250
rect 45560 16186 45612 16192
rect 45376 15632 45428 15638
rect 45376 15574 45428 15580
rect 44088 15020 44140 15026
rect 44088 14962 44140 14968
rect 44100 13530 44128 14962
rect 45192 14816 45244 14822
rect 45192 14758 45244 14764
rect 45468 14816 45520 14822
rect 45468 14758 45520 14764
rect 45204 14414 45232 14758
rect 45480 14414 45508 14758
rect 45192 14408 45244 14414
rect 45192 14350 45244 14356
rect 45468 14408 45520 14414
rect 45468 14350 45520 14356
rect 44180 14272 44232 14278
rect 44180 14214 44232 14220
rect 44088 13524 44140 13530
rect 44088 13466 44140 13472
rect 44192 13326 44220 14214
rect 45204 14006 45232 14350
rect 45192 14000 45244 14006
rect 45192 13942 45244 13948
rect 45480 13802 45508 14350
rect 44364 13796 44416 13802
rect 44364 13738 44416 13744
rect 45468 13796 45520 13802
rect 45468 13738 45520 13744
rect 44180 13320 44232 13326
rect 44180 13262 44232 13268
rect 44376 12918 44404 13738
rect 44364 12912 44416 12918
rect 44364 12854 44416 12860
rect 43824 12406 43944 12434
rect 43720 12232 43772 12238
rect 43720 12174 43772 12180
rect 42708 11552 42760 11558
rect 42708 11494 42760 11500
rect 42720 11150 42748 11494
rect 43824 11354 43852 12406
rect 44272 12232 44324 12238
rect 44272 12174 44324 12180
rect 45468 12232 45520 12238
rect 45468 12174 45520 12180
rect 43904 11688 43956 11694
rect 43904 11630 43956 11636
rect 43812 11348 43864 11354
rect 43812 11290 43864 11296
rect 43916 11218 43944 11630
rect 44180 11348 44232 11354
rect 44180 11290 44232 11296
rect 43904 11212 43956 11218
rect 43904 11154 43956 11160
rect 42708 11144 42760 11150
rect 42708 11086 42760 11092
rect 42720 10810 42748 11086
rect 42708 10804 42760 10810
rect 42708 10746 42760 10752
rect 43628 10600 43680 10606
rect 43628 10542 43680 10548
rect 43536 10532 43588 10538
rect 43536 10474 43588 10480
rect 42616 10464 42668 10470
rect 42616 10406 42668 10412
rect 41420 10124 41472 10130
rect 41420 10066 41472 10072
rect 40960 9376 41012 9382
rect 40960 9318 41012 9324
rect 40972 8906 41000 9318
rect 40960 8900 41012 8906
rect 40960 8842 41012 8848
rect 41696 8832 41748 8838
rect 41696 8774 41748 8780
rect 41708 8566 41736 8774
rect 41696 8560 41748 8566
rect 41696 8502 41748 8508
rect 40960 8424 41012 8430
rect 40960 8366 41012 8372
rect 40972 8090 41000 8366
rect 41144 8356 41196 8362
rect 41144 8298 41196 8304
rect 41236 8356 41288 8362
rect 41236 8298 41288 8304
rect 40960 8084 41012 8090
rect 40960 8026 41012 8032
rect 40868 8016 40920 8022
rect 40868 7958 40920 7964
rect 40880 7410 40908 7958
rect 40868 7404 40920 7410
rect 40972 7392 41000 8026
rect 41156 7954 41184 8298
rect 41144 7948 41196 7954
rect 41144 7890 41196 7896
rect 41156 7546 41184 7890
rect 41248 7750 41276 8298
rect 41708 8090 41736 8502
rect 41788 8424 41840 8430
rect 41788 8366 41840 8372
rect 41696 8084 41748 8090
rect 41696 8026 41748 8032
rect 41604 7880 41656 7886
rect 41604 7822 41656 7828
rect 41236 7744 41288 7750
rect 41236 7686 41288 7692
rect 41144 7540 41196 7546
rect 41144 7482 41196 7488
rect 41248 7410 41276 7686
rect 41616 7546 41644 7822
rect 41604 7540 41656 7546
rect 41604 7482 41656 7488
rect 41052 7404 41104 7410
rect 40972 7364 41052 7392
rect 40868 7346 40920 7352
rect 41052 7346 41104 7352
rect 41236 7404 41288 7410
rect 41708 7392 41736 8026
rect 41800 7546 41828 8366
rect 42628 7585 42656 10406
rect 43548 10130 43576 10474
rect 43536 10124 43588 10130
rect 43536 10066 43588 10072
rect 42984 9988 43036 9994
rect 42984 9930 43036 9936
rect 42996 9722 43024 9930
rect 43640 9926 43668 10542
rect 43628 9920 43680 9926
rect 43628 9862 43680 9868
rect 42984 9716 43036 9722
rect 42984 9658 43036 9664
rect 43640 9518 43668 9862
rect 44192 9654 44220 11290
rect 44284 11150 44312 12174
rect 45100 12096 45152 12102
rect 45100 12038 45152 12044
rect 44272 11144 44324 11150
rect 44272 11086 44324 11092
rect 45112 10742 45140 12038
rect 45480 11762 45508 12174
rect 46860 12102 46888 21490
rect 48700 14550 48728 23666
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 48688 14544 48740 14550
rect 48688 14486 48740 14492
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 48964 12912 49016 12918
rect 48964 12854 49016 12860
rect 48596 12844 48648 12850
rect 48596 12786 48648 12792
rect 47952 12368 48004 12374
rect 47952 12310 48004 12316
rect 45560 12096 45612 12102
rect 45560 12038 45612 12044
rect 46848 12096 46900 12102
rect 46848 12038 46900 12044
rect 45572 11898 45600 12038
rect 45560 11892 45612 11898
rect 45560 11834 45612 11840
rect 47964 11762 47992 12310
rect 48044 12232 48096 12238
rect 48044 12174 48096 12180
rect 48056 11898 48084 12174
rect 48136 12164 48188 12170
rect 48136 12106 48188 12112
rect 48044 11892 48096 11898
rect 48044 11834 48096 11840
rect 45468 11756 45520 11762
rect 45468 11698 45520 11704
rect 47952 11756 48004 11762
rect 47952 11698 48004 11704
rect 45100 10736 45152 10742
rect 45100 10678 45152 10684
rect 45480 10062 45508 11698
rect 46756 11620 46808 11626
rect 46756 11562 46808 11568
rect 46768 11354 46796 11562
rect 46940 11552 46992 11558
rect 46940 11494 46992 11500
rect 46756 11348 46808 11354
rect 46756 11290 46808 11296
rect 46952 10810 46980 11494
rect 47400 11144 47452 11150
rect 47400 11086 47452 11092
rect 47032 11076 47084 11082
rect 47032 11018 47084 11024
rect 47044 10810 47072 11018
rect 47412 10810 47440 11086
rect 46940 10804 46992 10810
rect 46940 10746 46992 10752
rect 47032 10804 47084 10810
rect 47032 10746 47084 10752
rect 47400 10804 47452 10810
rect 47400 10746 47452 10752
rect 46848 10668 46900 10674
rect 46848 10610 46900 10616
rect 46756 10600 46808 10606
rect 46756 10542 46808 10548
rect 46768 10130 46796 10542
rect 46860 10266 46888 10610
rect 46848 10260 46900 10266
rect 46848 10202 46900 10208
rect 46756 10124 46808 10130
rect 46756 10066 46808 10072
rect 45468 10056 45520 10062
rect 45468 9998 45520 10004
rect 45008 9920 45060 9926
rect 45008 9862 45060 9868
rect 44180 9648 44232 9654
rect 44180 9590 44232 9596
rect 43628 9512 43680 9518
rect 43628 9454 43680 9460
rect 43640 8650 43668 9454
rect 44192 8974 44220 9590
rect 45020 9586 45048 9862
rect 45008 9580 45060 9586
rect 45008 9522 45060 9528
rect 46768 9518 46796 10066
rect 47044 10062 47072 10746
rect 47032 10056 47084 10062
rect 47032 9998 47084 10004
rect 47584 9920 47636 9926
rect 47584 9862 47636 9868
rect 47596 9518 47624 9862
rect 46756 9512 46808 9518
rect 46756 9454 46808 9460
rect 47584 9512 47636 9518
rect 47584 9454 47636 9460
rect 47768 9376 47820 9382
rect 47768 9318 47820 9324
rect 46940 9172 46992 9178
rect 46940 9114 46992 9120
rect 44180 8968 44232 8974
rect 44180 8910 44232 8916
rect 44272 8832 44324 8838
rect 44272 8774 44324 8780
rect 43640 8634 43760 8650
rect 43640 8628 43772 8634
rect 43640 8622 43720 8628
rect 43720 8570 43772 8576
rect 43260 8492 43312 8498
rect 43260 8434 43312 8440
rect 43272 7886 43300 8434
rect 43260 7880 43312 7886
rect 43260 7822 43312 7828
rect 43076 7812 43128 7818
rect 43076 7754 43128 7760
rect 42614 7576 42670 7585
rect 41788 7540 41840 7546
rect 42614 7511 42670 7520
rect 41788 7482 41840 7488
rect 43088 7410 43116 7754
rect 43272 7410 43300 7822
rect 41788 7404 41840 7410
rect 41708 7364 41788 7392
rect 41236 7346 41288 7352
rect 41788 7346 41840 7352
rect 43076 7404 43128 7410
rect 43076 7346 43128 7352
rect 43260 7404 43312 7410
rect 43260 7346 43312 7352
rect 41236 7268 41288 7274
rect 41236 7210 41288 7216
rect 41144 6860 41196 6866
rect 41144 6802 41196 6808
rect 40684 6724 40736 6730
rect 40684 6666 40736 6672
rect 40960 6316 41012 6322
rect 40960 6258 41012 6264
rect 40590 5264 40646 5273
rect 40590 5199 40646 5208
rect 40604 4146 40632 5199
rect 40972 4826 41000 6258
rect 41156 5778 41184 6802
rect 41248 6322 41276 7210
rect 41236 6316 41288 6322
rect 41236 6258 41288 6264
rect 41800 6118 41828 7346
rect 43732 7342 43760 8570
rect 44284 8566 44312 8774
rect 44272 8560 44324 8566
rect 44272 8502 44324 8508
rect 46952 8022 46980 9114
rect 47780 8906 47808 9318
rect 47964 8974 47992 11698
rect 48056 11286 48084 11834
rect 48148 11830 48176 12106
rect 48320 12096 48372 12102
rect 48320 12038 48372 12044
rect 48136 11824 48188 11830
rect 48136 11766 48188 11772
rect 48148 11354 48176 11766
rect 48136 11348 48188 11354
rect 48136 11290 48188 11296
rect 48044 11280 48096 11286
rect 48044 11222 48096 11228
rect 48332 11218 48360 12038
rect 48504 11756 48556 11762
rect 48504 11698 48556 11704
rect 48320 11212 48372 11218
rect 48320 11154 48372 11160
rect 48332 11098 48360 11154
rect 48516 11150 48544 11698
rect 48608 11626 48636 12786
rect 48872 12436 48924 12442
rect 48872 12378 48924 12384
rect 48596 11620 48648 11626
rect 48596 11562 48648 11568
rect 48884 11558 48912 12378
rect 48976 12374 49004 12854
rect 49424 12776 49476 12782
rect 49424 12718 49476 12724
rect 49056 12640 49108 12646
rect 49056 12582 49108 12588
rect 48964 12368 49016 12374
rect 48964 12310 49016 12316
rect 48872 11552 48924 11558
rect 48872 11494 48924 11500
rect 48148 11070 48360 11098
rect 48504 11144 48556 11150
rect 48504 11086 48556 11092
rect 47952 8968 48004 8974
rect 47952 8910 48004 8916
rect 47768 8900 47820 8906
rect 47768 8842 47820 8848
rect 46940 8016 46992 8022
rect 46940 7958 46992 7964
rect 45008 7880 45060 7886
rect 45008 7822 45060 7828
rect 45560 7880 45612 7886
rect 45560 7822 45612 7828
rect 43996 7744 44048 7750
rect 43996 7686 44048 7692
rect 44088 7744 44140 7750
rect 44088 7686 44140 7692
rect 44008 7478 44036 7686
rect 44100 7546 44128 7686
rect 44088 7540 44140 7546
rect 44088 7482 44140 7488
rect 43996 7472 44048 7478
rect 43996 7414 44048 7420
rect 43720 7336 43772 7342
rect 43720 7278 43772 7284
rect 41880 6792 41932 6798
rect 41880 6734 41932 6740
rect 41892 6458 41920 6734
rect 43352 6656 43404 6662
rect 43352 6598 43404 6604
rect 43364 6458 43392 6598
rect 41880 6452 41932 6458
rect 41880 6394 41932 6400
rect 43352 6452 43404 6458
rect 43352 6394 43404 6400
rect 43732 6254 43760 7278
rect 43996 7200 44048 7206
rect 43996 7142 44048 7148
rect 44456 7200 44508 7206
rect 44456 7142 44508 7148
rect 44008 6798 44036 7142
rect 43996 6792 44048 6798
rect 43996 6734 44048 6740
rect 44272 6792 44324 6798
rect 44272 6734 44324 6740
rect 44180 6656 44232 6662
rect 44180 6598 44232 6604
rect 44192 6390 44220 6598
rect 44284 6458 44312 6734
rect 44272 6452 44324 6458
rect 44272 6394 44324 6400
rect 44180 6384 44232 6390
rect 44180 6326 44232 6332
rect 43720 6248 43772 6254
rect 43720 6190 43772 6196
rect 41788 6112 41840 6118
rect 41788 6054 41840 6060
rect 41144 5772 41196 5778
rect 41144 5714 41196 5720
rect 40960 4820 41012 4826
rect 40960 4762 41012 4768
rect 41156 4690 41184 5714
rect 41328 5364 41380 5370
rect 41328 5306 41380 5312
rect 41340 5250 41368 5306
rect 41248 5222 41368 5250
rect 42432 5296 42484 5302
rect 42432 5238 42484 5244
rect 41248 4758 41276 5222
rect 41328 5160 41380 5166
rect 41328 5102 41380 5108
rect 41236 4752 41288 4758
rect 41236 4694 41288 4700
rect 41144 4684 41196 4690
rect 41144 4626 41196 4632
rect 40866 4584 40922 4593
rect 40866 4519 40868 4528
rect 40920 4519 40922 4528
rect 40868 4490 40920 4496
rect 40592 4140 40644 4146
rect 40592 4082 40644 4088
rect 40604 4049 40632 4082
rect 40590 4040 40646 4049
rect 40408 4004 40460 4010
rect 40590 3975 40646 3984
rect 40408 3946 40460 3952
rect 40592 3936 40644 3942
rect 40592 3878 40644 3884
rect 40604 3466 40632 3878
rect 40592 3460 40644 3466
rect 40592 3402 40644 3408
rect 41144 3392 41196 3398
rect 41144 3334 41196 3340
rect 41156 3126 41184 3334
rect 41144 3120 41196 3126
rect 41144 3062 41196 3068
rect 41052 2916 41104 2922
rect 41052 2858 41104 2864
rect 40408 2576 40460 2582
rect 40408 2518 40460 2524
rect 39948 2508 40000 2514
rect 39948 2450 40000 2456
rect 40224 2440 40276 2446
rect 40224 2382 40276 2388
rect 39856 2304 39908 2310
rect 39856 2246 39908 2252
rect 40132 2304 40184 2310
rect 40132 2246 40184 2252
rect 39868 800 39896 2246
rect 40144 800 40172 2246
rect 40236 2106 40264 2382
rect 40224 2100 40276 2106
rect 40224 2042 40276 2048
rect 40420 800 40448 2518
rect 40960 2440 41012 2446
rect 40960 2382 41012 2388
rect 40868 2304 40920 2310
rect 40696 2264 40868 2292
rect 40696 800 40724 2264
rect 40868 2246 40920 2252
rect 40972 1970 41000 2382
rect 40960 1964 41012 1970
rect 40960 1906 41012 1912
rect 41064 1442 41092 2858
rect 41248 2774 41276 4694
rect 41340 4690 41368 5102
rect 41788 5024 41840 5030
rect 41788 4966 41840 4972
rect 41328 4684 41380 4690
rect 41328 4626 41380 4632
rect 41800 4078 41828 4966
rect 42154 4584 42210 4593
rect 42154 4519 42210 4528
rect 41878 4312 41934 4321
rect 41878 4247 41934 4256
rect 41788 4072 41840 4078
rect 41788 4014 41840 4020
rect 41788 3936 41840 3942
rect 41788 3878 41840 3884
rect 41604 3392 41656 3398
rect 41524 3352 41604 3380
rect 41524 3058 41552 3352
rect 41604 3334 41656 3340
rect 41512 3052 41564 3058
rect 41512 2994 41564 3000
rect 41248 2746 41368 2774
rect 41340 2038 41368 2746
rect 41604 2576 41656 2582
rect 41604 2518 41656 2524
rect 41328 2032 41380 2038
rect 41328 1974 41380 1980
rect 41236 1828 41288 1834
rect 41236 1770 41288 1776
rect 40972 1414 41092 1442
rect 40972 800 41000 1414
rect 41248 800 41276 1770
rect 41616 1170 41644 2518
rect 41524 1142 41644 1170
rect 41524 800 41552 1142
rect 41800 800 41828 3878
rect 41892 3058 41920 4247
rect 41972 3596 42024 3602
rect 41972 3538 42024 3544
rect 41880 3052 41932 3058
rect 41880 2994 41932 3000
rect 41984 2990 42012 3538
rect 42064 3120 42116 3126
rect 42064 3062 42116 3068
rect 41972 2984 42024 2990
rect 41972 2926 42024 2932
rect 42076 800 42104 3062
rect 42168 2446 42196 4519
rect 42340 4480 42392 4486
rect 42340 4422 42392 4428
rect 42248 4208 42300 4214
rect 42248 4150 42300 4156
rect 42260 2854 42288 4150
rect 42352 3398 42380 4422
rect 42444 4146 42472 5238
rect 42800 5228 42852 5234
rect 42800 5170 42852 5176
rect 42812 4622 42840 5170
rect 43352 5160 43404 5166
rect 43352 5102 43404 5108
rect 43364 4622 43392 5102
rect 42800 4616 42852 4622
rect 42800 4558 42852 4564
rect 42984 4616 43036 4622
rect 42984 4558 43036 4564
rect 43352 4616 43404 4622
rect 43352 4558 43404 4564
rect 42524 4548 42576 4554
rect 42524 4490 42576 4496
rect 42616 4548 42668 4554
rect 42616 4490 42668 4496
rect 42432 4140 42484 4146
rect 42432 4082 42484 4088
rect 42432 4004 42484 4010
rect 42432 3946 42484 3952
rect 42444 3602 42472 3946
rect 42536 3602 42564 4490
rect 42628 4282 42656 4490
rect 42800 4480 42852 4486
rect 42800 4422 42852 4428
rect 42616 4276 42668 4282
rect 42616 4218 42668 4224
rect 42616 3664 42668 3670
rect 42616 3606 42668 3612
rect 42432 3596 42484 3602
rect 42432 3538 42484 3544
rect 42524 3596 42576 3602
rect 42524 3538 42576 3544
rect 42536 3398 42564 3538
rect 42340 3392 42392 3398
rect 42524 3392 42576 3398
rect 42392 3352 42472 3380
rect 42340 3334 42392 3340
rect 42340 2984 42392 2990
rect 42340 2926 42392 2932
rect 42248 2848 42300 2854
rect 42248 2790 42300 2796
rect 42156 2440 42208 2446
rect 42156 2382 42208 2388
rect 42352 800 42380 2926
rect 42444 2417 42472 3352
rect 42524 3334 42576 3340
rect 42524 2848 42576 2854
rect 42524 2790 42576 2796
rect 42536 2446 42564 2790
rect 42524 2440 42576 2446
rect 42430 2408 42486 2417
rect 42524 2382 42576 2388
rect 42430 2343 42486 2352
rect 42628 800 42656 3606
rect 42812 3534 42840 4422
rect 42996 3738 43024 4558
rect 43364 3913 43392 4558
rect 43536 4480 43588 4486
rect 43536 4422 43588 4428
rect 43444 3936 43496 3942
rect 43350 3904 43406 3913
rect 43444 3878 43496 3884
rect 43350 3839 43406 3848
rect 42984 3732 43036 3738
rect 42984 3674 43036 3680
rect 43456 3602 43484 3878
rect 43444 3596 43496 3602
rect 43444 3538 43496 3544
rect 42800 3528 42852 3534
rect 42800 3470 42852 3476
rect 42708 3392 42760 3398
rect 42708 3334 42760 3340
rect 43444 3392 43496 3398
rect 43444 3334 43496 3340
rect 42720 3126 42748 3334
rect 42708 3120 42760 3126
rect 42708 3062 42760 3068
rect 43168 2916 43220 2922
rect 43168 2858 43220 2864
rect 42800 2848 42852 2854
rect 42800 2790 42852 2796
rect 42812 2514 42840 2790
rect 42800 2508 42852 2514
rect 42800 2450 42852 2456
rect 42892 2508 42944 2514
rect 42892 2450 42944 2456
rect 42798 2408 42854 2417
rect 42798 2343 42800 2352
rect 42852 2343 42854 2352
rect 42800 2314 42852 2320
rect 42708 2304 42760 2310
rect 42708 2246 42760 2252
rect 42720 1834 42748 2246
rect 42708 1828 42760 1834
rect 42708 1770 42760 1776
rect 42904 800 42932 2450
rect 43180 800 43208 2858
rect 43456 800 43484 3334
rect 43548 3126 43576 4422
rect 43626 3496 43682 3505
rect 43626 3431 43682 3440
rect 43536 3120 43588 3126
rect 43536 3062 43588 3068
rect 43536 2848 43588 2854
rect 43640 2836 43668 3431
rect 43732 3194 43760 6190
rect 44272 4616 44324 4622
rect 44272 4558 44324 4564
rect 44180 4480 44232 4486
rect 44180 4422 44232 4428
rect 44192 4214 44220 4422
rect 44180 4208 44232 4214
rect 44180 4150 44232 4156
rect 44284 4049 44312 4558
rect 44270 4040 44326 4049
rect 44270 3975 44326 3984
rect 43812 3732 43864 3738
rect 43812 3674 43864 3680
rect 43720 3188 43772 3194
rect 43720 3130 43772 3136
rect 43588 2808 43668 2836
rect 43536 2790 43588 2796
rect 43824 2774 43852 3674
rect 44272 2984 44324 2990
rect 43994 2952 44050 2961
rect 44272 2926 44324 2932
rect 43994 2887 44050 2896
rect 43732 2746 43852 2774
rect 43732 800 43760 2746
rect 43904 2440 43956 2446
rect 43904 2382 43956 2388
rect 43916 2038 43944 2382
rect 43904 2032 43956 2038
rect 43904 1974 43956 1980
rect 44008 800 44036 2887
rect 44284 2582 44312 2926
rect 44468 2774 44496 7142
rect 45020 6866 45048 7822
rect 45100 7744 45152 7750
rect 45100 7686 45152 7692
rect 45112 7410 45140 7686
rect 45100 7404 45152 7410
rect 45100 7346 45152 7352
rect 45192 6996 45244 7002
rect 45192 6938 45244 6944
rect 45008 6860 45060 6866
rect 45008 6802 45060 6808
rect 45204 6798 45232 6938
rect 45572 6934 45600 7822
rect 45560 6928 45612 6934
rect 45560 6870 45612 6876
rect 45192 6792 45244 6798
rect 45192 6734 45244 6740
rect 47492 6724 47544 6730
rect 47492 6666 47544 6672
rect 45744 6656 45796 6662
rect 45744 6598 45796 6604
rect 45756 6390 45784 6598
rect 45744 6384 45796 6390
rect 45744 6326 45796 6332
rect 47124 6248 47176 6254
rect 47124 6190 47176 6196
rect 46940 6112 46992 6118
rect 46940 6054 46992 6060
rect 46296 5908 46348 5914
rect 46296 5850 46348 5856
rect 46308 5166 46336 5850
rect 46952 5760 46980 6054
rect 46860 5732 46980 5760
rect 46480 5704 46532 5710
rect 46480 5646 46532 5652
rect 46296 5160 46348 5166
rect 46296 5102 46348 5108
rect 45652 5024 45704 5030
rect 45652 4966 45704 4972
rect 45928 5024 45980 5030
rect 45928 4966 45980 4972
rect 44824 4684 44876 4690
rect 44824 4626 44876 4632
rect 44548 3596 44600 3602
rect 44548 3538 44600 3544
rect 44376 2746 44496 2774
rect 44272 2576 44324 2582
rect 44272 2518 44324 2524
rect 44376 2106 44404 2746
rect 44364 2100 44416 2106
rect 44364 2042 44416 2048
rect 44272 2032 44324 2038
rect 44272 1974 44324 1980
rect 44284 800 44312 1974
rect 44560 800 44588 3538
rect 44836 800 44864 4626
rect 45100 4616 45152 4622
rect 45100 4558 45152 4564
rect 45376 4616 45428 4622
rect 45376 4558 45428 4564
rect 45008 4480 45060 4486
rect 45008 4422 45060 4428
rect 45020 4214 45048 4422
rect 45008 4208 45060 4214
rect 45008 4150 45060 4156
rect 45112 3738 45140 4558
rect 45192 4072 45244 4078
rect 45192 4014 45244 4020
rect 45100 3732 45152 3738
rect 45100 3674 45152 3680
rect 45204 3194 45232 4014
rect 45284 3392 45336 3398
rect 45284 3334 45336 3340
rect 45192 3188 45244 3194
rect 45192 3130 45244 3136
rect 45296 2922 45324 3334
rect 45284 2916 45336 2922
rect 45284 2858 45336 2864
rect 45282 2816 45338 2825
rect 45282 2751 45338 2760
rect 45008 2304 45060 2310
rect 45008 2246 45060 2252
rect 45020 800 45048 2246
rect 45100 1896 45152 1902
rect 45100 1838 45152 1844
rect 45112 800 45140 1838
rect 45296 800 45324 2751
rect 45388 800 45416 4558
rect 45560 3936 45612 3942
rect 45560 3878 45612 3884
rect 45572 3602 45600 3878
rect 45560 3596 45612 3602
rect 45560 3538 45612 3544
rect 45560 1828 45612 1834
rect 45560 1770 45612 1776
rect 45572 800 45600 1770
rect 45664 800 45692 4966
rect 45836 4140 45888 4146
rect 45836 4082 45888 4088
rect 45848 800 45876 4082
rect 45940 800 45968 4966
rect 46204 4684 46256 4690
rect 46204 4626 46256 4632
rect 46112 4004 46164 4010
rect 46112 3946 46164 3952
rect 46020 3664 46072 3670
rect 46020 3606 46072 3612
rect 46032 2854 46060 3606
rect 46020 2848 46072 2854
rect 46020 2790 46072 2796
rect 46124 800 46152 3946
rect 46216 800 46244 4626
rect 46308 4078 46336 5102
rect 46388 4276 46440 4282
rect 46388 4218 46440 4224
rect 46296 4072 46348 4078
rect 46296 4014 46348 4020
rect 46308 2582 46336 4014
rect 46400 3602 46428 4218
rect 46388 3596 46440 3602
rect 46388 3538 46440 3544
rect 46388 3460 46440 3466
rect 46388 3402 46440 3408
rect 46296 2576 46348 2582
rect 46296 2518 46348 2524
rect 46400 800 46428 3402
rect 46492 800 46520 5646
rect 46572 5568 46624 5574
rect 46572 5510 46624 5516
rect 46584 4146 46612 5510
rect 46860 5098 46888 5732
rect 47136 5386 47164 6190
rect 46952 5358 47164 5386
rect 46848 5092 46900 5098
rect 46848 5034 46900 5040
rect 46756 5024 46808 5030
rect 46756 4966 46808 4972
rect 46572 4140 46624 4146
rect 46572 4082 46624 4088
rect 46584 2310 46612 4082
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 46676 2582 46704 3878
rect 46664 2576 46716 2582
rect 46664 2518 46716 2524
rect 46664 2372 46716 2378
rect 46664 2314 46716 2320
rect 46572 2304 46624 2310
rect 46572 2246 46624 2252
rect 46676 2106 46704 2314
rect 46664 2100 46716 2106
rect 46664 2042 46716 2048
rect 46768 800 46796 4966
rect 46860 3942 46888 5034
rect 46952 4622 46980 5358
rect 47308 5092 47360 5098
rect 47308 5034 47360 5040
rect 47216 4752 47268 4758
rect 47216 4694 47268 4700
rect 46940 4616 46992 4622
rect 46940 4558 46992 4564
rect 46952 4010 46980 4558
rect 47032 4480 47084 4486
rect 47032 4422 47084 4428
rect 46940 4004 46992 4010
rect 46940 3946 46992 3952
rect 46848 3936 46900 3942
rect 46848 3878 46900 3884
rect 47044 3534 47072 4422
rect 47124 3936 47176 3942
rect 47124 3878 47176 3884
rect 47136 3602 47164 3878
rect 47124 3596 47176 3602
rect 47124 3538 47176 3544
rect 47032 3528 47084 3534
rect 47032 3470 47084 3476
rect 47228 2774 47256 4694
rect 47044 2746 47256 2774
rect 47044 800 47072 2746
rect 47216 1760 47268 1766
rect 47216 1702 47268 1708
rect 47228 800 47256 1702
rect 47320 800 47348 5034
rect 47400 3528 47452 3534
rect 47400 3470 47452 3476
rect 47412 1902 47440 3470
rect 47504 2514 47532 6666
rect 47676 4684 47728 4690
rect 47676 4626 47728 4632
rect 47582 2952 47638 2961
rect 47582 2887 47584 2896
rect 47636 2887 47638 2896
rect 47584 2858 47636 2864
rect 47492 2508 47544 2514
rect 47492 2450 47544 2456
rect 47400 1896 47452 1902
rect 47400 1838 47452 1844
rect 47688 1442 47716 4626
rect 47780 3738 47808 8842
rect 47860 7200 47912 7206
rect 47860 7142 47912 7148
rect 47768 3732 47820 3738
rect 47768 3674 47820 3680
rect 47872 2378 47900 7142
rect 48148 5370 48176 11070
rect 48596 10668 48648 10674
rect 48596 10610 48648 10616
rect 48412 10464 48464 10470
rect 48412 10406 48464 10412
rect 48228 10056 48280 10062
rect 48280 10004 48360 10010
rect 48228 9998 48360 10004
rect 48240 9982 48360 9998
rect 48332 8498 48360 9982
rect 48424 9450 48452 10406
rect 48608 10266 48636 10610
rect 48504 10260 48556 10266
rect 48504 10202 48556 10208
rect 48596 10260 48648 10266
rect 48596 10202 48648 10208
rect 48516 10146 48544 10202
rect 48884 10146 48912 11494
rect 48976 11286 49004 12310
rect 49068 12170 49096 12582
rect 49056 12164 49108 12170
rect 49056 12106 49108 12112
rect 49240 11892 49292 11898
rect 49240 11834 49292 11840
rect 49252 11762 49280 11834
rect 49436 11762 49464 12718
rect 50160 12640 50212 12646
rect 50160 12582 50212 12588
rect 49700 11892 49752 11898
rect 49700 11834 49752 11840
rect 49148 11756 49200 11762
rect 49148 11698 49200 11704
rect 49240 11756 49292 11762
rect 49240 11698 49292 11704
rect 49424 11756 49476 11762
rect 49424 11698 49476 11704
rect 48964 11280 49016 11286
rect 48964 11222 49016 11228
rect 48976 11150 49004 11222
rect 49160 11150 49188 11698
rect 48964 11144 49016 11150
rect 48964 11086 49016 11092
rect 49148 11144 49200 11150
rect 49148 11086 49200 11092
rect 49436 11014 49464 11698
rect 49424 11008 49476 11014
rect 49424 10950 49476 10956
rect 49436 10810 49464 10950
rect 49424 10804 49476 10810
rect 49424 10746 49476 10752
rect 49436 10538 49464 10746
rect 49424 10532 49476 10538
rect 49424 10474 49476 10480
rect 49608 10532 49660 10538
rect 49608 10474 49660 10480
rect 48516 10118 48912 10146
rect 49148 10192 49200 10198
rect 49148 10134 49200 10140
rect 49516 10192 49568 10198
rect 49516 10134 49568 10140
rect 48596 9988 48648 9994
rect 48596 9930 48648 9936
rect 48608 9586 48636 9930
rect 48596 9580 48648 9586
rect 48596 9522 48648 9528
rect 48412 9444 48464 9450
rect 48412 9386 48464 9392
rect 48504 8832 48556 8838
rect 48504 8774 48556 8780
rect 48320 8492 48372 8498
rect 48320 8434 48372 8440
rect 48332 7886 48360 8434
rect 48320 7880 48372 7886
rect 48320 7822 48372 7828
rect 48516 7410 48544 8774
rect 48608 8430 48636 9522
rect 48780 9376 48832 9382
rect 48780 9318 48832 9324
rect 48792 8974 48820 9318
rect 48884 9178 48912 10118
rect 49160 9926 49188 10134
rect 49332 10124 49384 10130
rect 49332 10066 49384 10072
rect 49240 10056 49292 10062
rect 49240 9998 49292 10004
rect 49148 9920 49200 9926
rect 49148 9862 49200 9868
rect 49160 9586 49188 9862
rect 49252 9722 49280 9998
rect 49240 9716 49292 9722
rect 49240 9658 49292 9664
rect 49148 9580 49200 9586
rect 49148 9522 49200 9528
rect 49344 9178 49372 10066
rect 49424 9648 49476 9654
rect 49424 9590 49476 9596
rect 48872 9172 48924 9178
rect 48872 9114 48924 9120
rect 49332 9172 49384 9178
rect 49332 9114 49384 9120
rect 48780 8968 48832 8974
rect 48780 8910 48832 8916
rect 48884 8566 48912 9114
rect 49436 9110 49464 9590
rect 49424 9104 49476 9110
rect 49424 9046 49476 9052
rect 48964 9036 49016 9042
rect 48964 8978 49016 8984
rect 48872 8560 48924 8566
rect 48872 8502 48924 8508
rect 48976 8498 49004 8978
rect 49332 8560 49384 8566
rect 49332 8502 49384 8508
rect 48964 8492 49016 8498
rect 48964 8434 49016 8440
rect 48596 8424 48648 8430
rect 48596 8366 48648 8372
rect 49344 8294 49372 8502
rect 49436 8498 49464 9046
rect 49528 8906 49556 10134
rect 49620 8974 49648 10474
rect 49712 9586 49740 11834
rect 49884 11756 49936 11762
rect 49884 11698 49936 11704
rect 49896 11354 49924 11698
rect 49884 11348 49936 11354
rect 49884 11290 49936 11296
rect 49976 11144 50028 11150
rect 49976 11086 50028 11092
rect 49792 10600 49844 10606
rect 49792 10542 49844 10548
rect 49804 10266 49832 10542
rect 49792 10260 49844 10266
rect 49792 10202 49844 10208
rect 49988 10130 50016 11086
rect 50172 11082 50200 12582
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 50620 11280 50672 11286
rect 50620 11222 50672 11228
rect 50160 11076 50212 11082
rect 50160 11018 50212 11024
rect 50068 10736 50120 10742
rect 50068 10678 50120 10684
rect 49792 10124 49844 10130
rect 49792 10066 49844 10072
rect 49976 10124 50028 10130
rect 49976 10066 50028 10072
rect 49700 9580 49752 9586
rect 49700 9522 49752 9528
rect 49712 9110 49740 9522
rect 49700 9104 49752 9110
rect 49700 9046 49752 9052
rect 49608 8968 49660 8974
rect 49608 8910 49660 8916
rect 49516 8900 49568 8906
rect 49516 8842 49568 8848
rect 49712 8498 49740 9046
rect 49424 8492 49476 8498
rect 49424 8434 49476 8440
rect 49700 8492 49752 8498
rect 49700 8434 49752 8440
rect 48596 8288 48648 8294
rect 48596 8230 48648 8236
rect 49332 8288 49384 8294
rect 49332 8230 49384 8236
rect 48608 7886 48636 8230
rect 49436 7970 49464 8434
rect 49804 8378 49832 10066
rect 49882 10024 49938 10033
rect 49882 9959 49938 9968
rect 49976 9988 50028 9994
rect 49896 9654 49924 9959
rect 49976 9930 50028 9936
rect 49988 9722 50016 9930
rect 49976 9716 50028 9722
rect 49976 9658 50028 9664
rect 49884 9648 49936 9654
rect 49884 9590 49936 9596
rect 49884 9512 49936 9518
rect 49884 9454 49936 9460
rect 49608 8356 49660 8362
rect 49608 8298 49660 8304
rect 49712 8350 49832 8378
rect 49344 7942 49464 7970
rect 49344 7886 49372 7942
rect 48596 7880 48648 7886
rect 48596 7822 48648 7828
rect 49332 7880 49384 7886
rect 49332 7822 49384 7828
rect 49620 7834 49648 8298
rect 49712 7954 49740 8350
rect 49700 7948 49752 7954
rect 49700 7890 49752 7896
rect 49620 7806 49832 7834
rect 48596 7744 48648 7750
rect 48596 7686 48648 7692
rect 49700 7744 49752 7750
rect 49700 7686 49752 7692
rect 48504 7404 48556 7410
rect 48504 7346 48556 7352
rect 48320 7200 48372 7206
rect 48320 7142 48372 7148
rect 48332 6798 48360 7142
rect 48608 6866 48636 7686
rect 48412 6860 48464 6866
rect 48412 6802 48464 6808
rect 48596 6860 48648 6866
rect 48596 6802 48648 6808
rect 48320 6792 48372 6798
rect 48320 6734 48372 6740
rect 48332 6322 48360 6734
rect 48320 6316 48372 6322
rect 48320 6258 48372 6264
rect 48424 5710 48452 6802
rect 49424 6792 49476 6798
rect 49424 6734 49476 6740
rect 48504 6656 48556 6662
rect 48504 6598 48556 6604
rect 48412 5704 48464 5710
rect 48412 5646 48464 5652
rect 48424 5574 48452 5646
rect 48412 5568 48464 5574
rect 48412 5510 48464 5516
rect 48136 5364 48188 5370
rect 48136 5306 48188 5312
rect 48136 4820 48188 4826
rect 48136 4762 48188 4768
rect 48044 4616 48096 4622
rect 48044 4558 48096 4564
rect 47952 3596 48004 3602
rect 47952 3538 48004 3544
rect 47860 2372 47912 2378
rect 47860 2314 47912 2320
rect 47872 1766 47900 2314
rect 47860 1760 47912 1766
rect 47860 1702 47912 1708
rect 47964 1442 47992 3538
rect 48056 3466 48084 4558
rect 48044 3460 48096 3466
rect 48044 3402 48096 3408
rect 47596 1414 47716 1442
rect 47872 1414 47992 1442
rect 47596 800 47624 1414
rect 47872 800 47900 1414
rect 48148 800 48176 4762
rect 48320 4616 48372 4622
rect 48240 4564 48320 4570
rect 48240 4558 48372 4564
rect 48240 4542 48360 4558
rect 48240 4146 48268 4542
rect 48412 4480 48464 4486
rect 48412 4422 48464 4428
rect 48424 4282 48452 4422
rect 48412 4276 48464 4282
rect 48412 4218 48464 4224
rect 48228 4140 48280 4146
rect 48228 4082 48280 4088
rect 48228 3936 48280 3942
rect 48228 3878 48280 3884
rect 48240 2990 48268 3878
rect 48412 3120 48464 3126
rect 48412 3062 48464 3068
rect 48228 2984 48280 2990
rect 48228 2926 48280 2932
rect 48228 2372 48280 2378
rect 48228 2314 48280 2320
rect 48240 2038 48268 2314
rect 48228 2032 48280 2038
rect 48228 1974 48280 1980
rect 48424 800 48452 3062
rect 48516 1970 48544 6598
rect 48964 6316 49016 6322
rect 48964 6258 49016 6264
rect 48596 6248 48648 6254
rect 48596 6190 48648 6196
rect 48608 5778 48636 6190
rect 48976 5914 49004 6258
rect 48964 5908 49016 5914
rect 48964 5850 49016 5856
rect 48596 5772 48648 5778
rect 48596 5714 48648 5720
rect 48688 5092 48740 5098
rect 48688 5034 48740 5040
rect 48596 4140 48648 4146
rect 48596 4082 48648 4088
rect 48608 3738 48636 4082
rect 48596 3732 48648 3738
rect 48596 3674 48648 3680
rect 48596 3188 48648 3194
rect 48596 3130 48648 3136
rect 48608 2446 48636 3130
rect 48596 2440 48648 2446
rect 48596 2382 48648 2388
rect 48504 1964 48556 1970
rect 48504 1906 48556 1912
rect 48700 800 48728 5034
rect 48780 3664 48832 3670
rect 48780 3606 48832 3612
rect 48976 3618 49004 5850
rect 49056 5024 49108 5030
rect 49056 4966 49108 4972
rect 49068 4146 49096 4966
rect 49436 4706 49464 6734
rect 49712 6730 49740 7686
rect 49804 7410 49832 7806
rect 49792 7404 49844 7410
rect 49792 7346 49844 7352
rect 49700 6724 49752 6730
rect 49700 6666 49752 6672
rect 49896 6322 49924 9454
rect 49988 8294 50016 9658
rect 50080 9178 50108 10678
rect 50172 10674 50200 11018
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 50632 10674 50660 11222
rect 50160 10668 50212 10674
rect 50160 10610 50212 10616
rect 50620 10668 50672 10674
rect 50620 10610 50672 10616
rect 50804 10668 50856 10674
rect 50804 10610 50856 10616
rect 50252 10260 50304 10266
rect 50172 10220 50252 10248
rect 50068 9172 50120 9178
rect 50068 9114 50120 9120
rect 50172 8634 50200 10220
rect 50252 10202 50304 10208
rect 50436 10124 50488 10130
rect 50436 10066 50488 10072
rect 50448 10033 50476 10066
rect 50434 10024 50490 10033
rect 50434 9959 50490 9968
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50632 9722 50660 10610
rect 50712 10600 50764 10606
rect 50712 10542 50764 10548
rect 50620 9716 50672 9722
rect 50620 9658 50672 9664
rect 50252 9648 50304 9654
rect 50252 9590 50304 9596
rect 50264 9450 50292 9590
rect 50252 9444 50304 9450
rect 50252 9386 50304 9392
rect 50528 9444 50580 9450
rect 50528 9386 50580 9392
rect 50540 8974 50568 9386
rect 50724 9382 50752 10542
rect 50816 9518 50844 10610
rect 50896 10464 50948 10470
rect 50896 10406 50948 10412
rect 50804 9512 50856 9518
rect 50804 9454 50856 9460
rect 50712 9376 50764 9382
rect 50712 9318 50764 9324
rect 50908 9178 50936 10406
rect 50986 10024 51042 10033
rect 50986 9959 51042 9968
rect 51000 9518 51028 9959
rect 51264 9920 51316 9926
rect 51264 9862 51316 9868
rect 51276 9654 51304 9862
rect 51264 9648 51316 9654
rect 51264 9590 51316 9596
rect 50988 9512 51040 9518
rect 50988 9454 51040 9460
rect 50988 9376 51040 9382
rect 50988 9318 51040 9324
rect 50896 9172 50948 9178
rect 50896 9114 50948 9120
rect 50804 9104 50856 9110
rect 50804 9046 50856 9052
rect 50528 8968 50580 8974
rect 50580 8916 50660 8922
rect 50528 8910 50660 8916
rect 50540 8894 50660 8910
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 50160 8628 50212 8634
rect 50160 8570 50212 8576
rect 49976 8288 50028 8294
rect 49976 8230 50028 8236
rect 50172 8090 50200 8570
rect 50632 8294 50660 8894
rect 50712 8832 50764 8838
rect 50712 8774 50764 8780
rect 50620 8288 50672 8294
rect 50620 8230 50672 8236
rect 50160 8084 50212 8090
rect 50160 8026 50212 8032
rect 50724 7886 50752 8774
rect 50816 8566 50844 9046
rect 50908 8974 50936 9114
rect 50896 8968 50948 8974
rect 50896 8910 50948 8916
rect 50908 8634 50936 8910
rect 51000 8906 51028 9318
rect 50988 8900 51040 8906
rect 50988 8842 51040 8848
rect 50896 8628 50948 8634
rect 50896 8570 50948 8576
rect 50804 8560 50856 8566
rect 50804 8502 50856 8508
rect 50712 7880 50764 7886
rect 50712 7822 50764 7828
rect 49976 7812 50028 7818
rect 49976 7754 50028 7760
rect 49988 7410 50016 7754
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 52736 7540 52788 7546
rect 52736 7482 52788 7488
rect 49976 7404 50028 7410
rect 49976 7346 50028 7352
rect 49988 6934 50016 7346
rect 49976 6928 50028 6934
rect 49976 6870 50028 6876
rect 49988 6746 50016 6870
rect 49988 6718 50108 6746
rect 49976 6656 50028 6662
rect 49976 6598 50028 6604
rect 49884 6316 49936 6322
rect 49884 6258 49936 6264
rect 49896 5574 49924 6258
rect 49884 5568 49936 5574
rect 49884 5510 49936 5516
rect 49516 5296 49568 5302
rect 49988 5250 50016 6598
rect 50080 6390 50108 6718
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50068 6384 50120 6390
rect 50068 6326 50120 6332
rect 51448 6316 51500 6322
rect 51448 6258 51500 6264
rect 50988 6180 51040 6186
rect 50988 6122 51040 6128
rect 50068 6112 50120 6118
rect 50068 6054 50120 6060
rect 50896 6112 50948 6118
rect 50896 6054 50948 6060
rect 50080 5778 50108 6054
rect 50068 5772 50120 5778
rect 50068 5714 50120 5720
rect 49516 5238 49568 5244
rect 49160 4678 49464 4706
rect 49056 4140 49108 4146
rect 49056 4082 49108 4088
rect 48792 3398 48820 3606
rect 48976 3602 49096 3618
rect 48872 3596 48924 3602
rect 48976 3596 49108 3602
rect 48976 3590 49056 3596
rect 48872 3538 48924 3544
rect 49056 3538 49108 3544
rect 48884 3505 48912 3538
rect 48870 3496 48926 3505
rect 48870 3431 48926 3440
rect 48780 3392 48832 3398
rect 48780 3334 48832 3340
rect 48962 2816 49018 2825
rect 48962 2751 49018 2760
rect 48976 2446 49004 2751
rect 48964 2440 49016 2446
rect 48964 2382 49016 2388
rect 49160 1834 49188 4678
rect 49528 4434 49556 5238
rect 49896 5234 50016 5250
rect 50080 5234 50108 5714
rect 50908 5710 50936 6054
rect 51000 5710 51028 6122
rect 51460 5914 51488 6258
rect 51448 5908 51500 5914
rect 51448 5850 51500 5856
rect 50896 5704 50948 5710
rect 50896 5646 50948 5652
rect 50988 5704 51040 5710
rect 50988 5646 51040 5652
rect 50160 5568 50212 5574
rect 50160 5510 50212 5516
rect 51356 5568 51408 5574
rect 51356 5510 51408 5516
rect 49884 5228 50016 5234
rect 49936 5222 50016 5228
rect 50068 5228 50120 5234
rect 49884 5170 49936 5176
rect 50068 5170 50120 5176
rect 49976 4752 50028 4758
rect 49976 4694 50028 4700
rect 49436 4406 49556 4434
rect 49332 4140 49384 4146
rect 49332 4082 49384 4088
rect 49344 3942 49372 4082
rect 49332 3936 49384 3942
rect 49332 3878 49384 3884
rect 49240 3596 49292 3602
rect 49240 3538 49292 3544
rect 49252 3126 49280 3538
rect 49240 3120 49292 3126
rect 49240 3062 49292 3068
rect 49344 3058 49372 3878
rect 49332 3052 49384 3058
rect 49332 2994 49384 3000
rect 49238 2816 49294 2825
rect 49238 2751 49294 2760
rect 49148 1828 49200 1834
rect 49148 1770 49200 1776
rect 48964 1624 49016 1630
rect 48964 1566 49016 1572
rect 48976 800 49004 1566
rect 49252 800 49280 2751
rect 49436 1442 49464 4406
rect 49516 4276 49568 4282
rect 49516 4218 49568 4224
rect 49528 3108 49556 4218
rect 49700 4072 49752 4078
rect 49700 4014 49752 4020
rect 49712 3194 49740 4014
rect 49792 3528 49844 3534
rect 49792 3470 49844 3476
rect 49700 3188 49752 3194
rect 49700 3130 49752 3136
rect 49608 3120 49660 3126
rect 49528 3080 49608 3108
rect 49528 2854 49556 3080
rect 49608 3062 49660 3068
rect 49516 2848 49568 2854
rect 49516 2790 49568 2796
rect 49608 2440 49660 2446
rect 49608 2382 49660 2388
rect 49620 1834 49648 2382
rect 49608 1828 49660 1834
rect 49608 1770 49660 1776
rect 49436 1414 49556 1442
rect 49528 800 49556 1414
rect 49804 800 49832 3470
rect 49988 2774 50016 4694
rect 50172 4128 50200 5510
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50620 5228 50672 5234
rect 50620 5170 50672 5176
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50080 4100 50292 4128
rect 50080 4010 50108 4100
rect 50068 4004 50120 4010
rect 50068 3946 50120 3952
rect 50160 4004 50212 4010
rect 50160 3946 50212 3952
rect 50080 3126 50108 3946
rect 50068 3120 50120 3126
rect 50068 3062 50120 3068
rect 49988 2746 50108 2774
rect 49884 2508 49936 2514
rect 49884 2450 49936 2456
rect 49896 2106 49924 2450
rect 49884 2100 49936 2106
rect 49884 2042 49936 2048
rect 50080 800 50108 2746
rect 50172 1442 50200 3946
rect 50264 3942 50292 4100
rect 50632 4078 50660 5170
rect 51172 4684 51224 4690
rect 51172 4626 51224 4632
rect 50896 4616 50948 4622
rect 50896 4558 50948 4564
rect 50712 4548 50764 4554
rect 50712 4490 50764 4496
rect 50620 4072 50672 4078
rect 50620 4014 50672 4020
rect 50252 3936 50304 3942
rect 50252 3878 50304 3884
rect 50344 3936 50396 3942
rect 50344 3878 50396 3884
rect 50356 3738 50384 3878
rect 50344 3732 50396 3738
rect 50344 3674 50396 3680
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 50724 3194 50752 4490
rect 50908 4282 50936 4558
rect 50896 4276 50948 4282
rect 50896 4218 50948 4224
rect 50804 4004 50856 4010
rect 50804 3946 50856 3952
rect 50816 3534 50844 3946
rect 50804 3528 50856 3534
rect 50804 3470 50856 3476
rect 50712 3188 50764 3194
rect 50712 3130 50764 3136
rect 51184 2922 51212 4626
rect 51264 3936 51316 3942
rect 51264 3878 51316 3884
rect 51276 3466 51304 3878
rect 51264 3460 51316 3466
rect 51264 3402 51316 3408
rect 50620 2916 50672 2922
rect 50620 2858 50672 2864
rect 51172 2916 51224 2922
rect 51172 2858 51224 2864
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 50172 1414 50384 1442
rect 50356 800 50384 1414
rect 50632 800 50660 2858
rect 51080 2848 51132 2854
rect 51080 2790 51132 2796
rect 51092 2514 51120 2790
rect 51080 2508 51132 2514
rect 51080 2450 51132 2456
rect 51276 2446 51304 3402
rect 51264 2440 51316 2446
rect 51264 2382 51316 2388
rect 51368 2378 51396 5510
rect 51724 5024 51776 5030
rect 51724 4966 51776 4972
rect 51632 4480 51684 4486
rect 51632 4422 51684 4428
rect 51448 2848 51500 2854
rect 51448 2790 51500 2796
rect 51356 2372 51408 2378
rect 51356 2314 51408 2320
rect 50896 2304 50948 2310
rect 50896 2246 50948 2252
rect 51172 2304 51224 2310
rect 51172 2246 51224 2252
rect 50908 800 50936 2246
rect 51184 800 51212 2246
rect 51460 800 51488 2790
rect 51644 2446 51672 4422
rect 51736 3602 51764 4966
rect 52092 4480 52144 4486
rect 52092 4422 52144 4428
rect 51908 3936 51960 3942
rect 51908 3878 51960 3884
rect 51816 3732 51868 3738
rect 51816 3674 51868 3680
rect 51724 3596 51776 3602
rect 51724 3538 51776 3544
rect 51828 3058 51856 3674
rect 51816 3052 51868 3058
rect 51816 2994 51868 3000
rect 51724 2984 51776 2990
rect 51724 2926 51776 2932
rect 51632 2440 51684 2446
rect 51632 2382 51684 2388
rect 51736 800 51764 2926
rect 51920 2825 51948 3878
rect 52104 3534 52132 4422
rect 52092 3528 52144 3534
rect 52092 3470 52144 3476
rect 52368 3528 52420 3534
rect 52368 3470 52420 3476
rect 52276 2848 52328 2854
rect 51906 2816 51962 2825
rect 52276 2790 52328 2796
rect 51906 2751 51962 2760
rect 52000 2304 52052 2310
rect 52000 2246 52052 2252
rect 52012 800 52040 2246
rect 52288 800 52316 2790
rect 52380 1630 52408 3470
rect 52748 3058 52776 7482
rect 54024 6248 54076 6254
rect 54024 6190 54076 6196
rect 53288 5024 53340 5030
rect 53288 4966 53340 4972
rect 52736 3052 52788 3058
rect 52736 2994 52788 3000
rect 52828 2916 52880 2922
rect 52828 2858 52880 2864
rect 52552 2576 52604 2582
rect 52552 2518 52604 2524
rect 52368 1624 52420 1630
rect 52368 1566 52420 1572
rect 52564 800 52592 2518
rect 52840 800 52868 2858
rect 53300 2446 53328 4966
rect 54036 4826 54064 6190
rect 54588 4826 54616 28494
rect 57716 23730 57744 31758
rect 65654 31036 65962 31045
rect 65654 31034 65660 31036
rect 65716 31034 65740 31036
rect 65796 31034 65820 31036
rect 65876 31034 65900 31036
rect 65956 31034 65962 31036
rect 65716 30982 65718 31034
rect 65898 30982 65900 31034
rect 65654 30980 65660 30982
rect 65716 30980 65740 30982
rect 65796 30980 65820 30982
rect 65876 30980 65900 30982
rect 65956 30980 65962 30982
rect 65654 30971 65962 30980
rect 65654 29948 65962 29957
rect 65654 29946 65660 29948
rect 65716 29946 65740 29948
rect 65796 29946 65820 29948
rect 65876 29946 65900 29948
rect 65956 29946 65962 29948
rect 65716 29894 65718 29946
rect 65898 29894 65900 29946
rect 65654 29892 65660 29894
rect 65716 29892 65740 29894
rect 65796 29892 65820 29894
rect 65876 29892 65900 29894
rect 65956 29892 65962 29894
rect 65654 29883 65962 29892
rect 61384 29640 61436 29646
rect 61384 29582 61436 29588
rect 60556 25288 60608 25294
rect 60556 25230 60608 25236
rect 57704 23724 57756 23730
rect 57704 23666 57756 23672
rect 60568 20262 60596 25230
rect 55128 20256 55180 20262
rect 55128 20198 55180 20204
rect 60556 20256 60608 20262
rect 60556 20198 60608 20204
rect 55140 18630 55168 20198
rect 55128 18624 55180 18630
rect 55128 18566 55180 18572
rect 55772 18624 55824 18630
rect 55772 18566 55824 18572
rect 54668 17672 54720 17678
rect 54668 17614 54720 17620
rect 54680 8022 54708 17614
rect 55312 17264 55364 17270
rect 55312 17206 55364 17212
rect 54668 8016 54720 8022
rect 54668 7958 54720 7964
rect 54024 4820 54076 4826
rect 54024 4762 54076 4768
rect 54576 4820 54628 4826
rect 54576 4762 54628 4768
rect 54036 4282 54064 4762
rect 54024 4276 54076 4282
rect 54024 4218 54076 4224
rect 53470 3496 53526 3505
rect 53470 3431 53472 3440
rect 53524 3431 53526 3440
rect 53472 3402 53524 3408
rect 53932 3392 53984 3398
rect 53932 3334 53984 3340
rect 53380 2848 53432 2854
rect 53380 2790 53432 2796
rect 53288 2440 53340 2446
rect 53288 2382 53340 2388
rect 53104 2304 53156 2310
rect 53104 2246 53156 2252
rect 53116 800 53144 2246
rect 53392 800 53420 2790
rect 53656 2372 53708 2378
rect 53656 2314 53708 2320
rect 53668 800 53696 2314
rect 53944 800 53972 3334
rect 54036 2514 54064 4218
rect 54484 3596 54536 3602
rect 54484 3538 54536 3544
rect 54208 2916 54260 2922
rect 54208 2858 54260 2864
rect 54024 2508 54076 2514
rect 54024 2450 54076 2456
rect 54220 800 54248 2858
rect 54496 800 54524 3538
rect 54588 3534 54616 4762
rect 54680 4146 54708 7958
rect 55220 5636 55272 5642
rect 55220 5578 55272 5584
rect 55232 4146 55260 5578
rect 55324 4826 55352 17206
rect 55312 4820 55364 4826
rect 55312 4762 55364 4768
rect 54668 4140 54720 4146
rect 55220 4140 55272 4146
rect 54668 4082 54720 4088
rect 55140 4100 55220 4128
rect 54576 3528 54628 3534
rect 54576 3470 54628 3476
rect 54680 3126 54708 4082
rect 54668 3120 54720 3126
rect 54668 3062 54720 3068
rect 54760 3120 54812 3126
rect 54760 3062 54812 3068
rect 54772 800 54800 3062
rect 55140 3058 55168 4100
rect 55220 4082 55272 4088
rect 55232 4017 55260 4082
rect 55324 3058 55352 4762
rect 55784 4146 55812 18566
rect 56324 14544 56376 14550
rect 56324 14486 56376 14492
rect 55956 4480 56008 4486
rect 55956 4422 56008 4428
rect 55772 4140 55824 4146
rect 55772 4082 55824 4088
rect 55404 3528 55456 3534
rect 55404 3470 55456 3476
rect 55128 3052 55180 3058
rect 55128 2994 55180 3000
rect 55312 3052 55364 3058
rect 55312 2994 55364 3000
rect 55128 2916 55180 2922
rect 55048 2876 55128 2904
rect 55048 800 55076 2876
rect 55128 2858 55180 2864
rect 55416 1850 55444 3470
rect 55588 2848 55640 2854
rect 55588 2790 55640 2796
rect 55496 2372 55548 2378
rect 55496 2314 55548 2320
rect 55324 1822 55444 1850
rect 55324 800 55352 1822
rect 55508 800 55536 2314
rect 55600 800 55628 2790
rect 55784 2514 55812 4082
rect 55864 3596 55916 3602
rect 55864 3538 55916 3544
rect 55772 2508 55824 2514
rect 55772 2450 55824 2456
rect 55876 800 55904 3538
rect 55968 2378 55996 4422
rect 56336 4146 56364 14486
rect 61396 5642 61424 29582
rect 65654 28860 65962 28869
rect 65654 28858 65660 28860
rect 65716 28858 65740 28860
rect 65796 28858 65820 28860
rect 65876 28858 65900 28860
rect 65956 28858 65962 28860
rect 65716 28806 65718 28858
rect 65898 28806 65900 28858
rect 65654 28804 65660 28806
rect 65716 28804 65740 28806
rect 65796 28804 65820 28806
rect 65876 28804 65900 28806
rect 65956 28804 65962 28806
rect 65654 28795 65962 28804
rect 67192 28558 67220 39374
rect 67284 31958 67312 41414
rect 67468 39642 67496 48690
rect 67546 48648 67602 48657
rect 67546 48583 67548 48592
rect 67600 48583 67602 48592
rect 67548 48554 67600 48560
rect 68008 41472 68060 41478
rect 68008 41414 68060 41420
rect 68020 41177 68048 41414
rect 68006 41168 68062 41177
rect 68006 41103 68062 41112
rect 67456 39636 67508 39642
rect 67456 39578 67508 39584
rect 67364 33992 67416 33998
rect 67364 33934 67416 33940
rect 67272 31952 67324 31958
rect 67272 31894 67324 31900
rect 67376 29850 67404 33934
rect 68008 33856 68060 33862
rect 68008 33798 68060 33804
rect 68020 33697 68048 33798
rect 68006 33688 68062 33697
rect 68006 33623 68062 33632
rect 67364 29844 67416 29850
rect 67364 29786 67416 29792
rect 67180 28552 67232 28558
rect 67180 28494 67232 28500
rect 65654 27772 65962 27781
rect 65654 27770 65660 27772
rect 65716 27770 65740 27772
rect 65796 27770 65820 27772
rect 65876 27770 65900 27772
rect 65956 27770 65962 27772
rect 65716 27718 65718 27770
rect 65898 27718 65900 27770
rect 65654 27716 65660 27718
rect 65716 27716 65740 27718
rect 65796 27716 65820 27718
rect 65876 27716 65900 27718
rect 65956 27716 65962 27718
rect 65654 27707 65962 27716
rect 65654 26684 65962 26693
rect 65654 26682 65660 26684
rect 65716 26682 65740 26684
rect 65796 26682 65820 26684
rect 65876 26682 65900 26684
rect 65956 26682 65962 26684
rect 65716 26630 65718 26682
rect 65898 26630 65900 26682
rect 65654 26628 65660 26630
rect 65716 26628 65740 26630
rect 65796 26628 65820 26630
rect 65876 26628 65900 26630
rect 65956 26628 65962 26630
rect 65654 26619 65962 26628
rect 68008 26512 68060 26518
rect 68008 26454 68060 26460
rect 67824 26376 67876 26382
rect 67824 26318 67876 26324
rect 65654 25596 65962 25605
rect 65654 25594 65660 25596
rect 65716 25594 65740 25596
rect 65796 25594 65820 25596
rect 65876 25594 65900 25596
rect 65956 25594 65962 25596
rect 65716 25542 65718 25594
rect 65898 25542 65900 25594
rect 65654 25540 65660 25542
rect 65716 25540 65740 25542
rect 65796 25540 65820 25542
rect 65876 25540 65900 25542
rect 65956 25540 65962 25542
rect 65654 25531 65962 25540
rect 67836 25226 67864 26318
rect 68020 26217 68048 26454
rect 68006 26208 68062 26217
rect 68006 26143 68062 26152
rect 67824 25220 67876 25226
rect 67824 25162 67876 25168
rect 65654 24508 65962 24517
rect 65654 24506 65660 24508
rect 65716 24506 65740 24508
rect 65796 24506 65820 24508
rect 65876 24506 65900 24508
rect 65956 24506 65962 24508
rect 65716 24454 65718 24506
rect 65898 24454 65900 24506
rect 65654 24452 65660 24454
rect 65716 24452 65740 24454
rect 65796 24452 65820 24454
rect 65876 24452 65900 24454
rect 65956 24452 65962 24454
rect 65654 24443 65962 24452
rect 65654 23420 65962 23429
rect 65654 23418 65660 23420
rect 65716 23418 65740 23420
rect 65796 23418 65820 23420
rect 65876 23418 65900 23420
rect 65956 23418 65962 23420
rect 65716 23366 65718 23418
rect 65898 23366 65900 23418
rect 65654 23364 65660 23366
rect 65716 23364 65740 23366
rect 65796 23364 65820 23366
rect 65876 23364 65900 23366
rect 65956 23364 65962 23366
rect 65654 23355 65962 23364
rect 65654 22332 65962 22341
rect 65654 22330 65660 22332
rect 65716 22330 65740 22332
rect 65796 22330 65820 22332
rect 65876 22330 65900 22332
rect 65956 22330 65962 22332
rect 65716 22278 65718 22330
rect 65898 22278 65900 22330
rect 65654 22276 65660 22278
rect 65716 22276 65740 22278
rect 65796 22276 65820 22278
rect 65876 22276 65900 22278
rect 65956 22276 65962 22278
rect 65654 22267 65962 22276
rect 65654 21244 65962 21253
rect 65654 21242 65660 21244
rect 65716 21242 65740 21244
rect 65796 21242 65820 21244
rect 65876 21242 65900 21244
rect 65956 21242 65962 21244
rect 65716 21190 65718 21242
rect 65898 21190 65900 21242
rect 65654 21188 65660 21190
rect 65716 21188 65740 21190
rect 65796 21188 65820 21190
rect 65876 21188 65900 21190
rect 65956 21188 65962 21190
rect 65654 21179 65962 21188
rect 65654 20156 65962 20165
rect 65654 20154 65660 20156
rect 65716 20154 65740 20156
rect 65796 20154 65820 20156
rect 65876 20154 65900 20156
rect 65956 20154 65962 20156
rect 65716 20102 65718 20154
rect 65898 20102 65900 20154
rect 65654 20100 65660 20102
rect 65716 20100 65740 20102
rect 65796 20100 65820 20102
rect 65876 20100 65900 20102
rect 65956 20100 65962 20102
rect 65654 20091 65962 20100
rect 65654 19068 65962 19077
rect 65654 19066 65660 19068
rect 65716 19066 65740 19068
rect 65796 19066 65820 19068
rect 65876 19066 65900 19068
rect 65956 19066 65962 19068
rect 65716 19014 65718 19066
rect 65898 19014 65900 19066
rect 65654 19012 65660 19014
rect 65716 19012 65740 19014
rect 65796 19012 65820 19014
rect 65876 19012 65900 19014
rect 65956 19012 65962 19014
rect 65654 19003 65962 19012
rect 67824 18760 67876 18766
rect 67824 18702 67876 18708
rect 68006 18728 68062 18737
rect 65654 17980 65962 17989
rect 65654 17978 65660 17980
rect 65716 17978 65740 17980
rect 65796 17978 65820 17980
rect 65876 17978 65900 17980
rect 65956 17978 65962 17980
rect 65716 17926 65718 17978
rect 65898 17926 65900 17978
rect 65654 17924 65660 17926
rect 65716 17924 65740 17926
rect 65796 17924 65820 17926
rect 65876 17924 65900 17926
rect 65956 17924 65962 17926
rect 65654 17915 65962 17924
rect 67836 17610 67864 18702
rect 68006 18663 68062 18672
rect 68020 18630 68048 18663
rect 68008 18624 68060 18630
rect 68008 18566 68060 18572
rect 67824 17604 67876 17610
rect 67824 17546 67876 17552
rect 65654 16892 65962 16901
rect 65654 16890 65660 16892
rect 65716 16890 65740 16892
rect 65796 16890 65820 16892
rect 65876 16890 65900 16892
rect 65956 16890 65962 16892
rect 65716 16838 65718 16890
rect 65898 16838 65900 16890
rect 65654 16836 65660 16838
rect 65716 16836 65740 16838
rect 65796 16836 65820 16838
rect 65876 16836 65900 16838
rect 65956 16836 65962 16838
rect 65654 16827 65962 16836
rect 65654 15804 65962 15813
rect 65654 15802 65660 15804
rect 65716 15802 65740 15804
rect 65796 15802 65820 15804
rect 65876 15802 65900 15804
rect 65956 15802 65962 15804
rect 65716 15750 65718 15802
rect 65898 15750 65900 15802
rect 65654 15748 65660 15750
rect 65716 15748 65740 15750
rect 65796 15748 65820 15750
rect 65876 15748 65900 15750
rect 65956 15748 65962 15750
rect 65654 15739 65962 15748
rect 65654 14716 65962 14725
rect 65654 14714 65660 14716
rect 65716 14714 65740 14716
rect 65796 14714 65820 14716
rect 65876 14714 65900 14716
rect 65956 14714 65962 14716
rect 65716 14662 65718 14714
rect 65898 14662 65900 14714
rect 65654 14660 65660 14662
rect 65716 14660 65740 14662
rect 65796 14660 65820 14662
rect 65876 14660 65900 14662
rect 65956 14660 65962 14662
rect 65654 14651 65962 14660
rect 65654 13628 65962 13637
rect 65654 13626 65660 13628
rect 65716 13626 65740 13628
rect 65796 13626 65820 13628
rect 65876 13626 65900 13628
rect 65956 13626 65962 13628
rect 65716 13574 65718 13626
rect 65898 13574 65900 13626
rect 65654 13572 65660 13574
rect 65716 13572 65740 13574
rect 65796 13572 65820 13574
rect 65876 13572 65900 13574
rect 65956 13572 65962 13574
rect 65654 13563 65962 13572
rect 65654 12540 65962 12549
rect 65654 12538 65660 12540
rect 65716 12538 65740 12540
rect 65796 12538 65820 12540
rect 65876 12538 65900 12540
rect 65956 12538 65962 12540
rect 65716 12486 65718 12538
rect 65898 12486 65900 12538
rect 65654 12484 65660 12486
rect 65716 12484 65740 12486
rect 65796 12484 65820 12486
rect 65876 12484 65900 12486
rect 65956 12484 65962 12486
rect 65654 12475 65962 12484
rect 67364 11756 67416 11762
rect 67364 11698 67416 11704
rect 65654 11452 65962 11461
rect 65654 11450 65660 11452
rect 65716 11450 65740 11452
rect 65796 11450 65820 11452
rect 65876 11450 65900 11452
rect 65956 11450 65962 11452
rect 65716 11398 65718 11450
rect 65898 11398 65900 11450
rect 65654 11396 65660 11398
rect 65716 11396 65740 11398
rect 65796 11396 65820 11398
rect 65876 11396 65900 11398
rect 65956 11396 65962 11398
rect 65654 11387 65962 11396
rect 67376 11354 67404 11698
rect 67548 11552 67600 11558
rect 67548 11494 67600 11500
rect 67364 11348 67416 11354
rect 67364 11290 67416 11296
rect 67560 11257 67588 11494
rect 67546 11248 67602 11257
rect 67546 11183 67602 11192
rect 65654 10364 65962 10373
rect 65654 10362 65660 10364
rect 65716 10362 65740 10364
rect 65796 10362 65820 10364
rect 65876 10362 65900 10364
rect 65956 10362 65962 10364
rect 65716 10310 65718 10362
rect 65898 10310 65900 10362
rect 65654 10308 65660 10310
rect 65716 10308 65740 10310
rect 65796 10308 65820 10310
rect 65876 10308 65900 10310
rect 65956 10308 65962 10310
rect 65654 10299 65962 10308
rect 65654 9276 65962 9285
rect 65654 9274 65660 9276
rect 65716 9274 65740 9276
rect 65796 9274 65820 9276
rect 65876 9274 65900 9276
rect 65956 9274 65962 9276
rect 65716 9222 65718 9274
rect 65898 9222 65900 9274
rect 65654 9220 65660 9222
rect 65716 9220 65740 9222
rect 65796 9220 65820 9222
rect 65876 9220 65900 9222
rect 65956 9220 65962 9222
rect 65654 9211 65962 9220
rect 65654 8188 65962 8197
rect 65654 8186 65660 8188
rect 65716 8186 65740 8188
rect 65796 8186 65820 8188
rect 65876 8186 65900 8188
rect 65956 8186 65962 8188
rect 65716 8134 65718 8186
rect 65898 8134 65900 8186
rect 65654 8132 65660 8134
rect 65716 8132 65740 8134
rect 65796 8132 65820 8134
rect 65876 8132 65900 8134
rect 65956 8132 65962 8134
rect 65654 8123 65962 8132
rect 65654 7100 65962 7109
rect 65654 7098 65660 7100
rect 65716 7098 65740 7100
rect 65796 7098 65820 7100
rect 65876 7098 65900 7100
rect 65956 7098 65962 7100
rect 65716 7046 65718 7098
rect 65898 7046 65900 7098
rect 65654 7044 65660 7046
rect 65716 7044 65740 7046
rect 65796 7044 65820 7046
rect 65876 7044 65900 7046
rect 65956 7044 65962 7046
rect 65654 7035 65962 7044
rect 65654 6012 65962 6021
rect 65654 6010 65660 6012
rect 65716 6010 65740 6012
rect 65796 6010 65820 6012
rect 65876 6010 65900 6012
rect 65956 6010 65962 6012
rect 65716 5958 65718 6010
rect 65898 5958 65900 6010
rect 65654 5956 65660 5958
rect 65716 5956 65740 5958
rect 65796 5956 65820 5958
rect 65876 5956 65900 5958
rect 65956 5956 65962 5958
rect 65654 5947 65962 5956
rect 61384 5636 61436 5642
rect 61384 5578 61436 5584
rect 65654 4924 65962 4933
rect 65654 4922 65660 4924
rect 65716 4922 65740 4924
rect 65796 4922 65820 4924
rect 65876 4922 65900 4924
rect 65956 4922 65962 4924
rect 65716 4870 65718 4922
rect 65898 4870 65900 4922
rect 65654 4868 65660 4870
rect 65716 4868 65740 4870
rect 65796 4868 65820 4870
rect 65876 4868 65900 4870
rect 65956 4868 65962 4870
rect 65654 4859 65962 4868
rect 67180 4276 67232 4282
rect 67180 4218 67232 4224
rect 56324 4140 56376 4146
rect 56324 4082 56376 4088
rect 56336 2446 56364 4082
rect 65654 3836 65962 3845
rect 65654 3834 65660 3836
rect 65716 3834 65740 3836
rect 65796 3834 65820 3836
rect 65876 3834 65900 3836
rect 65956 3834 65962 3836
rect 65716 3782 65718 3834
rect 65898 3782 65900 3834
rect 65654 3780 65660 3782
rect 65716 3780 65740 3782
rect 65796 3780 65820 3782
rect 65876 3780 65900 3782
rect 65956 3780 65962 3782
rect 65654 3771 65962 3780
rect 57244 3664 57296 3670
rect 57244 3606 57296 3612
rect 56416 3528 56468 3534
rect 56416 3470 56468 3476
rect 56324 2440 56376 2446
rect 56324 2382 56376 2388
rect 55956 2372 56008 2378
rect 55956 2314 56008 2320
rect 56140 2304 56192 2310
rect 56140 2246 56192 2252
rect 56152 800 56180 2246
rect 56428 800 56456 3470
rect 56784 3120 56836 3126
rect 56784 3062 56836 3068
rect 56796 2650 56824 3062
rect 56968 2984 57020 2990
rect 56968 2926 57020 2932
rect 56784 2644 56836 2650
rect 56784 2586 56836 2592
rect 56692 2576 56744 2582
rect 56692 2518 56744 2524
rect 56704 800 56732 2518
rect 56980 800 57008 2926
rect 57256 800 57284 3606
rect 57612 3596 57664 3602
rect 57612 3538 57664 3544
rect 57520 2916 57572 2922
rect 57520 2858 57572 2864
rect 57428 2508 57480 2514
rect 57428 2450 57480 2456
rect 57440 800 57468 2450
rect 57532 800 57560 2858
rect 57624 800 57652 3538
rect 67192 3534 67220 4218
rect 67364 4140 67416 4146
rect 67364 4082 67416 4088
rect 67376 3738 67404 4082
rect 67548 3936 67600 3942
rect 67548 3878 67600 3884
rect 67560 3777 67588 3878
rect 67546 3768 67602 3777
rect 67364 3732 67416 3738
rect 67546 3703 67602 3712
rect 67364 3674 67416 3680
rect 67180 3528 67232 3534
rect 67180 3470 67232 3476
rect 65654 2748 65962 2757
rect 65654 2746 65660 2748
rect 65716 2746 65740 2748
rect 65796 2746 65820 2748
rect 65876 2746 65900 2748
rect 65956 2746 65962 2748
rect 65716 2694 65718 2746
rect 65898 2694 65900 2746
rect 65654 2692 65660 2694
rect 65716 2692 65740 2694
rect 65796 2692 65820 2694
rect 65876 2692 65900 2694
rect 65956 2692 65962 2694
rect 65654 2683 65962 2692
rect 11808 734 12296 762
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 52918 0 52974 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53194 0 53250 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53470 0 53526 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53838 0 53894 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54114 0 54170 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 54390 0 54446 800
rect 54482 0 54538 800
rect 54574 0 54630 800
rect 54666 0 54722 800
rect 54758 0 54814 800
rect 54850 0 54906 800
rect 54942 0 54998 800
rect 55034 0 55090 800
rect 55126 0 55182 800
rect 55218 0 55274 800
rect 55310 0 55366 800
rect 55402 0 55458 800
rect 55494 0 55550 800
rect 55586 0 55642 800
rect 55678 0 55734 800
rect 55770 0 55826 800
rect 55862 0 55918 800
rect 55954 0 56010 800
rect 56046 0 56102 800
rect 56138 0 56194 800
rect 56230 0 56286 800
rect 56322 0 56378 800
rect 56414 0 56470 800
rect 56506 0 56562 800
rect 56598 0 56654 800
rect 56690 0 56746 800
rect 56782 0 56838 800
rect 56874 0 56930 800
rect 56966 0 57022 800
rect 57058 0 57114 800
rect 57150 0 57206 800
rect 57242 0 57298 800
rect 57334 0 57390 800
rect 57426 0 57482 800
rect 57518 0 57574 800
rect 57610 0 57666 800
<< via2 >>
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 65660 57146 65716 57148
rect 65740 57146 65796 57148
rect 65820 57146 65876 57148
rect 65900 57146 65956 57148
rect 65660 57094 65706 57146
rect 65706 57094 65716 57146
rect 65740 57094 65770 57146
rect 65770 57094 65782 57146
rect 65782 57094 65796 57146
rect 65820 57094 65834 57146
rect 65834 57094 65846 57146
rect 65846 57094 65876 57146
rect 65900 57094 65910 57146
rect 65910 57094 65956 57146
rect 65660 57092 65716 57094
rect 65740 57092 65796 57094
rect 65820 57092 65876 57094
rect 65900 57092 65956 57094
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 65660 56058 65716 56060
rect 65740 56058 65796 56060
rect 65820 56058 65876 56060
rect 65900 56058 65956 56060
rect 65660 56006 65706 56058
rect 65706 56006 65716 56058
rect 65740 56006 65770 56058
rect 65770 56006 65782 56058
rect 65782 56006 65796 56058
rect 65820 56006 65834 56058
rect 65834 56006 65846 56058
rect 65846 56006 65876 56058
rect 65900 56006 65910 56058
rect 65910 56006 65956 56058
rect 65660 56004 65716 56006
rect 65740 56004 65796 56006
rect 65820 56004 65876 56006
rect 65900 56004 65956 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 65660 54970 65716 54972
rect 65740 54970 65796 54972
rect 65820 54970 65876 54972
rect 65900 54970 65956 54972
rect 65660 54918 65706 54970
rect 65706 54918 65716 54970
rect 65740 54918 65770 54970
rect 65770 54918 65782 54970
rect 65782 54918 65796 54970
rect 65820 54918 65834 54970
rect 65834 54918 65846 54970
rect 65846 54918 65876 54970
rect 65900 54918 65910 54970
rect 65910 54918 65956 54970
rect 65660 54916 65716 54918
rect 65740 54916 65796 54918
rect 65820 54916 65876 54918
rect 65900 54916 65956 54918
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 65660 53882 65716 53884
rect 65740 53882 65796 53884
rect 65820 53882 65876 53884
rect 65900 53882 65956 53884
rect 65660 53830 65706 53882
rect 65706 53830 65716 53882
rect 65740 53830 65770 53882
rect 65770 53830 65782 53882
rect 65782 53830 65796 53882
rect 65820 53830 65834 53882
rect 65834 53830 65846 53882
rect 65846 53830 65876 53882
rect 65900 53830 65910 53882
rect 65910 53830 65956 53882
rect 65660 53828 65716 53830
rect 65740 53828 65796 53830
rect 65820 53828 65876 53830
rect 65900 53828 65956 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 65660 52794 65716 52796
rect 65740 52794 65796 52796
rect 65820 52794 65876 52796
rect 65900 52794 65956 52796
rect 65660 52742 65706 52794
rect 65706 52742 65716 52794
rect 65740 52742 65770 52794
rect 65770 52742 65782 52794
rect 65782 52742 65796 52794
rect 65820 52742 65834 52794
rect 65834 52742 65846 52794
rect 65846 52742 65876 52794
rect 65900 52742 65910 52794
rect 65910 52742 65956 52794
rect 65660 52740 65716 52742
rect 65740 52740 65796 52742
rect 65820 52740 65876 52742
rect 65900 52740 65956 52742
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 65660 51706 65716 51708
rect 65740 51706 65796 51708
rect 65820 51706 65876 51708
rect 65900 51706 65956 51708
rect 65660 51654 65706 51706
rect 65706 51654 65716 51706
rect 65740 51654 65770 51706
rect 65770 51654 65782 51706
rect 65782 51654 65796 51706
rect 65820 51654 65834 51706
rect 65834 51654 65846 51706
rect 65846 51654 65876 51706
rect 65900 51654 65910 51706
rect 65910 51654 65956 51706
rect 65660 51652 65716 51654
rect 65740 51652 65796 51654
rect 65820 51652 65876 51654
rect 65900 51652 65956 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 65660 50618 65716 50620
rect 65740 50618 65796 50620
rect 65820 50618 65876 50620
rect 65900 50618 65956 50620
rect 65660 50566 65706 50618
rect 65706 50566 65716 50618
rect 65740 50566 65770 50618
rect 65770 50566 65782 50618
rect 65782 50566 65796 50618
rect 65820 50566 65834 50618
rect 65834 50566 65846 50618
rect 65846 50566 65876 50618
rect 65900 50566 65910 50618
rect 65910 50566 65956 50618
rect 65660 50564 65716 50566
rect 65740 50564 65796 50566
rect 65820 50564 65876 50566
rect 65900 50564 65956 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 65660 49530 65716 49532
rect 65740 49530 65796 49532
rect 65820 49530 65876 49532
rect 65900 49530 65956 49532
rect 65660 49478 65706 49530
rect 65706 49478 65716 49530
rect 65740 49478 65770 49530
rect 65770 49478 65782 49530
rect 65782 49478 65796 49530
rect 65820 49478 65834 49530
rect 65834 49478 65846 49530
rect 65846 49478 65876 49530
rect 65900 49478 65910 49530
rect 65910 49478 65956 49530
rect 65660 49476 65716 49478
rect 65740 49476 65796 49478
rect 65820 49476 65876 49478
rect 65900 49476 65956 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 65660 48442 65716 48444
rect 65740 48442 65796 48444
rect 65820 48442 65876 48444
rect 65900 48442 65956 48444
rect 65660 48390 65706 48442
rect 65706 48390 65716 48442
rect 65740 48390 65770 48442
rect 65770 48390 65782 48442
rect 65782 48390 65796 48442
rect 65820 48390 65834 48442
rect 65834 48390 65846 48442
rect 65846 48390 65876 48442
rect 65900 48390 65910 48442
rect 65910 48390 65956 48442
rect 65660 48388 65716 48390
rect 65740 48388 65796 48390
rect 65820 48388 65876 48390
rect 65900 48388 65956 48390
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 65660 47354 65716 47356
rect 65740 47354 65796 47356
rect 65820 47354 65876 47356
rect 65900 47354 65956 47356
rect 65660 47302 65706 47354
rect 65706 47302 65716 47354
rect 65740 47302 65770 47354
rect 65770 47302 65782 47354
rect 65782 47302 65796 47354
rect 65820 47302 65834 47354
rect 65834 47302 65846 47354
rect 65846 47302 65876 47354
rect 65900 47302 65910 47354
rect 65910 47302 65956 47354
rect 65660 47300 65716 47302
rect 65740 47300 65796 47302
rect 65820 47300 65876 47302
rect 65900 47300 65956 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 65660 46266 65716 46268
rect 65740 46266 65796 46268
rect 65820 46266 65876 46268
rect 65900 46266 65956 46268
rect 65660 46214 65706 46266
rect 65706 46214 65716 46266
rect 65740 46214 65770 46266
rect 65770 46214 65782 46266
rect 65782 46214 65796 46266
rect 65820 46214 65834 46266
rect 65834 46214 65846 46266
rect 65846 46214 65876 46266
rect 65900 46214 65910 46266
rect 65910 46214 65956 46266
rect 65660 46212 65716 46214
rect 65740 46212 65796 46214
rect 65820 46212 65876 46214
rect 65900 46212 65956 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 67546 56108 67548 56128
rect 67548 56108 67600 56128
rect 67600 56108 67602 56128
rect 67546 56072 67602 56108
rect 65660 45178 65716 45180
rect 65740 45178 65796 45180
rect 65820 45178 65876 45180
rect 65900 45178 65956 45180
rect 65660 45126 65706 45178
rect 65706 45126 65716 45178
rect 65740 45126 65770 45178
rect 65770 45126 65782 45178
rect 65782 45126 65796 45178
rect 65820 45126 65834 45178
rect 65834 45126 65846 45178
rect 65846 45126 65876 45178
rect 65900 45126 65910 45178
rect 65910 45126 65956 45178
rect 65660 45124 65716 45126
rect 65740 45124 65796 45126
rect 65820 45124 65876 45126
rect 65900 45124 65956 45126
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 65660 44090 65716 44092
rect 65740 44090 65796 44092
rect 65820 44090 65876 44092
rect 65900 44090 65956 44092
rect 65660 44038 65706 44090
rect 65706 44038 65716 44090
rect 65740 44038 65770 44090
rect 65770 44038 65782 44090
rect 65782 44038 65796 44090
rect 65820 44038 65834 44090
rect 65834 44038 65846 44090
rect 65846 44038 65876 44090
rect 65900 44038 65910 44090
rect 65910 44038 65956 44090
rect 65660 44036 65716 44038
rect 65740 44036 65796 44038
rect 65820 44036 65876 44038
rect 65900 44036 65956 44038
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 65660 43002 65716 43004
rect 65740 43002 65796 43004
rect 65820 43002 65876 43004
rect 65900 43002 65956 43004
rect 65660 42950 65706 43002
rect 65706 42950 65716 43002
rect 65740 42950 65770 43002
rect 65770 42950 65782 43002
rect 65782 42950 65796 43002
rect 65820 42950 65834 43002
rect 65834 42950 65846 43002
rect 65846 42950 65876 43002
rect 65900 42950 65910 43002
rect 65910 42950 65956 43002
rect 65660 42948 65716 42950
rect 65740 42948 65796 42950
rect 65820 42948 65876 42950
rect 65900 42948 65956 42950
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 65660 41914 65716 41916
rect 65740 41914 65796 41916
rect 65820 41914 65876 41916
rect 65900 41914 65956 41916
rect 65660 41862 65706 41914
rect 65706 41862 65716 41914
rect 65740 41862 65770 41914
rect 65770 41862 65782 41914
rect 65782 41862 65796 41914
rect 65820 41862 65834 41914
rect 65834 41862 65846 41914
rect 65846 41862 65876 41914
rect 65900 41862 65910 41914
rect 65910 41862 65956 41914
rect 65660 41860 65716 41862
rect 65740 41860 65796 41862
rect 65820 41860 65876 41862
rect 65900 41860 65956 41862
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 65660 40826 65716 40828
rect 65740 40826 65796 40828
rect 65820 40826 65876 40828
rect 65900 40826 65956 40828
rect 65660 40774 65706 40826
rect 65706 40774 65716 40826
rect 65740 40774 65770 40826
rect 65770 40774 65782 40826
rect 65782 40774 65796 40826
rect 65820 40774 65834 40826
rect 65834 40774 65846 40826
rect 65846 40774 65876 40826
rect 65900 40774 65910 40826
rect 65910 40774 65956 40826
rect 65660 40772 65716 40774
rect 65740 40772 65796 40774
rect 65820 40772 65876 40774
rect 65900 40772 65956 40774
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 65660 39738 65716 39740
rect 65740 39738 65796 39740
rect 65820 39738 65876 39740
rect 65900 39738 65956 39740
rect 65660 39686 65706 39738
rect 65706 39686 65716 39738
rect 65740 39686 65770 39738
rect 65770 39686 65782 39738
rect 65782 39686 65796 39738
rect 65820 39686 65834 39738
rect 65834 39686 65846 39738
rect 65846 39686 65876 39738
rect 65900 39686 65910 39738
rect 65910 39686 65956 39738
rect 65660 39684 65716 39686
rect 65740 39684 65796 39686
rect 65820 39684 65876 39686
rect 65900 39684 65956 39686
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 65660 38650 65716 38652
rect 65740 38650 65796 38652
rect 65820 38650 65876 38652
rect 65900 38650 65956 38652
rect 65660 38598 65706 38650
rect 65706 38598 65716 38650
rect 65740 38598 65770 38650
rect 65770 38598 65782 38650
rect 65782 38598 65796 38650
rect 65820 38598 65834 38650
rect 65834 38598 65846 38650
rect 65846 38598 65876 38650
rect 65900 38598 65910 38650
rect 65910 38598 65956 38650
rect 65660 38596 65716 38598
rect 65740 38596 65796 38598
rect 65820 38596 65876 38598
rect 65900 38596 65956 38598
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 65660 37562 65716 37564
rect 65740 37562 65796 37564
rect 65820 37562 65876 37564
rect 65900 37562 65956 37564
rect 65660 37510 65706 37562
rect 65706 37510 65716 37562
rect 65740 37510 65770 37562
rect 65770 37510 65782 37562
rect 65782 37510 65796 37562
rect 65820 37510 65834 37562
rect 65834 37510 65846 37562
rect 65846 37510 65876 37562
rect 65900 37510 65910 37562
rect 65910 37510 65956 37562
rect 65660 37508 65716 37510
rect 65740 37508 65796 37510
rect 65820 37508 65876 37510
rect 65900 37508 65956 37510
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 65660 36474 65716 36476
rect 65740 36474 65796 36476
rect 65820 36474 65876 36476
rect 65900 36474 65956 36476
rect 65660 36422 65706 36474
rect 65706 36422 65716 36474
rect 65740 36422 65770 36474
rect 65770 36422 65782 36474
rect 65782 36422 65796 36474
rect 65820 36422 65834 36474
rect 65834 36422 65846 36474
rect 65846 36422 65876 36474
rect 65900 36422 65910 36474
rect 65910 36422 65956 36474
rect 65660 36420 65716 36422
rect 65740 36420 65796 36422
rect 65820 36420 65876 36422
rect 65900 36420 65956 36422
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 14922 31084 14924 31104
rect 14924 31084 14976 31104
rect 14976 31084 14978 31104
rect 14922 31048 14978 31084
rect 11058 11056 11114 11112
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 8666 4140 8722 4176
rect 8666 4120 8668 4140
rect 8668 4120 8720 4140
rect 8720 4120 8722 4140
rect 10322 3884 10324 3904
rect 10324 3884 10376 3904
rect 10376 3884 10378 3904
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 10322 3848 10378 3884
rect 8390 3460 8446 3496
rect 8390 3440 8392 3460
rect 8392 3440 8444 3460
rect 8444 3440 8446 3460
rect 8482 3304 8538 3360
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10138 2760 10194 2816
rect 9954 2352 10010 2408
rect 10874 3032 10930 3088
rect 10966 1400 11022 1456
rect 16762 28600 16818 28656
rect 14186 20848 14242 20904
rect 14186 17484 14188 17504
rect 14188 17484 14240 17504
rect 14240 17484 14242 17504
rect 14186 17448 14242 17484
rect 13542 8336 13598 8392
rect 12254 5072 12310 5128
rect 12070 3476 12072 3496
rect 12072 3476 12124 3496
rect 12124 3476 12126 3496
rect 12070 3440 12126 3476
rect 12070 2932 12072 2952
rect 12072 2932 12124 2952
rect 12124 2932 12126 2952
rect 12070 2896 12126 2932
rect 11886 1944 11942 2000
rect 12806 4140 12862 4176
rect 12806 4120 12808 4140
rect 12808 4120 12860 4140
rect 12860 4120 12862 4140
rect 12714 2624 12770 2680
rect 13542 2488 13598 2544
rect 15014 20884 15016 20904
rect 15016 20884 15068 20904
rect 15068 20884 15070 20904
rect 15014 20848 15070 20884
rect 17038 28484 17094 28520
rect 17038 28464 17040 28484
rect 17040 28464 17092 28484
rect 17092 28464 17094 28484
rect 14922 13932 14978 13968
rect 14922 13912 14924 13932
rect 14924 13912 14976 13932
rect 14976 13912 14978 13932
rect 15198 6316 15254 6352
rect 15198 6296 15200 6316
rect 15200 6296 15252 6316
rect 15252 6296 15254 6316
rect 14922 5072 14978 5128
rect 13910 3304 13966 3360
rect 13910 2760 13966 2816
rect 14738 3984 14794 4040
rect 14462 2760 14518 2816
rect 14646 3848 14702 3904
rect 14646 2760 14702 2816
rect 14646 2644 14702 2680
rect 14646 2624 14648 2644
rect 14648 2624 14700 2644
rect 14700 2624 14702 2644
rect 14922 1944 14978 2000
rect 16486 17448 16542 17504
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 17038 17176 17094 17232
rect 18142 23432 18198 23488
rect 15290 3576 15346 3632
rect 15198 2916 15254 2952
rect 15198 2896 15200 2916
rect 15200 2896 15252 2916
rect 15252 2896 15254 2916
rect 15106 2624 15162 2680
rect 15198 2488 15254 2544
rect 15382 2372 15438 2408
rect 15382 2352 15384 2372
rect 15384 2352 15436 2372
rect 15436 2352 15438 2372
rect 16210 3032 16266 3088
rect 16026 2644 16082 2680
rect 16026 2624 16028 2644
rect 16028 2624 16080 2644
rect 16080 2624 16082 2644
rect 16486 3596 16542 3632
rect 16486 3576 16488 3596
rect 16488 3576 16540 3596
rect 16540 3576 16542 3596
rect 17038 1400 17094 1456
rect 17498 2524 17500 2544
rect 17500 2524 17552 2544
rect 17552 2524 17554 2544
rect 17498 2488 17554 2524
rect 18510 6160 18566 6216
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19430 25900 19486 25936
rect 19430 25880 19432 25900
rect 19432 25880 19484 25900
rect 19484 25880 19486 25900
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 20534 26968 20590 27024
rect 20442 25880 20498 25936
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19522 22616 19578 22672
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 22742 17040 22798 17096
rect 25134 22500 25190 22536
rect 25134 22480 25136 22500
rect 25136 22480 25188 22500
rect 25188 22480 25190 22500
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 27710 33516 27766 33552
rect 27710 33496 27712 33516
rect 27712 33496 27764 33516
rect 27764 33496 27766 33516
rect 28906 33532 28908 33552
rect 28908 33532 28960 33552
rect 28960 33532 28962 33552
rect 28906 33496 28962 33532
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 23478 17060 23534 17096
rect 23478 17040 23480 17060
rect 23480 17040 23532 17060
rect 23532 17040 23534 17060
rect 20810 8880 20866 8936
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 26330 13912 26386 13968
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 27250 6160 27306 6216
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 28722 6316 28778 6352
rect 28722 6296 28724 6316
rect 28724 6296 28776 6316
rect 28776 6296 28778 6316
rect 32770 22616 32826 22672
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 33506 17040 33562 17096
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 37830 28600 37886 28656
rect 42246 28500 42248 28520
rect 42248 28500 42300 28520
rect 42300 28500 42302 28520
rect 42246 28464 42302 28500
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 33598 8880 33654 8936
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 65660 35386 65716 35388
rect 65740 35386 65796 35388
rect 65820 35386 65876 35388
rect 65900 35386 65956 35388
rect 65660 35334 65706 35386
rect 65706 35334 65716 35386
rect 65740 35334 65770 35386
rect 65770 35334 65782 35386
rect 65782 35334 65796 35386
rect 65820 35334 65834 35386
rect 65834 35334 65846 35386
rect 65846 35334 65876 35386
rect 65900 35334 65910 35386
rect 65910 35334 65956 35386
rect 65660 35332 65716 35334
rect 65740 35332 65796 35334
rect 65820 35332 65876 35334
rect 65900 35332 65956 35334
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 65660 34298 65716 34300
rect 65740 34298 65796 34300
rect 65820 34298 65876 34300
rect 65900 34298 65956 34300
rect 65660 34246 65706 34298
rect 65706 34246 65716 34298
rect 65740 34246 65770 34298
rect 65770 34246 65782 34298
rect 65782 34246 65796 34298
rect 65820 34246 65834 34298
rect 65834 34246 65846 34298
rect 65846 34246 65876 34298
rect 65900 34246 65910 34298
rect 65910 34246 65956 34298
rect 65660 34244 65716 34246
rect 65740 34244 65796 34246
rect 65820 34244 65876 34246
rect 65900 34244 65956 34246
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 65660 33210 65716 33212
rect 65740 33210 65796 33212
rect 65820 33210 65876 33212
rect 65900 33210 65956 33212
rect 65660 33158 65706 33210
rect 65706 33158 65716 33210
rect 65740 33158 65770 33210
rect 65770 33158 65782 33210
rect 65782 33158 65796 33210
rect 65820 33158 65834 33210
rect 65834 33158 65846 33210
rect 65846 33158 65876 33210
rect 65900 33158 65910 33210
rect 65910 33158 65956 33210
rect 65660 33156 65716 33158
rect 65740 33156 65796 33158
rect 65820 33156 65876 33158
rect 65900 33156 65956 33158
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 65660 32122 65716 32124
rect 65740 32122 65796 32124
rect 65820 32122 65876 32124
rect 65900 32122 65956 32124
rect 65660 32070 65706 32122
rect 65706 32070 65716 32122
rect 65740 32070 65770 32122
rect 65770 32070 65782 32122
rect 65782 32070 65796 32122
rect 65820 32070 65834 32122
rect 65834 32070 65846 32122
rect 65846 32070 65876 32122
rect 65900 32070 65910 32122
rect 65910 32070 65956 32122
rect 65660 32068 65716 32070
rect 65740 32068 65796 32070
rect 65820 32068 65876 32070
rect 65900 32068 65956 32070
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 41970 22480 42026 22536
rect 42614 22480 42670 22536
rect 36174 11076 36230 11112
rect 36174 11056 36176 11076
rect 36176 11056 36228 11076
rect 36228 11056 36230 11076
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 38014 7520 38070 7576
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 33046 4528 33102 4584
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 38658 5228 38714 5264
rect 38658 5208 38660 5228
rect 38660 5208 38712 5228
rect 38712 5208 38714 5228
rect 38658 4256 38714 4312
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 39946 4256 40002 4312
rect 39854 3848 39910 3904
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 42614 7520 42670 7576
rect 40590 5208 40646 5264
rect 40866 4548 40922 4584
rect 40866 4528 40868 4548
rect 40868 4528 40920 4548
rect 40920 4528 40922 4548
rect 40590 3984 40646 4040
rect 42154 4528 42210 4584
rect 41878 4256 41934 4312
rect 42430 2352 42486 2408
rect 43350 3848 43406 3904
rect 42798 2372 42854 2408
rect 42798 2352 42800 2372
rect 42800 2352 42852 2372
rect 42852 2352 42854 2372
rect 43626 3440 43682 3496
rect 44270 3984 44326 4040
rect 43994 2896 44050 2952
rect 45282 2760 45338 2816
rect 47582 2916 47638 2952
rect 47582 2896 47584 2916
rect 47584 2896 47636 2916
rect 47636 2896 47638 2916
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 49882 9968 49938 10024
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50434 9968 50490 10024
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50986 9968 51042 10024
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 48870 3440 48926 3496
rect 48962 2760 49018 2816
rect 49238 2760 49294 2816
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 51906 2760 51962 2816
rect 65660 31034 65716 31036
rect 65740 31034 65796 31036
rect 65820 31034 65876 31036
rect 65900 31034 65956 31036
rect 65660 30982 65706 31034
rect 65706 30982 65716 31034
rect 65740 30982 65770 31034
rect 65770 30982 65782 31034
rect 65782 30982 65796 31034
rect 65820 30982 65834 31034
rect 65834 30982 65846 31034
rect 65846 30982 65876 31034
rect 65900 30982 65910 31034
rect 65910 30982 65956 31034
rect 65660 30980 65716 30982
rect 65740 30980 65796 30982
rect 65820 30980 65876 30982
rect 65900 30980 65956 30982
rect 65660 29946 65716 29948
rect 65740 29946 65796 29948
rect 65820 29946 65876 29948
rect 65900 29946 65956 29948
rect 65660 29894 65706 29946
rect 65706 29894 65716 29946
rect 65740 29894 65770 29946
rect 65770 29894 65782 29946
rect 65782 29894 65796 29946
rect 65820 29894 65834 29946
rect 65834 29894 65846 29946
rect 65846 29894 65876 29946
rect 65900 29894 65910 29946
rect 65910 29894 65956 29946
rect 65660 29892 65716 29894
rect 65740 29892 65796 29894
rect 65820 29892 65876 29894
rect 65900 29892 65956 29894
rect 53470 3460 53526 3496
rect 53470 3440 53472 3460
rect 53472 3440 53524 3460
rect 53524 3440 53526 3460
rect 65660 28858 65716 28860
rect 65740 28858 65796 28860
rect 65820 28858 65876 28860
rect 65900 28858 65956 28860
rect 65660 28806 65706 28858
rect 65706 28806 65716 28858
rect 65740 28806 65770 28858
rect 65770 28806 65782 28858
rect 65782 28806 65796 28858
rect 65820 28806 65834 28858
rect 65834 28806 65846 28858
rect 65846 28806 65876 28858
rect 65900 28806 65910 28858
rect 65910 28806 65956 28858
rect 65660 28804 65716 28806
rect 65740 28804 65796 28806
rect 65820 28804 65876 28806
rect 65900 28804 65956 28806
rect 67546 48612 67602 48648
rect 67546 48592 67548 48612
rect 67548 48592 67600 48612
rect 67600 48592 67602 48612
rect 68006 41112 68062 41168
rect 68006 33632 68062 33688
rect 65660 27770 65716 27772
rect 65740 27770 65796 27772
rect 65820 27770 65876 27772
rect 65900 27770 65956 27772
rect 65660 27718 65706 27770
rect 65706 27718 65716 27770
rect 65740 27718 65770 27770
rect 65770 27718 65782 27770
rect 65782 27718 65796 27770
rect 65820 27718 65834 27770
rect 65834 27718 65846 27770
rect 65846 27718 65876 27770
rect 65900 27718 65910 27770
rect 65910 27718 65956 27770
rect 65660 27716 65716 27718
rect 65740 27716 65796 27718
rect 65820 27716 65876 27718
rect 65900 27716 65956 27718
rect 65660 26682 65716 26684
rect 65740 26682 65796 26684
rect 65820 26682 65876 26684
rect 65900 26682 65956 26684
rect 65660 26630 65706 26682
rect 65706 26630 65716 26682
rect 65740 26630 65770 26682
rect 65770 26630 65782 26682
rect 65782 26630 65796 26682
rect 65820 26630 65834 26682
rect 65834 26630 65846 26682
rect 65846 26630 65876 26682
rect 65900 26630 65910 26682
rect 65910 26630 65956 26682
rect 65660 26628 65716 26630
rect 65740 26628 65796 26630
rect 65820 26628 65876 26630
rect 65900 26628 65956 26630
rect 65660 25594 65716 25596
rect 65740 25594 65796 25596
rect 65820 25594 65876 25596
rect 65900 25594 65956 25596
rect 65660 25542 65706 25594
rect 65706 25542 65716 25594
rect 65740 25542 65770 25594
rect 65770 25542 65782 25594
rect 65782 25542 65796 25594
rect 65820 25542 65834 25594
rect 65834 25542 65846 25594
rect 65846 25542 65876 25594
rect 65900 25542 65910 25594
rect 65910 25542 65956 25594
rect 65660 25540 65716 25542
rect 65740 25540 65796 25542
rect 65820 25540 65876 25542
rect 65900 25540 65956 25542
rect 68006 26152 68062 26208
rect 65660 24506 65716 24508
rect 65740 24506 65796 24508
rect 65820 24506 65876 24508
rect 65900 24506 65956 24508
rect 65660 24454 65706 24506
rect 65706 24454 65716 24506
rect 65740 24454 65770 24506
rect 65770 24454 65782 24506
rect 65782 24454 65796 24506
rect 65820 24454 65834 24506
rect 65834 24454 65846 24506
rect 65846 24454 65876 24506
rect 65900 24454 65910 24506
rect 65910 24454 65956 24506
rect 65660 24452 65716 24454
rect 65740 24452 65796 24454
rect 65820 24452 65876 24454
rect 65900 24452 65956 24454
rect 65660 23418 65716 23420
rect 65740 23418 65796 23420
rect 65820 23418 65876 23420
rect 65900 23418 65956 23420
rect 65660 23366 65706 23418
rect 65706 23366 65716 23418
rect 65740 23366 65770 23418
rect 65770 23366 65782 23418
rect 65782 23366 65796 23418
rect 65820 23366 65834 23418
rect 65834 23366 65846 23418
rect 65846 23366 65876 23418
rect 65900 23366 65910 23418
rect 65910 23366 65956 23418
rect 65660 23364 65716 23366
rect 65740 23364 65796 23366
rect 65820 23364 65876 23366
rect 65900 23364 65956 23366
rect 65660 22330 65716 22332
rect 65740 22330 65796 22332
rect 65820 22330 65876 22332
rect 65900 22330 65956 22332
rect 65660 22278 65706 22330
rect 65706 22278 65716 22330
rect 65740 22278 65770 22330
rect 65770 22278 65782 22330
rect 65782 22278 65796 22330
rect 65820 22278 65834 22330
rect 65834 22278 65846 22330
rect 65846 22278 65876 22330
rect 65900 22278 65910 22330
rect 65910 22278 65956 22330
rect 65660 22276 65716 22278
rect 65740 22276 65796 22278
rect 65820 22276 65876 22278
rect 65900 22276 65956 22278
rect 65660 21242 65716 21244
rect 65740 21242 65796 21244
rect 65820 21242 65876 21244
rect 65900 21242 65956 21244
rect 65660 21190 65706 21242
rect 65706 21190 65716 21242
rect 65740 21190 65770 21242
rect 65770 21190 65782 21242
rect 65782 21190 65796 21242
rect 65820 21190 65834 21242
rect 65834 21190 65846 21242
rect 65846 21190 65876 21242
rect 65900 21190 65910 21242
rect 65910 21190 65956 21242
rect 65660 21188 65716 21190
rect 65740 21188 65796 21190
rect 65820 21188 65876 21190
rect 65900 21188 65956 21190
rect 65660 20154 65716 20156
rect 65740 20154 65796 20156
rect 65820 20154 65876 20156
rect 65900 20154 65956 20156
rect 65660 20102 65706 20154
rect 65706 20102 65716 20154
rect 65740 20102 65770 20154
rect 65770 20102 65782 20154
rect 65782 20102 65796 20154
rect 65820 20102 65834 20154
rect 65834 20102 65846 20154
rect 65846 20102 65876 20154
rect 65900 20102 65910 20154
rect 65910 20102 65956 20154
rect 65660 20100 65716 20102
rect 65740 20100 65796 20102
rect 65820 20100 65876 20102
rect 65900 20100 65956 20102
rect 65660 19066 65716 19068
rect 65740 19066 65796 19068
rect 65820 19066 65876 19068
rect 65900 19066 65956 19068
rect 65660 19014 65706 19066
rect 65706 19014 65716 19066
rect 65740 19014 65770 19066
rect 65770 19014 65782 19066
rect 65782 19014 65796 19066
rect 65820 19014 65834 19066
rect 65834 19014 65846 19066
rect 65846 19014 65876 19066
rect 65900 19014 65910 19066
rect 65910 19014 65956 19066
rect 65660 19012 65716 19014
rect 65740 19012 65796 19014
rect 65820 19012 65876 19014
rect 65900 19012 65956 19014
rect 65660 17978 65716 17980
rect 65740 17978 65796 17980
rect 65820 17978 65876 17980
rect 65900 17978 65956 17980
rect 65660 17926 65706 17978
rect 65706 17926 65716 17978
rect 65740 17926 65770 17978
rect 65770 17926 65782 17978
rect 65782 17926 65796 17978
rect 65820 17926 65834 17978
rect 65834 17926 65846 17978
rect 65846 17926 65876 17978
rect 65900 17926 65910 17978
rect 65910 17926 65956 17978
rect 65660 17924 65716 17926
rect 65740 17924 65796 17926
rect 65820 17924 65876 17926
rect 65900 17924 65956 17926
rect 68006 18672 68062 18728
rect 65660 16890 65716 16892
rect 65740 16890 65796 16892
rect 65820 16890 65876 16892
rect 65900 16890 65956 16892
rect 65660 16838 65706 16890
rect 65706 16838 65716 16890
rect 65740 16838 65770 16890
rect 65770 16838 65782 16890
rect 65782 16838 65796 16890
rect 65820 16838 65834 16890
rect 65834 16838 65846 16890
rect 65846 16838 65876 16890
rect 65900 16838 65910 16890
rect 65910 16838 65956 16890
rect 65660 16836 65716 16838
rect 65740 16836 65796 16838
rect 65820 16836 65876 16838
rect 65900 16836 65956 16838
rect 65660 15802 65716 15804
rect 65740 15802 65796 15804
rect 65820 15802 65876 15804
rect 65900 15802 65956 15804
rect 65660 15750 65706 15802
rect 65706 15750 65716 15802
rect 65740 15750 65770 15802
rect 65770 15750 65782 15802
rect 65782 15750 65796 15802
rect 65820 15750 65834 15802
rect 65834 15750 65846 15802
rect 65846 15750 65876 15802
rect 65900 15750 65910 15802
rect 65910 15750 65956 15802
rect 65660 15748 65716 15750
rect 65740 15748 65796 15750
rect 65820 15748 65876 15750
rect 65900 15748 65956 15750
rect 65660 14714 65716 14716
rect 65740 14714 65796 14716
rect 65820 14714 65876 14716
rect 65900 14714 65956 14716
rect 65660 14662 65706 14714
rect 65706 14662 65716 14714
rect 65740 14662 65770 14714
rect 65770 14662 65782 14714
rect 65782 14662 65796 14714
rect 65820 14662 65834 14714
rect 65834 14662 65846 14714
rect 65846 14662 65876 14714
rect 65900 14662 65910 14714
rect 65910 14662 65956 14714
rect 65660 14660 65716 14662
rect 65740 14660 65796 14662
rect 65820 14660 65876 14662
rect 65900 14660 65956 14662
rect 65660 13626 65716 13628
rect 65740 13626 65796 13628
rect 65820 13626 65876 13628
rect 65900 13626 65956 13628
rect 65660 13574 65706 13626
rect 65706 13574 65716 13626
rect 65740 13574 65770 13626
rect 65770 13574 65782 13626
rect 65782 13574 65796 13626
rect 65820 13574 65834 13626
rect 65834 13574 65846 13626
rect 65846 13574 65876 13626
rect 65900 13574 65910 13626
rect 65910 13574 65956 13626
rect 65660 13572 65716 13574
rect 65740 13572 65796 13574
rect 65820 13572 65876 13574
rect 65900 13572 65956 13574
rect 65660 12538 65716 12540
rect 65740 12538 65796 12540
rect 65820 12538 65876 12540
rect 65900 12538 65956 12540
rect 65660 12486 65706 12538
rect 65706 12486 65716 12538
rect 65740 12486 65770 12538
rect 65770 12486 65782 12538
rect 65782 12486 65796 12538
rect 65820 12486 65834 12538
rect 65834 12486 65846 12538
rect 65846 12486 65876 12538
rect 65900 12486 65910 12538
rect 65910 12486 65956 12538
rect 65660 12484 65716 12486
rect 65740 12484 65796 12486
rect 65820 12484 65876 12486
rect 65900 12484 65956 12486
rect 65660 11450 65716 11452
rect 65740 11450 65796 11452
rect 65820 11450 65876 11452
rect 65900 11450 65956 11452
rect 65660 11398 65706 11450
rect 65706 11398 65716 11450
rect 65740 11398 65770 11450
rect 65770 11398 65782 11450
rect 65782 11398 65796 11450
rect 65820 11398 65834 11450
rect 65834 11398 65846 11450
rect 65846 11398 65876 11450
rect 65900 11398 65910 11450
rect 65910 11398 65956 11450
rect 65660 11396 65716 11398
rect 65740 11396 65796 11398
rect 65820 11396 65876 11398
rect 65900 11396 65956 11398
rect 67546 11192 67602 11248
rect 65660 10362 65716 10364
rect 65740 10362 65796 10364
rect 65820 10362 65876 10364
rect 65900 10362 65956 10364
rect 65660 10310 65706 10362
rect 65706 10310 65716 10362
rect 65740 10310 65770 10362
rect 65770 10310 65782 10362
rect 65782 10310 65796 10362
rect 65820 10310 65834 10362
rect 65834 10310 65846 10362
rect 65846 10310 65876 10362
rect 65900 10310 65910 10362
rect 65910 10310 65956 10362
rect 65660 10308 65716 10310
rect 65740 10308 65796 10310
rect 65820 10308 65876 10310
rect 65900 10308 65956 10310
rect 65660 9274 65716 9276
rect 65740 9274 65796 9276
rect 65820 9274 65876 9276
rect 65900 9274 65956 9276
rect 65660 9222 65706 9274
rect 65706 9222 65716 9274
rect 65740 9222 65770 9274
rect 65770 9222 65782 9274
rect 65782 9222 65796 9274
rect 65820 9222 65834 9274
rect 65834 9222 65846 9274
rect 65846 9222 65876 9274
rect 65900 9222 65910 9274
rect 65910 9222 65956 9274
rect 65660 9220 65716 9222
rect 65740 9220 65796 9222
rect 65820 9220 65876 9222
rect 65900 9220 65956 9222
rect 65660 8186 65716 8188
rect 65740 8186 65796 8188
rect 65820 8186 65876 8188
rect 65900 8186 65956 8188
rect 65660 8134 65706 8186
rect 65706 8134 65716 8186
rect 65740 8134 65770 8186
rect 65770 8134 65782 8186
rect 65782 8134 65796 8186
rect 65820 8134 65834 8186
rect 65834 8134 65846 8186
rect 65846 8134 65876 8186
rect 65900 8134 65910 8186
rect 65910 8134 65956 8186
rect 65660 8132 65716 8134
rect 65740 8132 65796 8134
rect 65820 8132 65876 8134
rect 65900 8132 65956 8134
rect 65660 7098 65716 7100
rect 65740 7098 65796 7100
rect 65820 7098 65876 7100
rect 65900 7098 65956 7100
rect 65660 7046 65706 7098
rect 65706 7046 65716 7098
rect 65740 7046 65770 7098
rect 65770 7046 65782 7098
rect 65782 7046 65796 7098
rect 65820 7046 65834 7098
rect 65834 7046 65846 7098
rect 65846 7046 65876 7098
rect 65900 7046 65910 7098
rect 65910 7046 65956 7098
rect 65660 7044 65716 7046
rect 65740 7044 65796 7046
rect 65820 7044 65876 7046
rect 65900 7044 65956 7046
rect 65660 6010 65716 6012
rect 65740 6010 65796 6012
rect 65820 6010 65876 6012
rect 65900 6010 65956 6012
rect 65660 5958 65706 6010
rect 65706 5958 65716 6010
rect 65740 5958 65770 6010
rect 65770 5958 65782 6010
rect 65782 5958 65796 6010
rect 65820 5958 65834 6010
rect 65834 5958 65846 6010
rect 65846 5958 65876 6010
rect 65900 5958 65910 6010
rect 65910 5958 65956 6010
rect 65660 5956 65716 5958
rect 65740 5956 65796 5958
rect 65820 5956 65876 5958
rect 65900 5956 65956 5958
rect 65660 4922 65716 4924
rect 65740 4922 65796 4924
rect 65820 4922 65876 4924
rect 65900 4922 65956 4924
rect 65660 4870 65706 4922
rect 65706 4870 65716 4922
rect 65740 4870 65770 4922
rect 65770 4870 65782 4922
rect 65782 4870 65796 4922
rect 65820 4870 65834 4922
rect 65834 4870 65846 4922
rect 65846 4870 65876 4922
rect 65900 4870 65910 4922
rect 65910 4870 65956 4922
rect 65660 4868 65716 4870
rect 65740 4868 65796 4870
rect 65820 4868 65876 4870
rect 65900 4868 65956 4870
rect 65660 3834 65716 3836
rect 65740 3834 65796 3836
rect 65820 3834 65876 3836
rect 65900 3834 65956 3836
rect 65660 3782 65706 3834
rect 65706 3782 65716 3834
rect 65740 3782 65770 3834
rect 65770 3782 65782 3834
rect 65782 3782 65796 3834
rect 65820 3782 65834 3834
rect 65834 3782 65846 3834
rect 65846 3782 65876 3834
rect 65900 3782 65910 3834
rect 65910 3782 65956 3834
rect 65660 3780 65716 3782
rect 65740 3780 65796 3782
rect 65820 3780 65876 3782
rect 65900 3780 65956 3782
rect 67546 3712 67602 3768
rect 65660 2746 65716 2748
rect 65740 2746 65796 2748
rect 65820 2746 65876 2748
rect 65900 2746 65956 2748
rect 65660 2694 65706 2746
rect 65706 2694 65716 2746
rect 65740 2694 65770 2746
rect 65770 2694 65782 2746
rect 65782 2694 65796 2746
rect 65820 2694 65834 2746
rect 65834 2694 65846 2746
rect 65846 2694 65876 2746
rect 65900 2694 65910 2746
rect 65910 2694 65956 2746
rect 65660 2692 65716 2694
rect 65740 2692 65796 2694
rect 65820 2692 65876 2694
rect 65900 2692 65956 2694
<< metal3 >>
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 65650 57152 65966 57153
rect 65650 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65966 57152
rect 65650 57087 65966 57088
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 67541 56130 67607 56133
rect 69200 56130 70000 56160
rect 67541 56128 70000 56130
rect 67541 56072 67546 56128
rect 67602 56072 70000 56128
rect 67541 56070 70000 56072
rect 67541 56067 67607 56070
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 65650 56064 65966 56065
rect 65650 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65966 56064
rect 69200 56040 70000 56070
rect 65650 55999 65966 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 65650 54976 65966 54977
rect 65650 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65966 54976
rect 65650 54911 65966 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 65650 53888 65966 53889
rect 65650 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65966 53888
rect 65650 53823 65966 53824
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 34930 52735 35246 52736
rect 65650 52800 65966 52801
rect 65650 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65966 52800
rect 65650 52735 65966 52736
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 65650 51712 65966 51713
rect 65650 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65966 51712
rect 65650 51647 65966 51648
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 65650 50624 65966 50625
rect 65650 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65966 50624
rect 65650 50559 65966 50560
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 34930 49471 35246 49472
rect 65650 49536 65966 49537
rect 65650 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65966 49536
rect 65650 49471 65966 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 67541 48650 67607 48653
rect 69200 48650 70000 48680
rect 67541 48648 70000 48650
rect 67541 48592 67546 48648
rect 67602 48592 70000 48648
rect 67541 48590 70000 48592
rect 67541 48587 67607 48590
rect 69200 48560 70000 48590
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 65650 48448 65966 48449
rect 65650 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65966 48448
rect 65650 48383 65966 48384
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 65650 47360 65966 47361
rect 65650 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65966 47360
rect 65650 47295 65966 47296
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 34930 46207 35246 46208
rect 65650 46272 65966 46273
rect 65650 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65966 46272
rect 65650 46207 65966 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 65650 45184 65966 45185
rect 65650 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65966 45184
rect 65650 45119 65966 45120
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 50290 44575 50606 44576
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 65650 44096 65966 44097
rect 65650 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65966 44096
rect 65650 44031 65966 44032
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 65650 43008 65966 43009
rect 65650 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65966 43008
rect 65650 42943 65966 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 65650 41920 65966 41921
rect 65650 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65966 41920
rect 65650 41855 65966 41856
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 50290 41311 50606 41312
rect 68001 41170 68067 41173
rect 69200 41170 70000 41200
rect 68001 41168 70000 41170
rect 68001 41112 68006 41168
rect 68062 41112 70000 41168
rect 68001 41110 70000 41112
rect 68001 41107 68067 41110
rect 69200 41080 70000 41110
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 65650 40832 65966 40833
rect 65650 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65966 40832
rect 65650 40767 65966 40768
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 65650 39744 65966 39745
rect 65650 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65966 39744
rect 65650 39679 65966 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 65650 38656 65966 38657
rect 65650 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65966 38656
rect 65650 38591 65966 38592
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 65650 37568 65966 37569
rect 65650 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65966 37568
rect 65650 37503 65966 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 65650 36480 65966 36481
rect 65650 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65966 36480
rect 65650 36415 65966 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 65650 35392 65966 35393
rect 65650 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65966 35392
rect 65650 35327 65966 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 65650 34304 65966 34305
rect 65650 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65966 34304
rect 65650 34239 65966 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 68001 33690 68067 33693
rect 69200 33690 70000 33720
rect 68001 33688 70000 33690
rect 68001 33632 68006 33688
rect 68062 33632 70000 33688
rect 68001 33630 70000 33632
rect 68001 33627 68067 33630
rect 69200 33600 70000 33630
rect 27705 33554 27771 33557
rect 28901 33554 28967 33557
rect 27705 33552 28967 33554
rect 27705 33496 27710 33552
rect 27766 33496 28906 33552
rect 28962 33496 28967 33552
rect 27705 33494 28967 33496
rect 27705 33491 27771 33494
rect 28901 33491 28967 33494
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 65650 33216 65966 33217
rect 65650 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65966 33216
rect 65650 33151 65966 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 65650 32128 65966 32129
rect 65650 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65966 32128
rect 65650 32063 65966 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 50290 31519 50606 31520
rect 14917 31108 14983 31109
rect 14917 31106 14964 31108
rect 14872 31104 14964 31106
rect 14872 31048 14922 31104
rect 14872 31046 14964 31048
rect 14917 31044 14964 31046
rect 15028 31044 15034 31108
rect 14917 31043 14983 31044
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 65650 31040 65966 31041
rect 65650 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65966 31040
rect 65650 30975 65966 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 65650 29952 65966 29953
rect 65650 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65966 29952
rect 65650 29887 65966 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 65650 28864 65966 28865
rect 65650 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65966 28864
rect 65650 28799 65966 28800
rect 16757 28658 16823 28661
rect 37825 28658 37891 28661
rect 16757 28656 37891 28658
rect 16757 28600 16762 28656
rect 16818 28600 37830 28656
rect 37886 28600 37891 28656
rect 16757 28598 37891 28600
rect 16757 28595 16823 28598
rect 37825 28595 37891 28598
rect 17033 28522 17099 28525
rect 42241 28522 42307 28525
rect 17033 28520 42307 28522
rect 17033 28464 17038 28520
rect 17094 28464 42246 28520
rect 42302 28464 42307 28520
rect 17033 28462 42307 28464
rect 17033 28459 17099 28462
rect 42241 28459 42307 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 50290 28255 50606 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 65650 27776 65966 27777
rect 65650 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65966 27776
rect 65650 27711 65966 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 19374 26964 19380 27028
rect 19444 27026 19450 27028
rect 20529 27026 20595 27029
rect 19444 27024 20595 27026
rect 19444 26968 20534 27024
rect 20590 26968 20595 27024
rect 19444 26966 20595 26968
rect 19444 26964 19450 26966
rect 20529 26963 20595 26966
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 65650 26688 65966 26689
rect 65650 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65966 26688
rect 65650 26623 65966 26624
rect 68001 26210 68067 26213
rect 69200 26210 70000 26240
rect 68001 26208 70000 26210
rect 68001 26152 68006 26208
rect 68062 26152 70000 26208
rect 68001 26150 70000 26152
rect 68001 26147 68067 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 69200 26120 70000 26150
rect 50290 26079 50606 26080
rect 19425 25938 19491 25941
rect 20437 25938 20503 25941
rect 19425 25936 20503 25938
rect 19425 25880 19430 25936
rect 19486 25880 20442 25936
rect 20498 25880 20503 25936
rect 19425 25878 20503 25880
rect 19425 25875 19491 25878
rect 20437 25875 20503 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 65650 25600 65966 25601
rect 65650 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65966 25600
rect 65650 25535 65966 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 65650 24512 65966 24513
rect 65650 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65966 24512
rect 65650 24447 65966 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 18137 23490 18203 23493
rect 19374 23490 19380 23492
rect 18137 23488 19380 23490
rect 18137 23432 18142 23488
rect 18198 23432 19380 23488
rect 18137 23430 19380 23432
rect 18137 23427 18203 23430
rect 19374 23428 19380 23430
rect 19444 23428 19450 23492
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 65650 23424 65966 23425
rect 65650 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65966 23424
rect 65650 23359 65966 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 19517 22674 19583 22677
rect 32765 22674 32831 22677
rect 19517 22672 32831 22674
rect 19517 22616 19522 22672
rect 19578 22616 32770 22672
rect 32826 22616 32831 22672
rect 19517 22614 32831 22616
rect 19517 22611 19583 22614
rect 32765 22611 32831 22614
rect 25129 22538 25195 22541
rect 41965 22538 42031 22541
rect 42609 22538 42675 22541
rect 25129 22536 42675 22538
rect 25129 22480 25134 22536
rect 25190 22480 41970 22536
rect 42026 22480 42614 22536
rect 42670 22480 42675 22536
rect 25129 22478 42675 22480
rect 25129 22475 25195 22478
rect 41965 22475 42031 22478
rect 42609 22475 42675 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 65650 22336 65966 22337
rect 65650 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65966 22336
rect 65650 22271 65966 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 65650 21248 65966 21249
rect 65650 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65966 21248
rect 65650 21183 65966 21184
rect 14181 20906 14247 20909
rect 14590 20906 14596 20908
rect 14181 20904 14596 20906
rect 14181 20848 14186 20904
rect 14242 20848 14596 20904
rect 14181 20846 14596 20848
rect 14181 20843 14247 20846
rect 14590 20844 14596 20846
rect 14660 20906 14666 20908
rect 15009 20906 15075 20909
rect 14660 20904 15075 20906
rect 14660 20848 15014 20904
rect 15070 20848 15075 20904
rect 14660 20846 15075 20848
rect 14660 20844 14666 20846
rect 15009 20843 15075 20846
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 65650 20160 65966 20161
rect 65650 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65966 20160
rect 65650 20095 65966 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 65650 19072 65966 19073
rect 65650 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65966 19072
rect 65650 19007 65966 19008
rect 68001 18730 68067 18733
rect 69200 18730 70000 18760
rect 68001 18728 70000 18730
rect 68001 18672 68006 18728
rect 68062 18672 70000 18728
rect 68001 18670 70000 18672
rect 68001 18667 68067 18670
rect 69200 18640 70000 18670
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 50290 18463 50606 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 65650 17984 65966 17985
rect 65650 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65966 17984
rect 65650 17919 65966 17920
rect 14181 17506 14247 17509
rect 15694 17506 15700 17508
rect 14181 17504 15700 17506
rect 14181 17448 14186 17504
rect 14242 17448 15700 17504
rect 14181 17446 15700 17448
rect 14181 17443 14247 17446
rect 15694 17444 15700 17446
rect 15764 17506 15770 17508
rect 16481 17506 16547 17509
rect 15764 17504 16547 17506
rect 15764 17448 16486 17504
rect 16542 17448 16547 17504
rect 15764 17446 16547 17448
rect 15764 17444 15770 17446
rect 16481 17443 16547 17446
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 16062 17172 16068 17236
rect 16132 17234 16138 17236
rect 17033 17234 17099 17237
rect 16132 17232 17099 17234
rect 16132 17176 17038 17232
rect 17094 17176 17099 17232
rect 16132 17174 17099 17176
rect 16132 17172 16138 17174
rect 17033 17171 17099 17174
rect 14038 17036 14044 17100
rect 14108 17098 14114 17100
rect 22737 17098 22803 17101
rect 14108 17096 22803 17098
rect 14108 17040 22742 17096
rect 22798 17040 22803 17096
rect 14108 17038 22803 17040
rect 14108 17036 14114 17038
rect 22737 17035 22803 17038
rect 23473 17098 23539 17101
rect 33501 17098 33567 17101
rect 23473 17096 33567 17098
rect 23473 17040 23478 17096
rect 23534 17040 33506 17096
rect 33562 17040 33567 17096
rect 23473 17038 33567 17040
rect 23473 17035 23539 17038
rect 33501 17035 33567 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 65650 16896 65966 16897
rect 65650 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65966 16896
rect 65650 16831 65966 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 65650 15808 65966 15809
rect 65650 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65966 15808
rect 65650 15743 65966 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 65650 14720 65966 14721
rect 65650 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65966 14720
rect 65650 14655 65966 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 14917 13970 14983 13973
rect 26325 13970 26391 13973
rect 14917 13968 26391 13970
rect 14917 13912 14922 13968
rect 14978 13912 26330 13968
rect 26386 13912 26391 13968
rect 14917 13910 26391 13912
rect 14917 13907 14983 13910
rect 26325 13907 26391 13910
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 65650 13632 65966 13633
rect 65650 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65966 13632
rect 65650 13567 65966 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 65650 12544 65966 12545
rect 65650 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65966 12544
rect 65650 12479 65966 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 50290 11935 50606 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 65650 11456 65966 11457
rect 65650 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65966 11456
rect 65650 11391 65966 11392
rect 67541 11250 67607 11253
rect 69200 11250 70000 11280
rect 67541 11248 70000 11250
rect 67541 11192 67546 11248
rect 67602 11192 70000 11248
rect 67541 11190 70000 11192
rect 67541 11187 67607 11190
rect 69200 11160 70000 11190
rect 11053 11114 11119 11117
rect 36169 11114 36235 11117
rect 11053 11112 36235 11114
rect 11053 11056 11058 11112
rect 11114 11056 36174 11112
rect 36230 11056 36235 11112
rect 11053 11054 36235 11056
rect 11053 11051 11119 11054
rect 36169 11051 36235 11054
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 65650 10368 65966 10369
rect 65650 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65966 10368
rect 65650 10303 65966 10304
rect 49877 10026 49943 10029
rect 50429 10026 50495 10029
rect 50981 10026 51047 10029
rect 49877 10024 51047 10026
rect 49877 9968 49882 10024
rect 49938 9968 50434 10024
rect 50490 9968 50986 10024
rect 51042 9968 51047 10024
rect 49877 9966 51047 9968
rect 49877 9963 49943 9966
rect 50429 9963 50495 9966
rect 50981 9963 51047 9966
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 65650 9280 65966 9281
rect 65650 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65966 9280
rect 65650 9215 65966 9216
rect 20805 8938 20871 8941
rect 33593 8938 33659 8941
rect 20805 8936 33659 8938
rect 20805 8880 20810 8936
rect 20866 8880 33598 8936
rect 33654 8880 33659 8936
rect 20805 8878 33659 8880
rect 20805 8875 20871 8878
rect 33593 8875 33659 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 50290 8671 50606 8672
rect 13537 8394 13603 8397
rect 13854 8394 13860 8396
rect 13537 8392 13860 8394
rect 13537 8336 13542 8392
rect 13598 8336 13860 8392
rect 13537 8334 13860 8336
rect 13537 8331 13603 8334
rect 13854 8332 13860 8334
rect 13924 8332 13930 8396
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 65650 8192 65966 8193
rect 65650 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65966 8192
rect 65650 8127 65966 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 38009 7578 38075 7581
rect 42609 7578 42675 7581
rect 38009 7576 42675 7578
rect 38009 7520 38014 7576
rect 38070 7520 42614 7576
rect 42670 7520 42675 7576
rect 38009 7518 42675 7520
rect 38009 7515 38075 7518
rect 42609 7515 42675 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 65650 7104 65966 7105
rect 65650 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65966 7104
rect 65650 7039 65966 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 15193 6354 15259 6357
rect 28717 6354 28783 6357
rect 15193 6352 28783 6354
rect 15193 6296 15198 6352
rect 15254 6296 28722 6352
rect 28778 6296 28783 6352
rect 15193 6294 28783 6296
rect 15193 6291 15259 6294
rect 28717 6291 28783 6294
rect 18505 6218 18571 6221
rect 27245 6218 27311 6221
rect 18505 6216 27311 6218
rect 18505 6160 18510 6216
rect 18566 6160 27250 6216
rect 27306 6160 27311 6216
rect 18505 6158 27311 6160
rect 18505 6155 18571 6158
rect 27245 6155 27311 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 65650 6016 65966 6017
rect 65650 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65966 6016
rect 65650 5951 65966 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 38653 5266 38719 5269
rect 40585 5266 40651 5269
rect 38653 5264 40651 5266
rect 38653 5208 38658 5264
rect 38714 5208 40590 5264
rect 40646 5208 40651 5264
rect 38653 5206 40651 5208
rect 38653 5203 38719 5206
rect 40585 5203 40651 5206
rect 12249 5130 12315 5133
rect 14917 5130 14983 5133
rect 12249 5128 14983 5130
rect 12249 5072 12254 5128
rect 12310 5072 14922 5128
rect 14978 5072 14983 5128
rect 12249 5070 14983 5072
rect 12249 5067 12315 5070
rect 14917 5067 14983 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 65650 4928 65966 4929
rect 65650 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65966 4928
rect 65650 4863 65966 4864
rect 33041 4586 33107 4589
rect 40861 4586 40927 4589
rect 42149 4586 42215 4589
rect 33041 4584 42215 4586
rect 33041 4528 33046 4584
rect 33102 4528 40866 4584
rect 40922 4528 42154 4584
rect 42210 4528 42215 4584
rect 33041 4526 42215 4528
rect 33041 4523 33107 4526
rect 40861 4523 40927 4526
rect 42149 4523 42215 4526
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 38653 4314 38719 4317
rect 39941 4314 40007 4317
rect 41873 4314 41939 4317
rect 38653 4312 41939 4314
rect 38653 4256 38658 4312
rect 38714 4256 39946 4312
rect 40002 4256 41878 4312
rect 41934 4256 41939 4312
rect 38653 4254 41939 4256
rect 38653 4251 38719 4254
rect 39941 4251 40007 4254
rect 41873 4251 41939 4254
rect 8661 4178 8727 4181
rect 12801 4178 12867 4181
rect 8661 4176 12867 4178
rect 8661 4120 8666 4176
rect 8722 4120 12806 4176
rect 12862 4120 12867 4176
rect 8661 4118 12867 4120
rect 8661 4115 8727 4118
rect 12801 4115 12867 4118
rect 13854 3980 13860 4044
rect 13924 4042 13930 4044
rect 14733 4042 14799 4045
rect 13924 4040 14799 4042
rect 13924 3984 14738 4040
rect 14794 3984 14799 4040
rect 13924 3982 14799 3984
rect 13924 3980 13930 3982
rect 14733 3979 14799 3982
rect 40585 4042 40651 4045
rect 44265 4042 44331 4045
rect 40585 4040 44331 4042
rect 40585 3984 40590 4040
rect 40646 3984 44270 4040
rect 44326 3984 44331 4040
rect 40585 3982 44331 3984
rect 40585 3979 40651 3982
rect 44265 3979 44331 3982
rect 10317 3906 10383 3909
rect 14641 3906 14707 3909
rect 10317 3904 14707 3906
rect 10317 3848 10322 3904
rect 10378 3848 14646 3904
rect 14702 3848 14707 3904
rect 10317 3846 14707 3848
rect 10317 3843 10383 3846
rect 14641 3843 14707 3846
rect 39849 3906 39915 3909
rect 43345 3906 43411 3909
rect 39849 3904 43411 3906
rect 39849 3848 39854 3904
rect 39910 3848 43350 3904
rect 43406 3848 43411 3904
rect 39849 3846 43411 3848
rect 39849 3843 39915 3846
rect 43345 3843 43411 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 65650 3840 65966 3841
rect 65650 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65966 3840
rect 65650 3775 65966 3776
rect 67541 3770 67607 3773
rect 69200 3770 70000 3800
rect 67541 3768 70000 3770
rect 67541 3712 67546 3768
rect 67602 3712 70000 3768
rect 67541 3710 70000 3712
rect 67541 3707 67607 3710
rect 69200 3680 70000 3710
rect 15285 3634 15351 3637
rect 16481 3634 16547 3637
rect 15285 3632 16547 3634
rect 15285 3576 15290 3632
rect 15346 3576 16486 3632
rect 16542 3576 16547 3632
rect 15285 3574 16547 3576
rect 15285 3571 15351 3574
rect 16481 3571 16547 3574
rect 8385 3498 8451 3501
rect 12065 3498 12131 3501
rect 8385 3496 12131 3498
rect 8385 3440 8390 3496
rect 8446 3440 12070 3496
rect 12126 3440 12131 3496
rect 8385 3438 12131 3440
rect 8385 3435 8451 3438
rect 12065 3435 12131 3438
rect 43621 3498 43687 3501
rect 48865 3498 48931 3501
rect 53465 3498 53531 3501
rect 43621 3496 53531 3498
rect 43621 3440 43626 3496
rect 43682 3440 48870 3496
rect 48926 3440 53470 3496
rect 53526 3440 53531 3496
rect 43621 3438 53531 3440
rect 43621 3435 43687 3438
rect 48865 3435 48931 3438
rect 53465 3435 53531 3438
rect 8477 3362 8543 3365
rect 13905 3362 13971 3365
rect 14038 3362 14044 3364
rect 8477 3360 14044 3362
rect 8477 3304 8482 3360
rect 8538 3304 13910 3360
rect 13966 3304 14044 3360
rect 8477 3302 14044 3304
rect 8477 3299 8543 3302
rect 13905 3299 13971 3302
rect 14038 3300 14044 3302
rect 14108 3300 14114 3364
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 10869 3090 10935 3093
rect 16205 3090 16271 3093
rect 10869 3088 16271 3090
rect 10869 3032 10874 3088
rect 10930 3032 16210 3088
rect 16266 3032 16271 3088
rect 10869 3030 16271 3032
rect 10869 3027 10935 3030
rect 16205 3027 16271 3030
rect 12065 2954 12131 2957
rect 15193 2954 15259 2957
rect 12065 2952 15259 2954
rect 12065 2896 12070 2952
rect 12126 2896 15198 2952
rect 15254 2896 15259 2952
rect 12065 2894 15259 2896
rect 12065 2891 12131 2894
rect 15193 2891 15259 2894
rect 43989 2954 44055 2957
rect 47577 2954 47643 2957
rect 43989 2952 47643 2954
rect 43989 2896 43994 2952
rect 44050 2896 47582 2952
rect 47638 2896 47643 2952
rect 43989 2894 47643 2896
rect 43989 2891 44055 2894
rect 47577 2891 47643 2894
rect 10133 2818 10199 2821
rect 13905 2818 13971 2821
rect 10133 2816 13971 2818
rect 10133 2760 10138 2816
rect 10194 2760 13910 2816
rect 13966 2760 13971 2816
rect 10133 2758 13971 2760
rect 10133 2755 10199 2758
rect 13905 2755 13971 2758
rect 14038 2756 14044 2820
rect 14108 2756 14114 2820
rect 14457 2818 14523 2821
rect 14641 2818 14707 2821
rect 14457 2816 14707 2818
rect 14457 2760 14462 2816
rect 14518 2760 14646 2816
rect 14702 2760 14707 2816
rect 14457 2758 14707 2760
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 12709 2682 12775 2685
rect 14046 2682 14106 2756
rect 14457 2755 14523 2758
rect 14641 2755 14707 2758
rect 45277 2818 45343 2821
rect 48957 2818 49023 2821
rect 45277 2816 49023 2818
rect 45277 2760 45282 2816
rect 45338 2760 48962 2816
rect 49018 2760 49023 2816
rect 45277 2758 49023 2760
rect 45277 2755 45343 2758
rect 48957 2755 49023 2758
rect 49233 2818 49299 2821
rect 51901 2818 51967 2821
rect 49233 2816 51967 2818
rect 49233 2760 49238 2816
rect 49294 2760 51906 2816
rect 51962 2760 51967 2816
rect 49233 2758 51967 2760
rect 49233 2755 49299 2758
rect 51901 2755 51967 2758
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 65650 2752 65966 2753
rect 65650 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65966 2752
rect 65650 2687 65966 2688
rect 14641 2684 14707 2685
rect 12709 2680 14106 2682
rect 12709 2624 12714 2680
rect 12770 2624 14106 2680
rect 12709 2622 14106 2624
rect 12709 2619 12775 2622
rect 14590 2620 14596 2684
rect 14660 2682 14707 2684
rect 14660 2680 14752 2682
rect 14702 2624 14752 2680
rect 14660 2622 14752 2624
rect 14660 2620 14707 2622
rect 14958 2620 14964 2684
rect 15028 2682 15034 2684
rect 15101 2682 15167 2685
rect 16021 2684 16087 2685
rect 16021 2682 16068 2684
rect 15028 2680 15167 2682
rect 15028 2624 15106 2680
rect 15162 2624 15167 2680
rect 15028 2622 15167 2624
rect 15976 2680 16068 2682
rect 15976 2624 16026 2680
rect 15976 2622 16068 2624
rect 15028 2620 15034 2622
rect 14641 2619 14707 2620
rect 15101 2619 15167 2622
rect 16021 2620 16068 2622
rect 16132 2620 16138 2684
rect 16021 2619 16087 2620
rect 13537 2546 13603 2549
rect 15193 2546 15259 2549
rect 13537 2544 15259 2546
rect 13537 2488 13542 2544
rect 13598 2488 15198 2544
rect 15254 2488 15259 2544
rect 13537 2486 15259 2488
rect 13537 2483 13603 2486
rect 15193 2483 15259 2486
rect 15694 2484 15700 2548
rect 15764 2546 15770 2548
rect 17493 2546 17559 2549
rect 15764 2544 17559 2546
rect 15764 2488 17498 2544
rect 17554 2488 17559 2544
rect 15764 2486 17559 2488
rect 15764 2484 15770 2486
rect 17493 2483 17559 2486
rect 9949 2410 10015 2413
rect 15377 2410 15443 2413
rect 9949 2408 15443 2410
rect 9949 2352 9954 2408
rect 10010 2352 15382 2408
rect 15438 2352 15443 2408
rect 9949 2350 15443 2352
rect 9949 2347 10015 2350
rect 15377 2347 15443 2350
rect 42425 2410 42491 2413
rect 42793 2410 42859 2413
rect 42425 2408 42859 2410
rect 42425 2352 42430 2408
rect 42486 2352 42798 2408
rect 42854 2352 42859 2408
rect 42425 2350 42859 2352
rect 42425 2347 42491 2350
rect 42793 2347 42859 2350
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
rect 11881 2002 11947 2005
rect 14917 2002 14983 2005
rect 11881 2000 14983 2002
rect 11881 1944 11886 2000
rect 11942 1944 14922 2000
rect 14978 1944 14983 2000
rect 11881 1942 14983 1944
rect 11881 1939 11947 1942
rect 14917 1939 14983 1942
rect 10961 1458 11027 1461
rect 17033 1458 17099 1461
rect 10961 1456 17099 1458
rect 10961 1400 10966 1456
rect 11022 1400 17038 1456
rect 17094 1400 17099 1456
rect 10961 1398 17099 1400
rect 10961 1395 11027 1398
rect 17033 1395 17099 1398
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 65656 57148 65720 57152
rect 65656 57092 65660 57148
rect 65660 57092 65716 57148
rect 65716 57092 65720 57148
rect 65656 57088 65720 57092
rect 65736 57148 65800 57152
rect 65736 57092 65740 57148
rect 65740 57092 65796 57148
rect 65796 57092 65800 57148
rect 65736 57088 65800 57092
rect 65816 57148 65880 57152
rect 65816 57092 65820 57148
rect 65820 57092 65876 57148
rect 65876 57092 65880 57148
rect 65816 57088 65880 57092
rect 65896 57148 65960 57152
rect 65896 57092 65900 57148
rect 65900 57092 65956 57148
rect 65956 57092 65960 57148
rect 65896 57088 65960 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 65656 56060 65720 56064
rect 65656 56004 65660 56060
rect 65660 56004 65716 56060
rect 65716 56004 65720 56060
rect 65656 56000 65720 56004
rect 65736 56060 65800 56064
rect 65736 56004 65740 56060
rect 65740 56004 65796 56060
rect 65796 56004 65800 56060
rect 65736 56000 65800 56004
rect 65816 56060 65880 56064
rect 65816 56004 65820 56060
rect 65820 56004 65876 56060
rect 65876 56004 65880 56060
rect 65816 56000 65880 56004
rect 65896 56060 65960 56064
rect 65896 56004 65900 56060
rect 65900 56004 65956 56060
rect 65956 56004 65960 56060
rect 65896 56000 65960 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 65656 54972 65720 54976
rect 65656 54916 65660 54972
rect 65660 54916 65716 54972
rect 65716 54916 65720 54972
rect 65656 54912 65720 54916
rect 65736 54972 65800 54976
rect 65736 54916 65740 54972
rect 65740 54916 65796 54972
rect 65796 54916 65800 54972
rect 65736 54912 65800 54916
rect 65816 54972 65880 54976
rect 65816 54916 65820 54972
rect 65820 54916 65876 54972
rect 65876 54916 65880 54972
rect 65816 54912 65880 54916
rect 65896 54972 65960 54976
rect 65896 54916 65900 54972
rect 65900 54916 65956 54972
rect 65956 54916 65960 54972
rect 65896 54912 65960 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 65656 53884 65720 53888
rect 65656 53828 65660 53884
rect 65660 53828 65716 53884
rect 65716 53828 65720 53884
rect 65656 53824 65720 53828
rect 65736 53884 65800 53888
rect 65736 53828 65740 53884
rect 65740 53828 65796 53884
rect 65796 53828 65800 53884
rect 65736 53824 65800 53828
rect 65816 53884 65880 53888
rect 65816 53828 65820 53884
rect 65820 53828 65876 53884
rect 65876 53828 65880 53884
rect 65816 53824 65880 53828
rect 65896 53884 65960 53888
rect 65896 53828 65900 53884
rect 65900 53828 65956 53884
rect 65956 53828 65960 53884
rect 65896 53824 65960 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 65656 52796 65720 52800
rect 65656 52740 65660 52796
rect 65660 52740 65716 52796
rect 65716 52740 65720 52796
rect 65656 52736 65720 52740
rect 65736 52796 65800 52800
rect 65736 52740 65740 52796
rect 65740 52740 65796 52796
rect 65796 52740 65800 52796
rect 65736 52736 65800 52740
rect 65816 52796 65880 52800
rect 65816 52740 65820 52796
rect 65820 52740 65876 52796
rect 65876 52740 65880 52796
rect 65816 52736 65880 52740
rect 65896 52796 65960 52800
rect 65896 52740 65900 52796
rect 65900 52740 65956 52796
rect 65956 52740 65960 52796
rect 65896 52736 65960 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 65656 51708 65720 51712
rect 65656 51652 65660 51708
rect 65660 51652 65716 51708
rect 65716 51652 65720 51708
rect 65656 51648 65720 51652
rect 65736 51708 65800 51712
rect 65736 51652 65740 51708
rect 65740 51652 65796 51708
rect 65796 51652 65800 51708
rect 65736 51648 65800 51652
rect 65816 51708 65880 51712
rect 65816 51652 65820 51708
rect 65820 51652 65876 51708
rect 65876 51652 65880 51708
rect 65816 51648 65880 51652
rect 65896 51708 65960 51712
rect 65896 51652 65900 51708
rect 65900 51652 65956 51708
rect 65956 51652 65960 51708
rect 65896 51648 65960 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 65656 50620 65720 50624
rect 65656 50564 65660 50620
rect 65660 50564 65716 50620
rect 65716 50564 65720 50620
rect 65656 50560 65720 50564
rect 65736 50620 65800 50624
rect 65736 50564 65740 50620
rect 65740 50564 65796 50620
rect 65796 50564 65800 50620
rect 65736 50560 65800 50564
rect 65816 50620 65880 50624
rect 65816 50564 65820 50620
rect 65820 50564 65876 50620
rect 65876 50564 65880 50620
rect 65816 50560 65880 50564
rect 65896 50620 65960 50624
rect 65896 50564 65900 50620
rect 65900 50564 65956 50620
rect 65956 50564 65960 50620
rect 65896 50560 65960 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 65656 49532 65720 49536
rect 65656 49476 65660 49532
rect 65660 49476 65716 49532
rect 65716 49476 65720 49532
rect 65656 49472 65720 49476
rect 65736 49532 65800 49536
rect 65736 49476 65740 49532
rect 65740 49476 65796 49532
rect 65796 49476 65800 49532
rect 65736 49472 65800 49476
rect 65816 49532 65880 49536
rect 65816 49476 65820 49532
rect 65820 49476 65876 49532
rect 65876 49476 65880 49532
rect 65816 49472 65880 49476
rect 65896 49532 65960 49536
rect 65896 49476 65900 49532
rect 65900 49476 65956 49532
rect 65956 49476 65960 49532
rect 65896 49472 65960 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 65656 48444 65720 48448
rect 65656 48388 65660 48444
rect 65660 48388 65716 48444
rect 65716 48388 65720 48444
rect 65656 48384 65720 48388
rect 65736 48444 65800 48448
rect 65736 48388 65740 48444
rect 65740 48388 65796 48444
rect 65796 48388 65800 48444
rect 65736 48384 65800 48388
rect 65816 48444 65880 48448
rect 65816 48388 65820 48444
rect 65820 48388 65876 48444
rect 65876 48388 65880 48444
rect 65816 48384 65880 48388
rect 65896 48444 65960 48448
rect 65896 48388 65900 48444
rect 65900 48388 65956 48444
rect 65956 48388 65960 48444
rect 65896 48384 65960 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 65656 47356 65720 47360
rect 65656 47300 65660 47356
rect 65660 47300 65716 47356
rect 65716 47300 65720 47356
rect 65656 47296 65720 47300
rect 65736 47356 65800 47360
rect 65736 47300 65740 47356
rect 65740 47300 65796 47356
rect 65796 47300 65800 47356
rect 65736 47296 65800 47300
rect 65816 47356 65880 47360
rect 65816 47300 65820 47356
rect 65820 47300 65876 47356
rect 65876 47300 65880 47356
rect 65816 47296 65880 47300
rect 65896 47356 65960 47360
rect 65896 47300 65900 47356
rect 65900 47300 65956 47356
rect 65956 47300 65960 47356
rect 65896 47296 65960 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 65656 46268 65720 46272
rect 65656 46212 65660 46268
rect 65660 46212 65716 46268
rect 65716 46212 65720 46268
rect 65656 46208 65720 46212
rect 65736 46268 65800 46272
rect 65736 46212 65740 46268
rect 65740 46212 65796 46268
rect 65796 46212 65800 46268
rect 65736 46208 65800 46212
rect 65816 46268 65880 46272
rect 65816 46212 65820 46268
rect 65820 46212 65876 46268
rect 65876 46212 65880 46268
rect 65816 46208 65880 46212
rect 65896 46268 65960 46272
rect 65896 46212 65900 46268
rect 65900 46212 65956 46268
rect 65956 46212 65960 46268
rect 65896 46208 65960 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 65656 45180 65720 45184
rect 65656 45124 65660 45180
rect 65660 45124 65716 45180
rect 65716 45124 65720 45180
rect 65656 45120 65720 45124
rect 65736 45180 65800 45184
rect 65736 45124 65740 45180
rect 65740 45124 65796 45180
rect 65796 45124 65800 45180
rect 65736 45120 65800 45124
rect 65816 45180 65880 45184
rect 65816 45124 65820 45180
rect 65820 45124 65876 45180
rect 65876 45124 65880 45180
rect 65816 45120 65880 45124
rect 65896 45180 65960 45184
rect 65896 45124 65900 45180
rect 65900 45124 65956 45180
rect 65956 45124 65960 45180
rect 65896 45120 65960 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 65656 44092 65720 44096
rect 65656 44036 65660 44092
rect 65660 44036 65716 44092
rect 65716 44036 65720 44092
rect 65656 44032 65720 44036
rect 65736 44092 65800 44096
rect 65736 44036 65740 44092
rect 65740 44036 65796 44092
rect 65796 44036 65800 44092
rect 65736 44032 65800 44036
rect 65816 44092 65880 44096
rect 65816 44036 65820 44092
rect 65820 44036 65876 44092
rect 65876 44036 65880 44092
rect 65816 44032 65880 44036
rect 65896 44092 65960 44096
rect 65896 44036 65900 44092
rect 65900 44036 65956 44092
rect 65956 44036 65960 44092
rect 65896 44032 65960 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 65656 43004 65720 43008
rect 65656 42948 65660 43004
rect 65660 42948 65716 43004
rect 65716 42948 65720 43004
rect 65656 42944 65720 42948
rect 65736 43004 65800 43008
rect 65736 42948 65740 43004
rect 65740 42948 65796 43004
rect 65796 42948 65800 43004
rect 65736 42944 65800 42948
rect 65816 43004 65880 43008
rect 65816 42948 65820 43004
rect 65820 42948 65876 43004
rect 65876 42948 65880 43004
rect 65816 42944 65880 42948
rect 65896 43004 65960 43008
rect 65896 42948 65900 43004
rect 65900 42948 65956 43004
rect 65956 42948 65960 43004
rect 65896 42944 65960 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 65656 41916 65720 41920
rect 65656 41860 65660 41916
rect 65660 41860 65716 41916
rect 65716 41860 65720 41916
rect 65656 41856 65720 41860
rect 65736 41916 65800 41920
rect 65736 41860 65740 41916
rect 65740 41860 65796 41916
rect 65796 41860 65800 41916
rect 65736 41856 65800 41860
rect 65816 41916 65880 41920
rect 65816 41860 65820 41916
rect 65820 41860 65876 41916
rect 65876 41860 65880 41916
rect 65816 41856 65880 41860
rect 65896 41916 65960 41920
rect 65896 41860 65900 41916
rect 65900 41860 65956 41916
rect 65956 41860 65960 41916
rect 65896 41856 65960 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 65656 40828 65720 40832
rect 65656 40772 65660 40828
rect 65660 40772 65716 40828
rect 65716 40772 65720 40828
rect 65656 40768 65720 40772
rect 65736 40828 65800 40832
rect 65736 40772 65740 40828
rect 65740 40772 65796 40828
rect 65796 40772 65800 40828
rect 65736 40768 65800 40772
rect 65816 40828 65880 40832
rect 65816 40772 65820 40828
rect 65820 40772 65876 40828
rect 65876 40772 65880 40828
rect 65816 40768 65880 40772
rect 65896 40828 65960 40832
rect 65896 40772 65900 40828
rect 65900 40772 65956 40828
rect 65956 40772 65960 40828
rect 65896 40768 65960 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 65656 39740 65720 39744
rect 65656 39684 65660 39740
rect 65660 39684 65716 39740
rect 65716 39684 65720 39740
rect 65656 39680 65720 39684
rect 65736 39740 65800 39744
rect 65736 39684 65740 39740
rect 65740 39684 65796 39740
rect 65796 39684 65800 39740
rect 65736 39680 65800 39684
rect 65816 39740 65880 39744
rect 65816 39684 65820 39740
rect 65820 39684 65876 39740
rect 65876 39684 65880 39740
rect 65816 39680 65880 39684
rect 65896 39740 65960 39744
rect 65896 39684 65900 39740
rect 65900 39684 65956 39740
rect 65956 39684 65960 39740
rect 65896 39680 65960 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 65656 38652 65720 38656
rect 65656 38596 65660 38652
rect 65660 38596 65716 38652
rect 65716 38596 65720 38652
rect 65656 38592 65720 38596
rect 65736 38652 65800 38656
rect 65736 38596 65740 38652
rect 65740 38596 65796 38652
rect 65796 38596 65800 38652
rect 65736 38592 65800 38596
rect 65816 38652 65880 38656
rect 65816 38596 65820 38652
rect 65820 38596 65876 38652
rect 65876 38596 65880 38652
rect 65816 38592 65880 38596
rect 65896 38652 65960 38656
rect 65896 38596 65900 38652
rect 65900 38596 65956 38652
rect 65956 38596 65960 38652
rect 65896 38592 65960 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 65656 37564 65720 37568
rect 65656 37508 65660 37564
rect 65660 37508 65716 37564
rect 65716 37508 65720 37564
rect 65656 37504 65720 37508
rect 65736 37564 65800 37568
rect 65736 37508 65740 37564
rect 65740 37508 65796 37564
rect 65796 37508 65800 37564
rect 65736 37504 65800 37508
rect 65816 37564 65880 37568
rect 65816 37508 65820 37564
rect 65820 37508 65876 37564
rect 65876 37508 65880 37564
rect 65816 37504 65880 37508
rect 65896 37564 65960 37568
rect 65896 37508 65900 37564
rect 65900 37508 65956 37564
rect 65956 37508 65960 37564
rect 65896 37504 65960 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 65656 36476 65720 36480
rect 65656 36420 65660 36476
rect 65660 36420 65716 36476
rect 65716 36420 65720 36476
rect 65656 36416 65720 36420
rect 65736 36476 65800 36480
rect 65736 36420 65740 36476
rect 65740 36420 65796 36476
rect 65796 36420 65800 36476
rect 65736 36416 65800 36420
rect 65816 36476 65880 36480
rect 65816 36420 65820 36476
rect 65820 36420 65876 36476
rect 65876 36420 65880 36476
rect 65816 36416 65880 36420
rect 65896 36476 65960 36480
rect 65896 36420 65900 36476
rect 65900 36420 65956 36476
rect 65956 36420 65960 36476
rect 65896 36416 65960 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 65656 35388 65720 35392
rect 65656 35332 65660 35388
rect 65660 35332 65716 35388
rect 65716 35332 65720 35388
rect 65656 35328 65720 35332
rect 65736 35388 65800 35392
rect 65736 35332 65740 35388
rect 65740 35332 65796 35388
rect 65796 35332 65800 35388
rect 65736 35328 65800 35332
rect 65816 35388 65880 35392
rect 65816 35332 65820 35388
rect 65820 35332 65876 35388
rect 65876 35332 65880 35388
rect 65816 35328 65880 35332
rect 65896 35388 65960 35392
rect 65896 35332 65900 35388
rect 65900 35332 65956 35388
rect 65956 35332 65960 35388
rect 65896 35328 65960 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 65656 34300 65720 34304
rect 65656 34244 65660 34300
rect 65660 34244 65716 34300
rect 65716 34244 65720 34300
rect 65656 34240 65720 34244
rect 65736 34300 65800 34304
rect 65736 34244 65740 34300
rect 65740 34244 65796 34300
rect 65796 34244 65800 34300
rect 65736 34240 65800 34244
rect 65816 34300 65880 34304
rect 65816 34244 65820 34300
rect 65820 34244 65876 34300
rect 65876 34244 65880 34300
rect 65816 34240 65880 34244
rect 65896 34300 65960 34304
rect 65896 34244 65900 34300
rect 65900 34244 65956 34300
rect 65956 34244 65960 34300
rect 65896 34240 65960 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 65656 33212 65720 33216
rect 65656 33156 65660 33212
rect 65660 33156 65716 33212
rect 65716 33156 65720 33212
rect 65656 33152 65720 33156
rect 65736 33212 65800 33216
rect 65736 33156 65740 33212
rect 65740 33156 65796 33212
rect 65796 33156 65800 33212
rect 65736 33152 65800 33156
rect 65816 33212 65880 33216
rect 65816 33156 65820 33212
rect 65820 33156 65876 33212
rect 65876 33156 65880 33212
rect 65816 33152 65880 33156
rect 65896 33212 65960 33216
rect 65896 33156 65900 33212
rect 65900 33156 65956 33212
rect 65956 33156 65960 33212
rect 65896 33152 65960 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 65656 32124 65720 32128
rect 65656 32068 65660 32124
rect 65660 32068 65716 32124
rect 65716 32068 65720 32124
rect 65656 32064 65720 32068
rect 65736 32124 65800 32128
rect 65736 32068 65740 32124
rect 65740 32068 65796 32124
rect 65796 32068 65800 32124
rect 65736 32064 65800 32068
rect 65816 32124 65880 32128
rect 65816 32068 65820 32124
rect 65820 32068 65876 32124
rect 65876 32068 65880 32124
rect 65816 32064 65880 32068
rect 65896 32124 65960 32128
rect 65896 32068 65900 32124
rect 65900 32068 65956 32124
rect 65956 32068 65960 32124
rect 65896 32064 65960 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 14964 31104 15028 31108
rect 14964 31048 14978 31104
rect 14978 31048 15028 31104
rect 14964 31044 15028 31048
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 65656 31036 65720 31040
rect 65656 30980 65660 31036
rect 65660 30980 65716 31036
rect 65716 30980 65720 31036
rect 65656 30976 65720 30980
rect 65736 31036 65800 31040
rect 65736 30980 65740 31036
rect 65740 30980 65796 31036
rect 65796 30980 65800 31036
rect 65736 30976 65800 30980
rect 65816 31036 65880 31040
rect 65816 30980 65820 31036
rect 65820 30980 65876 31036
rect 65876 30980 65880 31036
rect 65816 30976 65880 30980
rect 65896 31036 65960 31040
rect 65896 30980 65900 31036
rect 65900 30980 65956 31036
rect 65956 30980 65960 31036
rect 65896 30976 65960 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 65656 29948 65720 29952
rect 65656 29892 65660 29948
rect 65660 29892 65716 29948
rect 65716 29892 65720 29948
rect 65656 29888 65720 29892
rect 65736 29948 65800 29952
rect 65736 29892 65740 29948
rect 65740 29892 65796 29948
rect 65796 29892 65800 29948
rect 65736 29888 65800 29892
rect 65816 29948 65880 29952
rect 65816 29892 65820 29948
rect 65820 29892 65876 29948
rect 65876 29892 65880 29948
rect 65816 29888 65880 29892
rect 65896 29948 65960 29952
rect 65896 29892 65900 29948
rect 65900 29892 65956 29948
rect 65956 29892 65960 29948
rect 65896 29888 65960 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 65656 28860 65720 28864
rect 65656 28804 65660 28860
rect 65660 28804 65716 28860
rect 65716 28804 65720 28860
rect 65656 28800 65720 28804
rect 65736 28860 65800 28864
rect 65736 28804 65740 28860
rect 65740 28804 65796 28860
rect 65796 28804 65800 28860
rect 65736 28800 65800 28804
rect 65816 28860 65880 28864
rect 65816 28804 65820 28860
rect 65820 28804 65876 28860
rect 65876 28804 65880 28860
rect 65816 28800 65880 28804
rect 65896 28860 65960 28864
rect 65896 28804 65900 28860
rect 65900 28804 65956 28860
rect 65956 28804 65960 28860
rect 65896 28800 65960 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 65656 27772 65720 27776
rect 65656 27716 65660 27772
rect 65660 27716 65716 27772
rect 65716 27716 65720 27772
rect 65656 27712 65720 27716
rect 65736 27772 65800 27776
rect 65736 27716 65740 27772
rect 65740 27716 65796 27772
rect 65796 27716 65800 27772
rect 65736 27712 65800 27716
rect 65816 27772 65880 27776
rect 65816 27716 65820 27772
rect 65820 27716 65876 27772
rect 65876 27716 65880 27772
rect 65816 27712 65880 27716
rect 65896 27772 65960 27776
rect 65896 27716 65900 27772
rect 65900 27716 65956 27772
rect 65956 27716 65960 27772
rect 65896 27712 65960 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 19380 26964 19444 27028
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 65656 26684 65720 26688
rect 65656 26628 65660 26684
rect 65660 26628 65716 26684
rect 65716 26628 65720 26684
rect 65656 26624 65720 26628
rect 65736 26684 65800 26688
rect 65736 26628 65740 26684
rect 65740 26628 65796 26684
rect 65796 26628 65800 26684
rect 65736 26624 65800 26628
rect 65816 26684 65880 26688
rect 65816 26628 65820 26684
rect 65820 26628 65876 26684
rect 65876 26628 65880 26684
rect 65816 26624 65880 26628
rect 65896 26684 65960 26688
rect 65896 26628 65900 26684
rect 65900 26628 65956 26684
rect 65956 26628 65960 26684
rect 65896 26624 65960 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 65656 25596 65720 25600
rect 65656 25540 65660 25596
rect 65660 25540 65716 25596
rect 65716 25540 65720 25596
rect 65656 25536 65720 25540
rect 65736 25596 65800 25600
rect 65736 25540 65740 25596
rect 65740 25540 65796 25596
rect 65796 25540 65800 25596
rect 65736 25536 65800 25540
rect 65816 25596 65880 25600
rect 65816 25540 65820 25596
rect 65820 25540 65876 25596
rect 65876 25540 65880 25596
rect 65816 25536 65880 25540
rect 65896 25596 65960 25600
rect 65896 25540 65900 25596
rect 65900 25540 65956 25596
rect 65956 25540 65960 25596
rect 65896 25536 65960 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 65656 24508 65720 24512
rect 65656 24452 65660 24508
rect 65660 24452 65716 24508
rect 65716 24452 65720 24508
rect 65656 24448 65720 24452
rect 65736 24508 65800 24512
rect 65736 24452 65740 24508
rect 65740 24452 65796 24508
rect 65796 24452 65800 24508
rect 65736 24448 65800 24452
rect 65816 24508 65880 24512
rect 65816 24452 65820 24508
rect 65820 24452 65876 24508
rect 65876 24452 65880 24508
rect 65816 24448 65880 24452
rect 65896 24508 65960 24512
rect 65896 24452 65900 24508
rect 65900 24452 65956 24508
rect 65956 24452 65960 24508
rect 65896 24448 65960 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 19380 23428 19444 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 65656 23420 65720 23424
rect 65656 23364 65660 23420
rect 65660 23364 65716 23420
rect 65716 23364 65720 23420
rect 65656 23360 65720 23364
rect 65736 23420 65800 23424
rect 65736 23364 65740 23420
rect 65740 23364 65796 23420
rect 65796 23364 65800 23420
rect 65736 23360 65800 23364
rect 65816 23420 65880 23424
rect 65816 23364 65820 23420
rect 65820 23364 65876 23420
rect 65876 23364 65880 23420
rect 65816 23360 65880 23364
rect 65896 23420 65960 23424
rect 65896 23364 65900 23420
rect 65900 23364 65956 23420
rect 65956 23364 65960 23420
rect 65896 23360 65960 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 65656 22332 65720 22336
rect 65656 22276 65660 22332
rect 65660 22276 65716 22332
rect 65716 22276 65720 22332
rect 65656 22272 65720 22276
rect 65736 22332 65800 22336
rect 65736 22276 65740 22332
rect 65740 22276 65796 22332
rect 65796 22276 65800 22332
rect 65736 22272 65800 22276
rect 65816 22332 65880 22336
rect 65816 22276 65820 22332
rect 65820 22276 65876 22332
rect 65876 22276 65880 22332
rect 65816 22272 65880 22276
rect 65896 22332 65960 22336
rect 65896 22276 65900 22332
rect 65900 22276 65956 22332
rect 65956 22276 65960 22332
rect 65896 22272 65960 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 65656 21244 65720 21248
rect 65656 21188 65660 21244
rect 65660 21188 65716 21244
rect 65716 21188 65720 21244
rect 65656 21184 65720 21188
rect 65736 21244 65800 21248
rect 65736 21188 65740 21244
rect 65740 21188 65796 21244
rect 65796 21188 65800 21244
rect 65736 21184 65800 21188
rect 65816 21244 65880 21248
rect 65816 21188 65820 21244
rect 65820 21188 65876 21244
rect 65876 21188 65880 21244
rect 65816 21184 65880 21188
rect 65896 21244 65960 21248
rect 65896 21188 65900 21244
rect 65900 21188 65956 21244
rect 65956 21188 65960 21244
rect 65896 21184 65960 21188
rect 14596 20844 14660 20908
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 65656 20156 65720 20160
rect 65656 20100 65660 20156
rect 65660 20100 65716 20156
rect 65716 20100 65720 20156
rect 65656 20096 65720 20100
rect 65736 20156 65800 20160
rect 65736 20100 65740 20156
rect 65740 20100 65796 20156
rect 65796 20100 65800 20156
rect 65736 20096 65800 20100
rect 65816 20156 65880 20160
rect 65816 20100 65820 20156
rect 65820 20100 65876 20156
rect 65876 20100 65880 20156
rect 65816 20096 65880 20100
rect 65896 20156 65960 20160
rect 65896 20100 65900 20156
rect 65900 20100 65956 20156
rect 65956 20100 65960 20156
rect 65896 20096 65960 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 65656 19068 65720 19072
rect 65656 19012 65660 19068
rect 65660 19012 65716 19068
rect 65716 19012 65720 19068
rect 65656 19008 65720 19012
rect 65736 19068 65800 19072
rect 65736 19012 65740 19068
rect 65740 19012 65796 19068
rect 65796 19012 65800 19068
rect 65736 19008 65800 19012
rect 65816 19068 65880 19072
rect 65816 19012 65820 19068
rect 65820 19012 65876 19068
rect 65876 19012 65880 19068
rect 65816 19008 65880 19012
rect 65896 19068 65960 19072
rect 65896 19012 65900 19068
rect 65900 19012 65956 19068
rect 65956 19012 65960 19068
rect 65896 19008 65960 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 65656 17980 65720 17984
rect 65656 17924 65660 17980
rect 65660 17924 65716 17980
rect 65716 17924 65720 17980
rect 65656 17920 65720 17924
rect 65736 17980 65800 17984
rect 65736 17924 65740 17980
rect 65740 17924 65796 17980
rect 65796 17924 65800 17980
rect 65736 17920 65800 17924
rect 65816 17980 65880 17984
rect 65816 17924 65820 17980
rect 65820 17924 65876 17980
rect 65876 17924 65880 17980
rect 65816 17920 65880 17924
rect 65896 17980 65960 17984
rect 65896 17924 65900 17980
rect 65900 17924 65956 17980
rect 65956 17924 65960 17980
rect 65896 17920 65960 17924
rect 15700 17444 15764 17508
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 16068 17172 16132 17236
rect 14044 17036 14108 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 65656 16892 65720 16896
rect 65656 16836 65660 16892
rect 65660 16836 65716 16892
rect 65716 16836 65720 16892
rect 65656 16832 65720 16836
rect 65736 16892 65800 16896
rect 65736 16836 65740 16892
rect 65740 16836 65796 16892
rect 65796 16836 65800 16892
rect 65736 16832 65800 16836
rect 65816 16892 65880 16896
rect 65816 16836 65820 16892
rect 65820 16836 65876 16892
rect 65876 16836 65880 16892
rect 65816 16832 65880 16836
rect 65896 16892 65960 16896
rect 65896 16836 65900 16892
rect 65900 16836 65956 16892
rect 65956 16836 65960 16892
rect 65896 16832 65960 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 65656 15804 65720 15808
rect 65656 15748 65660 15804
rect 65660 15748 65716 15804
rect 65716 15748 65720 15804
rect 65656 15744 65720 15748
rect 65736 15804 65800 15808
rect 65736 15748 65740 15804
rect 65740 15748 65796 15804
rect 65796 15748 65800 15804
rect 65736 15744 65800 15748
rect 65816 15804 65880 15808
rect 65816 15748 65820 15804
rect 65820 15748 65876 15804
rect 65876 15748 65880 15804
rect 65816 15744 65880 15748
rect 65896 15804 65960 15808
rect 65896 15748 65900 15804
rect 65900 15748 65956 15804
rect 65956 15748 65960 15804
rect 65896 15744 65960 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 65656 14716 65720 14720
rect 65656 14660 65660 14716
rect 65660 14660 65716 14716
rect 65716 14660 65720 14716
rect 65656 14656 65720 14660
rect 65736 14716 65800 14720
rect 65736 14660 65740 14716
rect 65740 14660 65796 14716
rect 65796 14660 65800 14716
rect 65736 14656 65800 14660
rect 65816 14716 65880 14720
rect 65816 14660 65820 14716
rect 65820 14660 65876 14716
rect 65876 14660 65880 14716
rect 65816 14656 65880 14660
rect 65896 14716 65960 14720
rect 65896 14660 65900 14716
rect 65900 14660 65956 14716
rect 65956 14660 65960 14716
rect 65896 14656 65960 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 65656 13628 65720 13632
rect 65656 13572 65660 13628
rect 65660 13572 65716 13628
rect 65716 13572 65720 13628
rect 65656 13568 65720 13572
rect 65736 13628 65800 13632
rect 65736 13572 65740 13628
rect 65740 13572 65796 13628
rect 65796 13572 65800 13628
rect 65736 13568 65800 13572
rect 65816 13628 65880 13632
rect 65816 13572 65820 13628
rect 65820 13572 65876 13628
rect 65876 13572 65880 13628
rect 65816 13568 65880 13572
rect 65896 13628 65960 13632
rect 65896 13572 65900 13628
rect 65900 13572 65956 13628
rect 65956 13572 65960 13628
rect 65896 13568 65960 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 65656 12540 65720 12544
rect 65656 12484 65660 12540
rect 65660 12484 65716 12540
rect 65716 12484 65720 12540
rect 65656 12480 65720 12484
rect 65736 12540 65800 12544
rect 65736 12484 65740 12540
rect 65740 12484 65796 12540
rect 65796 12484 65800 12540
rect 65736 12480 65800 12484
rect 65816 12540 65880 12544
rect 65816 12484 65820 12540
rect 65820 12484 65876 12540
rect 65876 12484 65880 12540
rect 65816 12480 65880 12484
rect 65896 12540 65960 12544
rect 65896 12484 65900 12540
rect 65900 12484 65956 12540
rect 65956 12484 65960 12540
rect 65896 12480 65960 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 65656 11452 65720 11456
rect 65656 11396 65660 11452
rect 65660 11396 65716 11452
rect 65716 11396 65720 11452
rect 65656 11392 65720 11396
rect 65736 11452 65800 11456
rect 65736 11396 65740 11452
rect 65740 11396 65796 11452
rect 65796 11396 65800 11452
rect 65736 11392 65800 11396
rect 65816 11452 65880 11456
rect 65816 11396 65820 11452
rect 65820 11396 65876 11452
rect 65876 11396 65880 11452
rect 65816 11392 65880 11396
rect 65896 11452 65960 11456
rect 65896 11396 65900 11452
rect 65900 11396 65956 11452
rect 65956 11396 65960 11452
rect 65896 11392 65960 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 65656 10364 65720 10368
rect 65656 10308 65660 10364
rect 65660 10308 65716 10364
rect 65716 10308 65720 10364
rect 65656 10304 65720 10308
rect 65736 10364 65800 10368
rect 65736 10308 65740 10364
rect 65740 10308 65796 10364
rect 65796 10308 65800 10364
rect 65736 10304 65800 10308
rect 65816 10364 65880 10368
rect 65816 10308 65820 10364
rect 65820 10308 65876 10364
rect 65876 10308 65880 10364
rect 65816 10304 65880 10308
rect 65896 10364 65960 10368
rect 65896 10308 65900 10364
rect 65900 10308 65956 10364
rect 65956 10308 65960 10364
rect 65896 10304 65960 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 65656 9276 65720 9280
rect 65656 9220 65660 9276
rect 65660 9220 65716 9276
rect 65716 9220 65720 9276
rect 65656 9216 65720 9220
rect 65736 9276 65800 9280
rect 65736 9220 65740 9276
rect 65740 9220 65796 9276
rect 65796 9220 65800 9276
rect 65736 9216 65800 9220
rect 65816 9276 65880 9280
rect 65816 9220 65820 9276
rect 65820 9220 65876 9276
rect 65876 9220 65880 9276
rect 65816 9216 65880 9220
rect 65896 9276 65960 9280
rect 65896 9220 65900 9276
rect 65900 9220 65956 9276
rect 65956 9220 65960 9276
rect 65896 9216 65960 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 13860 8332 13924 8396
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 65656 8188 65720 8192
rect 65656 8132 65660 8188
rect 65660 8132 65716 8188
rect 65716 8132 65720 8188
rect 65656 8128 65720 8132
rect 65736 8188 65800 8192
rect 65736 8132 65740 8188
rect 65740 8132 65796 8188
rect 65796 8132 65800 8188
rect 65736 8128 65800 8132
rect 65816 8188 65880 8192
rect 65816 8132 65820 8188
rect 65820 8132 65876 8188
rect 65876 8132 65880 8188
rect 65816 8128 65880 8132
rect 65896 8188 65960 8192
rect 65896 8132 65900 8188
rect 65900 8132 65956 8188
rect 65956 8132 65960 8188
rect 65896 8128 65960 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 65656 7100 65720 7104
rect 65656 7044 65660 7100
rect 65660 7044 65716 7100
rect 65716 7044 65720 7100
rect 65656 7040 65720 7044
rect 65736 7100 65800 7104
rect 65736 7044 65740 7100
rect 65740 7044 65796 7100
rect 65796 7044 65800 7100
rect 65736 7040 65800 7044
rect 65816 7100 65880 7104
rect 65816 7044 65820 7100
rect 65820 7044 65876 7100
rect 65876 7044 65880 7100
rect 65816 7040 65880 7044
rect 65896 7100 65960 7104
rect 65896 7044 65900 7100
rect 65900 7044 65956 7100
rect 65956 7044 65960 7100
rect 65896 7040 65960 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 65656 6012 65720 6016
rect 65656 5956 65660 6012
rect 65660 5956 65716 6012
rect 65716 5956 65720 6012
rect 65656 5952 65720 5956
rect 65736 6012 65800 6016
rect 65736 5956 65740 6012
rect 65740 5956 65796 6012
rect 65796 5956 65800 6012
rect 65736 5952 65800 5956
rect 65816 6012 65880 6016
rect 65816 5956 65820 6012
rect 65820 5956 65876 6012
rect 65876 5956 65880 6012
rect 65816 5952 65880 5956
rect 65896 6012 65960 6016
rect 65896 5956 65900 6012
rect 65900 5956 65956 6012
rect 65956 5956 65960 6012
rect 65896 5952 65960 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 65656 4924 65720 4928
rect 65656 4868 65660 4924
rect 65660 4868 65716 4924
rect 65716 4868 65720 4924
rect 65656 4864 65720 4868
rect 65736 4924 65800 4928
rect 65736 4868 65740 4924
rect 65740 4868 65796 4924
rect 65796 4868 65800 4924
rect 65736 4864 65800 4868
rect 65816 4924 65880 4928
rect 65816 4868 65820 4924
rect 65820 4868 65876 4924
rect 65876 4868 65880 4924
rect 65816 4864 65880 4868
rect 65896 4924 65960 4928
rect 65896 4868 65900 4924
rect 65900 4868 65956 4924
rect 65956 4868 65960 4924
rect 65896 4864 65960 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 13860 3980 13924 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 65656 3836 65720 3840
rect 65656 3780 65660 3836
rect 65660 3780 65716 3836
rect 65716 3780 65720 3836
rect 65656 3776 65720 3780
rect 65736 3836 65800 3840
rect 65736 3780 65740 3836
rect 65740 3780 65796 3836
rect 65796 3780 65800 3836
rect 65736 3776 65800 3780
rect 65816 3836 65880 3840
rect 65816 3780 65820 3836
rect 65820 3780 65876 3836
rect 65876 3780 65880 3836
rect 65816 3776 65880 3780
rect 65896 3836 65960 3840
rect 65896 3780 65900 3836
rect 65900 3780 65956 3836
rect 65956 3780 65960 3836
rect 65896 3776 65960 3780
rect 14044 3300 14108 3364
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 14044 2756 14108 2820
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 65656 2748 65720 2752
rect 65656 2692 65660 2748
rect 65660 2692 65716 2748
rect 65716 2692 65720 2748
rect 65656 2688 65720 2692
rect 65736 2748 65800 2752
rect 65736 2692 65740 2748
rect 65740 2692 65796 2748
rect 65796 2692 65800 2748
rect 65736 2688 65800 2692
rect 65816 2748 65880 2752
rect 65816 2692 65820 2748
rect 65820 2692 65876 2748
rect 65876 2692 65880 2748
rect 65816 2688 65880 2692
rect 65896 2748 65960 2752
rect 65896 2692 65900 2748
rect 65900 2692 65956 2748
rect 65956 2692 65960 2748
rect 65896 2688 65960 2692
rect 14596 2680 14660 2684
rect 14596 2624 14646 2680
rect 14646 2624 14660 2680
rect 14596 2620 14660 2624
rect 14964 2620 15028 2684
rect 16068 2680 16132 2684
rect 16068 2624 16082 2680
rect 16082 2624 16132 2680
rect 16068 2620 16132 2624
rect 15700 2484 15764 2548
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 14963 31108 15029 31109
rect 14963 31044 14964 31108
rect 15028 31044 15029 31108
rect 14963 31043 15029 31044
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 14595 20908 14661 20909
rect 14595 20844 14596 20908
rect 14660 20844 14661 20908
rect 14595 20843 14661 20844
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 14043 17100 14109 17101
rect 14043 17036 14044 17100
rect 14108 17036 14109 17100
rect 14043 17035 14109 17036
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 13859 8396 13925 8397
rect 13859 8332 13860 8396
rect 13924 8332 13925 8396
rect 13859 8331 13925 8332
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 13862 4045 13922 8331
rect 13859 4044 13925 4045
rect 13859 3980 13860 4044
rect 13924 3980 13925 4044
rect 13859 3979 13925 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 14046 3365 14106 17035
rect 14043 3364 14109 3365
rect 14043 3300 14044 3364
rect 14108 3300 14109 3364
rect 14043 3299 14109 3300
rect 14046 2821 14106 3299
rect 14043 2820 14109 2821
rect 14043 2756 14044 2820
rect 14108 2756 14109 2820
rect 14043 2755 14109 2756
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 14598 2685 14658 20843
rect 14966 2685 15026 31043
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19379 27028 19445 27029
rect 19379 26964 19380 27028
rect 19444 26964 19445 27028
rect 19379 26963 19445 26964
rect 19382 23493 19442 26963
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19379 23492 19445 23493
rect 19379 23428 19380 23492
rect 19444 23428 19445 23492
rect 19379 23427 19445 23428
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 15699 17508 15765 17509
rect 15699 17444 15700 17508
rect 15764 17444 15765 17508
rect 15699 17443 15765 17444
rect 14595 2684 14661 2685
rect 14595 2620 14596 2684
rect 14660 2620 14661 2684
rect 14595 2619 14661 2620
rect 14963 2684 15029 2685
rect 14963 2620 14964 2684
rect 15028 2620 15029 2684
rect 14963 2619 15029 2620
rect 15702 2549 15762 17443
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 16067 17236 16133 17237
rect 16067 17172 16068 17236
rect 16132 17172 16133 17236
rect 16067 17171 16133 17172
rect 16070 2685 16130 17171
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 16067 2684 16133 2685
rect 16067 2620 16068 2684
rect 16132 2620 16133 2684
rect 16067 2619 16133 2620
rect 15699 2548 15765 2549
rect 15699 2484 15700 2548
rect 15764 2484 15765 2548
rect 15699 2483 15765 2484
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
rect 65648 57152 65968 57712
rect 65648 57088 65656 57152
rect 65720 57088 65736 57152
rect 65800 57088 65816 57152
rect 65880 57088 65896 57152
rect 65960 57088 65968 57152
rect 65648 56064 65968 57088
rect 65648 56000 65656 56064
rect 65720 56000 65736 56064
rect 65800 56000 65816 56064
rect 65880 56000 65896 56064
rect 65960 56000 65968 56064
rect 65648 54976 65968 56000
rect 65648 54912 65656 54976
rect 65720 54912 65736 54976
rect 65800 54912 65816 54976
rect 65880 54912 65896 54976
rect 65960 54912 65968 54976
rect 65648 53888 65968 54912
rect 65648 53824 65656 53888
rect 65720 53824 65736 53888
rect 65800 53824 65816 53888
rect 65880 53824 65896 53888
rect 65960 53824 65968 53888
rect 65648 52800 65968 53824
rect 65648 52736 65656 52800
rect 65720 52736 65736 52800
rect 65800 52736 65816 52800
rect 65880 52736 65896 52800
rect 65960 52736 65968 52800
rect 65648 51712 65968 52736
rect 65648 51648 65656 51712
rect 65720 51648 65736 51712
rect 65800 51648 65816 51712
rect 65880 51648 65896 51712
rect 65960 51648 65968 51712
rect 65648 50624 65968 51648
rect 65648 50560 65656 50624
rect 65720 50560 65736 50624
rect 65800 50560 65816 50624
rect 65880 50560 65896 50624
rect 65960 50560 65968 50624
rect 65648 49536 65968 50560
rect 65648 49472 65656 49536
rect 65720 49472 65736 49536
rect 65800 49472 65816 49536
rect 65880 49472 65896 49536
rect 65960 49472 65968 49536
rect 65648 48448 65968 49472
rect 65648 48384 65656 48448
rect 65720 48384 65736 48448
rect 65800 48384 65816 48448
rect 65880 48384 65896 48448
rect 65960 48384 65968 48448
rect 65648 47360 65968 48384
rect 65648 47296 65656 47360
rect 65720 47296 65736 47360
rect 65800 47296 65816 47360
rect 65880 47296 65896 47360
rect 65960 47296 65968 47360
rect 65648 46272 65968 47296
rect 65648 46208 65656 46272
rect 65720 46208 65736 46272
rect 65800 46208 65816 46272
rect 65880 46208 65896 46272
rect 65960 46208 65968 46272
rect 65648 45184 65968 46208
rect 65648 45120 65656 45184
rect 65720 45120 65736 45184
rect 65800 45120 65816 45184
rect 65880 45120 65896 45184
rect 65960 45120 65968 45184
rect 65648 44096 65968 45120
rect 65648 44032 65656 44096
rect 65720 44032 65736 44096
rect 65800 44032 65816 44096
rect 65880 44032 65896 44096
rect 65960 44032 65968 44096
rect 65648 43008 65968 44032
rect 65648 42944 65656 43008
rect 65720 42944 65736 43008
rect 65800 42944 65816 43008
rect 65880 42944 65896 43008
rect 65960 42944 65968 43008
rect 65648 41920 65968 42944
rect 65648 41856 65656 41920
rect 65720 41856 65736 41920
rect 65800 41856 65816 41920
rect 65880 41856 65896 41920
rect 65960 41856 65968 41920
rect 65648 40832 65968 41856
rect 65648 40768 65656 40832
rect 65720 40768 65736 40832
rect 65800 40768 65816 40832
rect 65880 40768 65896 40832
rect 65960 40768 65968 40832
rect 65648 39744 65968 40768
rect 65648 39680 65656 39744
rect 65720 39680 65736 39744
rect 65800 39680 65816 39744
rect 65880 39680 65896 39744
rect 65960 39680 65968 39744
rect 65648 38656 65968 39680
rect 65648 38592 65656 38656
rect 65720 38592 65736 38656
rect 65800 38592 65816 38656
rect 65880 38592 65896 38656
rect 65960 38592 65968 38656
rect 65648 37568 65968 38592
rect 65648 37504 65656 37568
rect 65720 37504 65736 37568
rect 65800 37504 65816 37568
rect 65880 37504 65896 37568
rect 65960 37504 65968 37568
rect 65648 36480 65968 37504
rect 65648 36416 65656 36480
rect 65720 36416 65736 36480
rect 65800 36416 65816 36480
rect 65880 36416 65896 36480
rect 65960 36416 65968 36480
rect 65648 35392 65968 36416
rect 65648 35328 65656 35392
rect 65720 35328 65736 35392
rect 65800 35328 65816 35392
rect 65880 35328 65896 35392
rect 65960 35328 65968 35392
rect 65648 34304 65968 35328
rect 65648 34240 65656 34304
rect 65720 34240 65736 34304
rect 65800 34240 65816 34304
rect 65880 34240 65896 34304
rect 65960 34240 65968 34304
rect 65648 33216 65968 34240
rect 65648 33152 65656 33216
rect 65720 33152 65736 33216
rect 65800 33152 65816 33216
rect 65880 33152 65896 33216
rect 65960 33152 65968 33216
rect 65648 32128 65968 33152
rect 65648 32064 65656 32128
rect 65720 32064 65736 32128
rect 65800 32064 65816 32128
rect 65880 32064 65896 32128
rect 65960 32064 65968 32128
rect 65648 31040 65968 32064
rect 65648 30976 65656 31040
rect 65720 30976 65736 31040
rect 65800 30976 65816 31040
rect 65880 30976 65896 31040
rect 65960 30976 65968 31040
rect 65648 29952 65968 30976
rect 65648 29888 65656 29952
rect 65720 29888 65736 29952
rect 65800 29888 65816 29952
rect 65880 29888 65896 29952
rect 65960 29888 65968 29952
rect 65648 28864 65968 29888
rect 65648 28800 65656 28864
rect 65720 28800 65736 28864
rect 65800 28800 65816 28864
rect 65880 28800 65896 28864
rect 65960 28800 65968 28864
rect 65648 27776 65968 28800
rect 65648 27712 65656 27776
rect 65720 27712 65736 27776
rect 65800 27712 65816 27776
rect 65880 27712 65896 27776
rect 65960 27712 65968 27776
rect 65648 26688 65968 27712
rect 65648 26624 65656 26688
rect 65720 26624 65736 26688
rect 65800 26624 65816 26688
rect 65880 26624 65896 26688
rect 65960 26624 65968 26688
rect 65648 25600 65968 26624
rect 65648 25536 65656 25600
rect 65720 25536 65736 25600
rect 65800 25536 65816 25600
rect 65880 25536 65896 25600
rect 65960 25536 65968 25600
rect 65648 24512 65968 25536
rect 65648 24448 65656 24512
rect 65720 24448 65736 24512
rect 65800 24448 65816 24512
rect 65880 24448 65896 24512
rect 65960 24448 65968 24512
rect 65648 23424 65968 24448
rect 65648 23360 65656 23424
rect 65720 23360 65736 23424
rect 65800 23360 65816 23424
rect 65880 23360 65896 23424
rect 65960 23360 65968 23424
rect 65648 22336 65968 23360
rect 65648 22272 65656 22336
rect 65720 22272 65736 22336
rect 65800 22272 65816 22336
rect 65880 22272 65896 22336
rect 65960 22272 65968 22336
rect 65648 21248 65968 22272
rect 65648 21184 65656 21248
rect 65720 21184 65736 21248
rect 65800 21184 65816 21248
rect 65880 21184 65896 21248
rect 65960 21184 65968 21248
rect 65648 20160 65968 21184
rect 65648 20096 65656 20160
rect 65720 20096 65736 20160
rect 65800 20096 65816 20160
rect 65880 20096 65896 20160
rect 65960 20096 65968 20160
rect 65648 19072 65968 20096
rect 65648 19008 65656 19072
rect 65720 19008 65736 19072
rect 65800 19008 65816 19072
rect 65880 19008 65896 19072
rect 65960 19008 65968 19072
rect 65648 17984 65968 19008
rect 65648 17920 65656 17984
rect 65720 17920 65736 17984
rect 65800 17920 65816 17984
rect 65880 17920 65896 17984
rect 65960 17920 65968 17984
rect 65648 16896 65968 17920
rect 65648 16832 65656 16896
rect 65720 16832 65736 16896
rect 65800 16832 65816 16896
rect 65880 16832 65896 16896
rect 65960 16832 65968 16896
rect 65648 15808 65968 16832
rect 65648 15744 65656 15808
rect 65720 15744 65736 15808
rect 65800 15744 65816 15808
rect 65880 15744 65896 15808
rect 65960 15744 65968 15808
rect 65648 14720 65968 15744
rect 65648 14656 65656 14720
rect 65720 14656 65736 14720
rect 65800 14656 65816 14720
rect 65880 14656 65896 14720
rect 65960 14656 65968 14720
rect 65648 13632 65968 14656
rect 65648 13568 65656 13632
rect 65720 13568 65736 13632
rect 65800 13568 65816 13632
rect 65880 13568 65896 13632
rect 65960 13568 65968 13632
rect 65648 12544 65968 13568
rect 65648 12480 65656 12544
rect 65720 12480 65736 12544
rect 65800 12480 65816 12544
rect 65880 12480 65896 12544
rect 65960 12480 65968 12544
rect 65648 11456 65968 12480
rect 65648 11392 65656 11456
rect 65720 11392 65736 11456
rect 65800 11392 65816 11456
rect 65880 11392 65896 11456
rect 65960 11392 65968 11456
rect 65648 10368 65968 11392
rect 65648 10304 65656 10368
rect 65720 10304 65736 10368
rect 65800 10304 65816 10368
rect 65880 10304 65896 10368
rect 65960 10304 65968 10368
rect 65648 9280 65968 10304
rect 65648 9216 65656 9280
rect 65720 9216 65736 9280
rect 65800 9216 65816 9280
rect 65880 9216 65896 9280
rect 65960 9216 65968 9280
rect 65648 8192 65968 9216
rect 65648 8128 65656 8192
rect 65720 8128 65736 8192
rect 65800 8128 65816 8192
rect 65880 8128 65896 8192
rect 65960 8128 65968 8192
rect 65648 7104 65968 8128
rect 65648 7040 65656 7104
rect 65720 7040 65736 7104
rect 65800 7040 65816 7104
rect 65880 7040 65896 7104
rect 65960 7040 65968 7104
rect 65648 6016 65968 7040
rect 65648 5952 65656 6016
rect 65720 5952 65736 6016
rect 65800 5952 65816 6016
rect 65880 5952 65896 6016
rect 65960 5952 65968 6016
rect 65648 4928 65968 5952
rect 65648 4864 65656 4928
rect 65720 4864 65736 4928
rect 65800 4864 65816 4928
rect 65880 4864 65896 4928
rect 65960 4864 65968 4928
rect 65648 3840 65968 4864
rect 65648 3776 65656 3840
rect 65720 3776 65736 3840
rect 65800 3776 65816 3840
rect 65880 3776 65896 3840
rect 65960 3776 65968 3840
rect 65648 2752 65968 3776
rect 65648 2688 65656 2752
rect 65720 2688 65736 2752
rect 65800 2688 65816 2752
rect 65880 2688 65896 2752
rect 65960 2688 65968 2752
rect 65648 2128 65968 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 46000 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A_N
timestamp 1649977179
transform 1 0 43332 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__S
timestamp 1649977179
transform -1 0 32292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A1
timestamp 1649977179
transform 1 0 33856 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__S
timestamp 1649977179
transform 1 0 33488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A0
timestamp 1649977179
transform -1 0 53636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__S
timestamp 1649977179
transform 1 0 45172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A
timestamp 1649977179
transform -1 0 18124 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1649977179
transform 1 0 21528 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A
timestamp 1649977179
transform 1 0 26312 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1649977179
transform 1 0 19044 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A
timestamp 1649977179
transform 1 0 23736 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A
timestamp 1649977179
transform 1 0 17664 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1649977179
transform -1 0 20056 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A
timestamp 1649977179
transform -1 0 26496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A
timestamp 1649977179
transform 1 0 23368 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1649977179
transform 1 0 18492 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1649977179
transform 1 0 33028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A
timestamp 1649977179
transform 1 0 25024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__B
timestamp 1649977179
transform -1 0 23460 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__C
timestamp 1649977179
transform -1 0 24656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A
timestamp 1649977179
transform 1 0 18768 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A
timestamp 1649977179
transform -1 0 16744 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1649977179
transform -1 0 27048 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A
timestamp 1649977179
transform 1 0 40388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A1
timestamp 1649977179
transform 1 0 23736 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A2
timestamp 1649977179
transform 1 0 22724 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__B1
timestamp 1649977179
transform -1 0 22356 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A
timestamp 1649977179
transform 1 0 30544 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__B
timestamp 1649977179
transform -1 0 31280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A0
timestamp 1649977179
transform -1 0 40020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A2
timestamp 1649977179
transform -1 0 43424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A
timestamp 1649977179
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__B_N
timestamp 1649977179
transform 1 0 22264 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A
timestamp 1649977179
transform -1 0 21988 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__B2
timestamp 1649977179
transform 1 0 21160 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A
timestamp 1649977179
transform -1 0 21620 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A
timestamp 1649977179
transform -1 0 21068 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A1
timestamp 1649977179
transform -1 0 22632 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A
timestamp 1649977179
transform 1 0 15456 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__A
timestamp 1649977179
transform 1 0 27232 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__A
timestamp 1649977179
transform -1 0 34224 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__A
timestamp 1649977179
transform -1 0 19412 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__A
timestamp 1649977179
transform 1 0 34592 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__A
timestamp 1649977179
transform 1 0 35788 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__A_N
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__B
timestamp 1649977179
transform -1 0 36984 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__A_N
timestamp 1649977179
transform -1 0 41032 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__A
timestamp 1649977179
transform 1 0 35144 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A
timestamp 1649977179
transform 1 0 37996 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__A
timestamp 1649977179
transform -1 0 39100 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A
timestamp 1649977179
transform 1 0 35604 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__A
timestamp 1649977179
transform -1 0 41676 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A
timestamp 1649977179
transform -1 0 45816 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A
timestamp 1649977179
transform -1 0 43884 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__B
timestamp 1649977179
transform 1 0 45172 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__B
timestamp 1649977179
transform -1 0 36800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1
timestamp 1649977179
transform 1 0 40664 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A1
timestamp 1649977179
transform 1 0 39192 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B_N
timestamp 1649977179
transform -1 0 31280 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__B_N
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__A_N
timestamp 1649977179
transform 1 0 37260 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A
timestamp 1649977179
transform -1 0 37444 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1284__A
timestamp 1649977179
transform 1 0 22448 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A
timestamp 1649977179
transform 1 0 38732 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__A
timestamp 1649977179
transform 1 0 38548 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A1
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__A1
timestamp 1649977179
transform -1 0 36616 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__A
timestamp 1649977179
transform 1 0 19780 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1308__A
timestamp 1649977179
transform -1 0 37444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A
timestamp 1649977179
transform 1 0 9752 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1312__A
timestamp 1649977179
transform -1 0 8464 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A
timestamp 1649977179
transform 1 0 12696 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1317__A
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__A_N
timestamp 1649977179
transform 1 0 13156 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1319__B
timestamp 1649977179
transform 1 0 14260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__A
timestamp 1649977179
transform -1 0 8280 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__A
timestamp 1649977179
transform 1 0 5428 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__A_N
timestamp 1649977179
transform 1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__B
timestamp 1649977179
transform -1 0 9016 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__A_N
timestamp 1649977179
transform 1 0 9568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__B
timestamp 1649977179
transform 1 0 7636 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__A_N
timestamp 1649977179
transform -1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__A
timestamp 1649977179
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__B
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__C_N
timestamp 1649977179
transform -1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__B1
timestamp 1649977179
transform -1 0 36892 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__B_N
timestamp 1649977179
transform -1 0 10488 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__A
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__A
timestamp 1649977179
transform 1 0 10304 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__B_N
timestamp 1649977179
transform 1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__B_N
timestamp 1649977179
transform 1 0 6992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__A_N
timestamp 1649977179
transform 1 0 6900 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__A
timestamp 1649977179
transform 1 0 10672 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__A
timestamp 1649977179
transform 1 0 12512 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__A3
timestamp 1649977179
transform 1 0 35604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__B1
timestamp 1649977179
transform 1 0 35420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__A
timestamp 1649977179
transform -1 0 24748 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__A
timestamp 1649977179
transform 1 0 24748 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__A
timestamp 1649977179
transform 1 0 23920 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__A
timestamp 1649977179
transform -1 0 34132 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__A_N
timestamp 1649977179
transform -1 0 33212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__A
timestamp 1649977179
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__A
timestamp 1649977179
transform 1 0 29808 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__A_N
timestamp 1649977179
transform 1 0 31372 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__B
timestamp 1649977179
transform 1 0 30820 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__A
timestamp 1649977179
transform 1 0 24472 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A
timestamp 1649977179
transform 1 0 23276 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__A
timestamp 1649977179
transform 1 0 28888 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__A
timestamp 1649977179
transform -1 0 26220 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__B
timestamp 1649977179
transform -1 0 29992 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__A1
timestamp 1649977179
transform -1 0 28980 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__A
timestamp 1649977179
transform 1 0 22724 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__B_N
timestamp 1649977179
transform -1 0 26588 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__B_N
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__A_N
timestamp 1649977179
transform -1 0 25208 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A
timestamp 1649977179
transform 1 0 22724 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__A1
timestamp 1649977179
transform -1 0 28888 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__A1
timestamp 1649977179
transform -1 0 27784 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__A
timestamp 1649977179
transform 1 0 30452 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__A
timestamp 1649977179
transform -1 0 17204 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__A
timestamp 1649977179
transform 1 0 15640 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__A
timestamp 1649977179
transform -1 0 13340 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__A
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__A
timestamp 1649977179
transform 1 0 7360 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__A
timestamp 1649977179
transform 1 0 10948 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__A
timestamp 1649977179
transform 1 0 18308 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__A_N
timestamp 1649977179
transform -1 0 14444 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__B
timestamp 1649977179
transform -1 0 14996 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__A_N
timestamp 1649977179
transform 1 0 37812 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__D
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__A
timestamp 1649977179
transform 1 0 17848 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__A
timestamp 1649977179
transform -1 0 15640 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__A_N
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__A
timestamp 1649977179
transform 1 0 17664 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__A
timestamp 1649977179
transform -1 0 15364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__C
timestamp 1649977179
transform -1 0 16100 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__D
timestamp 1649977179
transform 1 0 17112 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__B
timestamp 1649977179
transform 1 0 42228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__B
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1509__B
timestamp 1649977179
transform -1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__A1
timestamp 1649977179
transform 1 0 17572 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__A
timestamp 1649977179
transform 1 0 12788 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__A
timestamp 1649977179
transform 1 0 17296 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__B_N
timestamp 1649977179
transform 1 0 12052 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__B_N
timestamp 1649977179
transform -1 0 9016 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__A_N
timestamp 1649977179
transform 1 0 10488 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__A
timestamp 1649977179
transform -1 0 12328 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1520__A2
timestamp 1649977179
transform 1 0 13248 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__A1
timestamp 1649977179
transform 1 0 15180 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1522__A1
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1523__A1
timestamp 1649977179
transform 1 0 15088 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1524__A
timestamp 1649977179
transform 1 0 15456 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1525__A2
timestamp 1649977179
transform 1 0 10856 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1539__B
timestamp 1649977179
transform 1 0 9936 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1551__A2
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1555__A
timestamp 1649977179
transform -1 0 14812 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__A2
timestamp 1649977179
transform 1 0 42688 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1558__B1
timestamp 1649977179
transform -1 0 43240 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1562__A
timestamp 1649977179
transform 1 0 20148 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1564__A
timestamp 1649977179
transform 1 0 24564 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1567__A
timestamp 1649977179
transform 1 0 34868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1568__A
timestamp 1649977179
transform 1 0 26956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1569__A_N
timestamp 1649977179
transform 1 0 27784 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1570__B_N
timestamp 1649977179
transform 1 0 28704 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1573__A
timestamp 1649977179
transform 1 0 27876 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__A
timestamp 1649977179
transform 1 0 27508 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1578__A
timestamp 1649977179
transform 1 0 25576 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1580__A
timestamp 1649977179
transform -1 0 27140 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1581__A_N
timestamp 1649977179
transform 1 0 25760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__A
timestamp 1649977179
transform 1 0 24748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1589__B_N
timestamp 1649977179
transform 1 0 25208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1594__A
timestamp 1649977179
transform -1 0 28980 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1595__A
timestamp 1649977179
transform 1 0 30176 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1596__B_N
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1598__A
timestamp 1649977179
transform 1 0 29716 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1605__A
timestamp 1649977179
transform 1 0 33764 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1655__A
timestamp 1649977179
transform 1 0 42412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1656__A
timestamp 1649977179
transform -1 0 43148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1662__A
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1663__D
timestamp 1649977179
transform -1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1670__B
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1674__A
timestamp 1649977179
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1675__A1
timestamp 1649977179
transform -1 0 18768 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1677__A
timestamp 1649977179
transform 1 0 15456 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1678__A1
timestamp 1649977179
transform 1 0 19412 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1680__A
timestamp 1649977179
transform 1 0 14996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1681__A1
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1683__A
timestamp 1649977179
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1684__A1
timestamp 1649977179
transform -1 0 18952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1686__A
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1688__A1
timestamp 1649977179
transform -1 0 14904 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1690__A
timestamp 1649977179
transform 1 0 15088 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1691__A1
timestamp 1649977179
transform -1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1693__A
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1696__A
timestamp 1649977179
transform 1 0 17296 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1697__A1
timestamp 1649977179
transform -1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1699__A
timestamp 1649977179
transform 1 0 14904 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1700__A1
timestamp 1649977179
transform -1 0 17296 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1702__A
timestamp 1649977179
transform 1 0 16008 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1703__A1
timestamp 1649977179
transform 1 0 17848 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1705__A
timestamp 1649977179
transform 1 0 30636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1706__A
timestamp 1649977179
transform 1 0 22724 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1709__B
timestamp 1649977179
transform -1 0 28704 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1709__C
timestamp 1649977179
transform -1 0 27140 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1710__A
timestamp 1649977179
transform -1 0 36616 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1711__A0
timestamp 1649977179
transform 1 0 42688 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1713__A
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1714__A0
timestamp 1649977179
transform -1 0 43700 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1716__A
timestamp 1649977179
transform -1 0 28980 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1717__A0
timestamp 1649977179
transform -1 0 36892 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1719__A
timestamp 1649977179
transform -1 0 27600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1722__A
timestamp 1649977179
transform 1 0 24656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1725__A
timestamp 1649977179
transform -1 0 25852 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1726__A
timestamp 1649977179
transform 1 0 36340 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1729__A
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1730__A0
timestamp 1649977179
transform 1 0 40664 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1732__A
timestamp 1649977179
transform 1 0 20424 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1733__A0
timestamp 1649977179
transform 1 0 40848 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1735__A
timestamp 1649977179
transform -1 0 20056 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1736__A0
timestamp 1649977179
transform 1 0 40204 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1738__A
timestamp 1649977179
transform 1 0 19412 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1739__A0
timestamp 1649977179
transform 1 0 35880 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1741__A
timestamp 1649977179
transform 1 0 18584 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1742__A0
timestamp 1649977179
transform 1 0 34040 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1742__S
timestamp 1649977179
transform 1 0 34684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1746__B
timestamp 1649977179
transform -1 0 23460 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1746__C_N
timestamp 1649977179
transform 1 0 22632 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1748__A0
timestamp 1649977179
transform 1 0 42228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1750__A0
timestamp 1649977179
transform 1 0 43148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1752__A0
timestamp 1649977179
transform 1 0 37536 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1761__A0
timestamp 1649977179
transform 1 0 37812 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1763__A0
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1765__A0
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1767__A0
timestamp 1649977179
transform 1 0 36524 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1769__A0
timestamp 1649977179
transform 1 0 34592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1772__B
timestamp 1649977179
transform 1 0 14168 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1776__A1
timestamp 1649977179
transform 1 0 7728 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1778__A1
timestamp 1649977179
transform 1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1780__A1
timestamp 1649977179
transform -1 0 4600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1782__A1
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1785__A1
timestamp 1649977179
transform 1 0 6164 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1787__A1
timestamp 1649977179
transform 1 0 12604 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1791__A1
timestamp 1649977179
transform 1 0 8464 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1793__A1
timestamp 1649977179
transform 1 0 11868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1795__A1
timestamp 1649977179
transform 1 0 13156 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1798__A
timestamp 1649977179
transform -1 0 13708 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1802__A1
timestamp 1649977179
transform 1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1804__A1
timestamp 1649977179
transform 1 0 7544 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1806__A1
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1808__A1
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1811__A1
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1813__A1
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1817__A1
timestamp 1649977179
transform 1 0 7176 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1819__A1
timestamp 1649977179
transform 1 0 5612 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1821__A1
timestamp 1649977179
transform -1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1823__B
timestamp 1649977179
transform -1 0 24564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1823__C
timestamp 1649977179
transform 1 0 23828 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1825__A0
timestamp 1649977179
transform 1 0 33580 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1827__A0
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1829__A0
timestamp 1649977179
transform 1 0 31464 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1838__A0
timestamp 1649977179
transform 1 0 27324 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1840__A0
timestamp 1649977179
transform -1 0 23920 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1842__A0
timestamp 1649977179
transform 1 0 27048 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1844__A0
timestamp 1649977179
transform 1 0 25116 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1846__A0
timestamp 1649977179
transform -1 0 31372 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1848__A
timestamp 1649977179
transform 1 0 24748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1848__B
timestamp 1649977179
transform -1 0 27784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1848__C_N
timestamp 1649977179
transform 1 0 25024 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1849__A
timestamp 1649977179
transform 1 0 26864 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1850__A0
timestamp 1649977179
transform -1 0 30452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1852__A0
timestamp 1649977179
transform -1 0 29440 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1854__A0
timestamp 1649977179
transform -1 0 28428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1860__A
timestamp 1649977179
transform 1 0 25852 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1863__A0
timestamp 1649977179
transform 1 0 21620 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1865__A0
timestamp 1649977179
transform 1 0 23276 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1867__A0
timestamp 1649977179
transform -1 0 22632 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1869__A0
timestamp 1649977179
transform 1 0 23000 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1871__A0
timestamp 1649977179
transform 1 0 27048 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1871__S
timestamp 1649977179
transform 1 0 25668 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1874__B
timestamp 1649977179
transform -1 0 12880 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1875__A
timestamp 1649977179
transform -1 0 12880 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1878__A1
timestamp 1649977179
transform -1 0 10120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1880__A1
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1882__A1
timestamp 1649977179
transform 1 0 13432 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1884__A1
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1886__A
timestamp 1649977179
transform -1 0 8464 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1887__A1
timestamp 1649977179
transform 1 0 7544 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1889__A1
timestamp 1649977179
transform -1 0 4692 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1893__A1
timestamp 1649977179
transform -1 0 9108 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1895__A1
timestamp 1649977179
transform -1 0 8464 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1897__A1
timestamp 1649977179
transform -1 0 11868 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1897__S
timestamp 1649977179
transform -1 0 11316 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1899__B
timestamp 1649977179
transform 1 0 16928 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1901__A1
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1903__A1
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1905__A1
timestamp 1649977179
transform -1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1907__A1
timestamp 1649977179
transform -1 0 13432 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1909__A1
timestamp 1649977179
transform -1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1912__A1
timestamp 1649977179
transform 1 0 11040 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1914__A1
timestamp 1649977179
transform -1 0 14996 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1916__A1
timestamp 1649977179
transform -1 0 13156 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1918__A1
timestamp 1649977179
transform -1 0 14996 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1920__A1
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1922__A1
timestamp 1649977179
transform 1 0 14904 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1924__B
timestamp 1649977179
transform 1 0 22908 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1924__C
timestamp 1649977179
transform -1 0 22356 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1925__A
timestamp 1649977179
transform 1 0 33396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1926__A0
timestamp 1649977179
transform 1 0 31188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1928__A0
timestamp 1649977179
transform 1 0 32568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1930__A0
timestamp 1649977179
transform 1 0 33304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1936__A
timestamp 1649977179
transform 1 0 30636 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1939__A0
timestamp 1649977179
transform 1 0 31464 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1941__A0
timestamp 1649977179
transform 1 0 30268 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1943__A0
timestamp 1649977179
transform 1 0 33304 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1945__A0
timestamp 1649977179
transform 1 0 28888 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1947__A0
timestamp 1649977179
transform 1 0 34592 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1947__S
timestamp 1649977179
transform 1 0 34776 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1949__A
timestamp 1649977179
transform 1 0 20792 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1949__C_N
timestamp 1649977179
transform 1 0 22080 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1953__A0
timestamp 1649977179
transform 1 0 21896 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1955__A0
timestamp 1649977179
transform 1 0 21988 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1957__A0
timestamp 1649977179
transform 1 0 21804 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1959__A0
timestamp 1649977179
transform -1 0 25760 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1962__A0
timestamp 1649977179
transform 1 0 15456 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1964__A0
timestamp 1649977179
transform -1 0 16836 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1968__A0
timestamp 1649977179
transform -1 0 21252 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1970__A0
timestamp 1649977179
transform -1 0 18032 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1972__A0
timestamp 1649977179
transform 1 0 21160 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1978__A0
timestamp 1649977179
transform 1 0 30360 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1978__A1
timestamp 1649977179
transform 1 0 28704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1980__A0
timestamp 1649977179
transform -1 0 27968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1980__A1
timestamp 1649977179
transform 1 0 28336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1982__A1
timestamp 1649977179
transform 1 0 26312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1984__A1
timestamp 1649977179
transform 1 0 26312 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1986__A1
timestamp 1649977179
transform 1 0 23368 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1989__A1
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1991__A1
timestamp 1649977179
transform 1 0 18216 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1993__A1
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1995__A1
timestamp 1649977179
transform 1 0 18584 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1997__A1
timestamp 1649977179
transform 1 0 16744 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1999__A1
timestamp 1649977179
transform 1 0 18216 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2001__A0
timestamp 1649977179
transform -1 0 18676 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2004__A
timestamp 1649977179
transform -1 0 43332 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2005__A
timestamp 1649977179
transform -1 0 43424 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2011__A
timestamp 1649977179
transform 1 0 41952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2017__A
timestamp 1649977179
transform -1 0 38180 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2023__A
timestamp 1649977179
transform -1 0 24380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2029__A
timestamp 1649977179
transform 1 0 25024 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2035__A
timestamp 1649977179
transform 1 0 41308 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2036__A
timestamp 1649977179
transform -1 0 21344 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2037__A
timestamp 1649977179
transform -1 0 44068 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2038__A
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2039__A
timestamp 1649977179
transform 1 0 30728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2040__A
timestamp 1649977179
transform 1 0 39836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2041__A
timestamp 1649977179
transform -1 0 40664 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2208__D
timestamp 1649977179
transform 1 0 36156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2470__A
timestamp 1649977179
transform 1 0 53360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2471__A
timestamp 1649977179
transform -1 0 56120 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2472__A
timestamp 1649977179
transform -1 0 61364 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2473__A
timestamp 1649977179
transform -1 0 67988 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2474__A
timestamp 1649977179
transform -1 0 58512 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2475__A
timestamp 1649977179
transform -1 0 67988 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2476__A
timestamp 1649977179
transform 1 0 66608 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2477__A
timestamp 1649977179
transform -1 0 67988 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2478__A
timestamp 1649977179
transform -1 0 67988 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 26036 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 13248 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 18216 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 18676 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 13984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 13432 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 20424 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 20240 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 33856 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 33488 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 38180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 40020 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 32660 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 37536 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_wb_clk_i_A
timestamp 1649977179
transform 1 0 37352 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 56028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 51152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 51796 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 50968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 49680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 46920 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 50324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 47932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 8464 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 19412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 21988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 21988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 7452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 10488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 7268 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 17296 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 8004 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 9844 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 9200 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 10396 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 24564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 9108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 9752 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 6716 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 8188 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output41_A
timestamp 1649977179
transform 1 0 54004 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output44_A
timestamp 1649977179
transform 1 0 54648 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output45_A
timestamp 1649977179
transform 1 0 55752 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output46_A
timestamp 1649977179
transform 1 0 55200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output47_A
timestamp 1649977179
transform 1 0 56304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output48_A
timestamp 1649977179
transform 1 0 54556 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output49_A
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output52_A
timestamp 1649977179
transform 1 0 39192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1649977179
transform -1 0 67436 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101
timestamp 1649977179
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1649977179
transform 1 0 12144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_130
timestamp 1649977179
transform 1 0 13064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1649977179
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_181 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_227
timestamp 1649977179
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1649977179
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1649977179
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_255
timestamp 1649977179
transform 1 0 24564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_269
timestamp 1649977179
transform 1 0 25852 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_281 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_290
timestamp 1649977179
transform 1 0 27784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_318
timestamp 1649977179
transform 1 0 30360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_325
timestamp 1649977179
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_339
timestamp 1649977179
transform 1 0 32292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_346
timestamp 1649977179
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_353
timestamp 1649977179
transform 1 0 33580 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_369
timestamp 1649977179
transform 1 0 35052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_376
timestamp 1649977179
transform 1 0 35696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1649977179
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1649977179
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1649977179
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_421
timestamp 1649977179
transform 1 0 39836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_426
timestamp 1649977179
transform 1 0 40296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_434
timestamp 1649977179
transform 1 0 41032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_442
timestamp 1649977179
transform 1 0 41768 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_453
timestamp 1649977179
transform 1 0 42780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1649977179
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_469
timestamp 1649977179
transform 1 0 44252 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1649977179
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_481
timestamp 1649977179
transform 1 0 45356 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_489
timestamp 1649977179
transform 1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_497
timestamp 1649977179
transform 1 0 46828 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_503
timestamp 1649977179
transform 1 0 47380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_505
timestamp 1649977179
transform 1 0 47564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_513
timestamp 1649977179
transform 1 0 48300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_520
timestamp 1649977179
transform 1 0 48944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_527
timestamp 1649977179
transform 1 0 49588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_531
timestamp 1649977179
transform 1 0 49956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_546
timestamp 1649977179
transform 1 0 51336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_554
timestamp 1649977179
transform 1 0 52072 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_565
timestamp 1649977179
transform 1 0 53084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_573
timestamp 1649977179
transform 1 0 53820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_581
timestamp 1649977179
transform 1 0 54556 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_587
timestamp 1649977179
transform 1 0 55108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_593
timestamp 1649977179
transform 1 0 55660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_601
timestamp 1649977179
transform 1 0 56396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_608
timestamp 1649977179
transform 1 0 57040 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_627
timestamp 1649977179
transform 1 0 58788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_634
timestamp 1649977179
transform 1 0 59432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_642
timestamp 1649977179
transform 1 0 60168 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_645
timestamp 1649977179
transform 1 0 60444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_657
timestamp 1649977179
transform 1 0 61548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_669
timestamp 1649977179
transform 1 0 62652 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_673
timestamp 1649977179
transform 1 0 63020 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_685
timestamp 1649977179
transform 1 0 64124 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_697
timestamp 1649977179
transform 1 0 65228 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_701
timestamp 1649977179
transform 1 0 65596 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_713
timestamp 1649977179
transform 1 0 66700 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_725
timestamp 1649977179
transform 1 0 67804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_729
timestamp 1649977179
transform 1 0 68172 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_65
timestamp 1649977179
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_75
timestamp 1649977179
transform 1 0 8004 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_87
timestamp 1649977179
transform 1 0 9108 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_94
timestamp 1649977179
transform 1 0 9752 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_101
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_120
timestamp 1649977179
transform 1 0 12144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_128
timestamp 1649977179
transform 1 0 12880 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_146
timestamp 1649977179
transform 1 0 14536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_150
timestamp 1649977179
transform 1 0 14904 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1649977179
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_177
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_185
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_227
timestamp 1649977179
transform 1 0 21988 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1649977179
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_241
timestamp 1649977179
transform 1 0 23276 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_255
timestamp 1649977179
transform 1 0 24564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_269
timestamp 1649977179
transform 1 0 25852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1649977179
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_286
timestamp 1649977179
transform 1 0 27416 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_300
timestamp 1649977179
transform 1 0 28704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_324
timestamp 1649977179
transform 1 0 30912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_328
timestamp 1649977179
transform 1 0 31280 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_346
timestamp 1649977179
transform 1 0 32936 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_352
timestamp 1649977179
transform 1 0 33488 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_356
timestamp 1649977179
transform 1 0 33856 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_363
timestamp 1649977179
transform 1 0 34500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_370
timestamp 1649977179
transform 1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_377
timestamp 1649977179
transform 1 0 35788 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_386
timestamp 1649977179
transform 1 0 36616 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_396
timestamp 1649977179
transform 1 0 37536 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1649977179
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1649977179
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_453
timestamp 1649977179
transform 1 0 42780 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_481
timestamp 1649977179
transform 1 0 45356 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_489
timestamp 1649977179
transform 1 0 46092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_496
timestamp 1649977179
transform 1 0 46736 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_515
timestamp 1649977179
transform 1 0 48484 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_521
timestamp 1649977179
transform 1 0 49036 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_529
timestamp 1649977179
transform 1 0 49772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_538
timestamp 1649977179
transform 1 0 50600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_544
timestamp 1649977179
transform 1 0 51152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_552
timestamp 1649977179
transform 1 0 51888 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_565
timestamp 1649977179
transform 1 0 53084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_573
timestamp 1649977179
transform 1 0 53820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_581
timestamp 1649977179
transform 1 0 54556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_589
timestamp 1649977179
transform 1 0 55292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_596
timestamp 1649977179
transform 1 0 55936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_603
timestamp 1649977179
transform 1 0 56580 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_610
timestamp 1649977179
transform 1 0 57224 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_627
timestamp 1649977179
transform 1 0 58788 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_639
timestamp 1649977179
transform 1 0 59892 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_651
timestamp 1649977179
transform 1 0 60996 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_663
timestamp 1649977179
transform 1 0 62100 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_671
timestamp 1649977179
transform 1 0 62836 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_673
timestamp 1649977179
transform 1 0 63020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_685
timestamp 1649977179
transform 1 0 64124 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_697
timestamp 1649977179
transform 1 0 65228 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_709
timestamp 1649977179
transform 1 0 66332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_721
timestamp 1649977179
transform 1 0 67436 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_727
timestamp 1649977179
transform 1 0 67988 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_729
timestamp 1649977179
transform 1 0 68172 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_71
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1649977179
transform 1 0 9200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_94
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_108
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_115
timestamp 1649977179
transform 1 0 11684 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1649977179
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1649977179
transform 1 0 14720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_163
timestamp 1649977179
transform 1 0 16100 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_174
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_203
timestamp 1649977179
transform 1 0 19780 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_215
timestamp 1649977179
transform 1 0 20884 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_223
timestamp 1649977179
transform 1 0 21620 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_227
timestamp 1649977179
transform 1 0 21988 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1649977179
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1649977179
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1649977179
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_269
timestamp 1649977179
transform 1 0 25852 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_276
timestamp 1649977179
transform 1 0 26496 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_283
timestamp 1649977179
transform 1 0 27140 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_290
timestamp 1649977179
transform 1 0 27784 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_297
timestamp 1649977179
transform 1 0 28428 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1649977179
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_318
timestamp 1649977179
transform 1 0 30360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_342
timestamp 1649977179
transform 1 0 32568 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_353
timestamp 1649977179
transform 1 0 33580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1649977179
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_371
timestamp 1649977179
transform 1 0 35236 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_375
timestamp 1649977179
transform 1 0 35604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_399
timestamp 1649977179
transform 1 0 37812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_406
timestamp 1649977179
transform 1 0 38456 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_410
timestamp 1649977179
transform 1 0 38824 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_414
timestamp 1649977179
transform 1 0 39192 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_441
timestamp 1649977179
transform 1 0 41676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_454
timestamp 1649977179
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_462
timestamp 1649977179
transform 1 0 43608 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_470
timestamp 1649977179
transform 1 0 44344 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_486
timestamp 1649977179
transform 1 0 45816 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_493
timestamp 1649977179
transform 1 0 46460 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_504
timestamp 1649977179
transform 1 0 47472 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_511
timestamp 1649977179
transform 1 0 48116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_515
timestamp 1649977179
transform 1 0 48484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1649977179
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_535
timestamp 1649977179
transform 1 0 50324 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_551
timestamp 1649977179
transform 1 0 51796 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_558
timestamp 1649977179
transform 1 0 52440 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_565
timestamp 1649977179
transform 1 0 53084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_571
timestamp 1649977179
transform 1 0 53636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_579
timestamp 1649977179
transform 1 0 54372 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1649977179
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_592
timestamp 1649977179
transform 1 0 55568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_599
timestamp 1649977179
transform 1 0 56212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_606
timestamp 1649977179
transform 1 0 56856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_613
timestamp 1649977179
transform 1 0 57500 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_620
timestamp 1649977179
transform 1 0 58144 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_627
timestamp 1649977179
transform 1 0 58788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_639
timestamp 1649977179
transform 1 0 59892 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_643
timestamp 1649977179
transform 1 0 60260 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_645
timestamp 1649977179
transform 1 0 60444 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_657
timestamp 1649977179
transform 1 0 61548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_669
timestamp 1649977179
transform 1 0 62652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_681
timestamp 1649977179
transform 1 0 63756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_693
timestamp 1649977179
transform 1 0 64860 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_699
timestamp 1649977179
transform 1 0 65412 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_701
timestamp 1649977179
transform 1 0 65596 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_713
timestamp 1649977179
transform 1 0 66700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_717
timestamp 1649977179
transform 1 0 67068 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_721
timestamp 1649977179
transform 1 0 67436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_727
timestamp 1649977179
transform 1 0 67988 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_77
timestamp 1649977179
transform 1 0 8188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_83
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_89
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_95
timestamp 1649977179
transform 1 0 9844 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_101
timestamp 1649977179
transform 1 0 10396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_120
timestamp 1649977179
transform 1 0 12144 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1649977179
transform 1 0 12788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_134
timestamp 1649977179
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_142
timestamp 1649977179
transform 1 0 14168 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_150
timestamp 1649977179
transform 1 0 14904 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_177
timestamp 1649977179
transform 1 0 17388 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_186
timestamp 1649977179
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_192
timestamp 1649977179
transform 1 0 18768 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_213
timestamp 1649977179
transform 1 0 20700 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_228
timestamp 1649977179
transform 1 0 22080 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_236
timestamp 1649977179
transform 1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_242
timestamp 1649977179
transform 1 0 23368 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_255
timestamp 1649977179
transform 1 0 24564 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_272
timestamp 1649977179
transform 1 0 26128 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_289
timestamp 1649977179
transform 1 0 27692 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_304
timestamp 1649977179
transform 1 0 29072 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_311
timestamp 1649977179
transform 1 0 29716 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_318
timestamp 1649977179
transform 1 0 30360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_324
timestamp 1649977179
transform 1 0 30912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_331
timestamp 1649977179
transform 1 0 31556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_339
timestamp 1649977179
transform 1 0 32292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_352
timestamp 1649977179
transform 1 0 33488 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_358
timestamp 1649977179
transform 1 0 34040 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_370
timestamp 1649977179
transform 1 0 35144 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_382
timestamp 1649977179
transform 1 0 36248 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1649977179
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_396
timestamp 1649977179
transform 1 0 37536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1649977179
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_410
timestamp 1649977179
transform 1 0 38824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_417
timestamp 1649977179
transform 1 0 39468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_423
timestamp 1649977179
transform 1 0 40020 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_430
timestamp 1649977179
transform 1 0 40664 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_434
timestamp 1649977179
transform 1 0 41032 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_444
timestamp 1649977179
transform 1 0 41952 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_453
timestamp 1649977179
transform 1 0 42780 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_459
timestamp 1649977179
transform 1 0 43332 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_480
timestamp 1649977179
transform 1 0 45264 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_3_495
timestamp 1649977179
transform 1 0 46644 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_508
timestamp 1649977179
transform 1 0 47840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_515
timestamp 1649977179
transform 1 0 48484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_521
timestamp 1649977179
transform 1 0 49036 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_529
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_539
timestamp 1649977179
transform 1 0 50692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_546
timestamp 1649977179
transform 1 0 51336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_564
timestamp 1649977179
transform 1 0 52992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_571
timestamp 1649977179
transform 1 0 53636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_578
timestamp 1649977179
transform 1 0 54280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_584
timestamp 1649977179
transform 1 0 54832 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_590
timestamp 1649977179
transform 1 0 55384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_596
timestamp 1649977179
transform 1 0 55936 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_602
timestamp 1649977179
transform 1 0 56488 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_614
timestamp 1649977179
transform 1 0 57592 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_617
timestamp 1649977179
transform 1 0 57868 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_629
timestamp 1649977179
transform 1 0 58972 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_641
timestamp 1649977179
transform 1 0 60076 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_653
timestamp 1649977179
transform 1 0 61180 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_665
timestamp 1649977179
transform 1 0 62284 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_671
timestamp 1649977179
transform 1 0 62836 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_673
timestamp 1649977179
transform 1 0 63020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_685
timestamp 1649977179
transform 1 0 64124 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_697
timestamp 1649977179
transform 1 0 65228 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_709
timestamp 1649977179
transform 1 0 66332 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_717
timestamp 1649977179
transform 1 0 67068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_724
timestamp 1649977179
transform 1 0 67712 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_729
timestamp 1649977179
transform 1 0 68172 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1649977179
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_96
timestamp 1649977179
transform 1 0 9936 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_102
timestamp 1649977179
transform 1 0 10488 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_108
timestamp 1649977179
transform 1 0 11040 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_115
timestamp 1649977179
transform 1 0 11684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_122
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_129
timestamp 1649977179
transform 1 0 12972 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_146
timestamp 1649977179
transform 1 0 14536 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_155
timestamp 1649977179
transform 1 0 15364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_174
timestamp 1649977179
transform 1 0 17112 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_185
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1649977179
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_213
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_220
timestamp 1649977179
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_226
timestamp 1649977179
transform 1 0 21896 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1649977179
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_258
timestamp 1649977179
transform 1 0 24840 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_270
timestamp 1649977179
transform 1 0 25944 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_282
timestamp 1649977179
transform 1 0 27048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_286
timestamp 1649977179
transform 1 0 27416 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_290
timestamp 1649977179
transform 1 0 27784 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_302
timestamp 1649977179
transform 1 0 28888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_313
timestamp 1649977179
transform 1 0 29900 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_317
timestamp 1649977179
transform 1 0 30268 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_325
timestamp 1649977179
transform 1 0 31004 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_329
timestamp 1649977179
transform 1 0 31372 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_338
timestamp 1649977179
transform 1 0 32200 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_350
timestamp 1649977179
transform 1 0 33304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_354
timestamp 1649977179
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_362
timestamp 1649977179
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_397
timestamp 1649977179
transform 1 0 37628 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_406
timestamp 1649977179
transform 1 0 38456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_423
timestamp 1649977179
transform 1 0 40020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_436
timestamp 1649977179
transform 1 0 41216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_449
timestamp 1649977179
transform 1 0 42412 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_456
timestamp 1649977179
transform 1 0 43056 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_463
timestamp 1649977179
transform 1 0 43700 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_470
timestamp 1649977179
transform 1 0 44344 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_480
timestamp 1649977179
transform 1 0 45264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_487
timestamp 1649977179
transform 1 0 45908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_494
timestamp 1649977179
transform 1 0 46552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_501
timestamp 1649977179
transform 1 0 47196 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_508
timestamp 1649977179
transform 1 0 47840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_515
timestamp 1649977179
transform 1 0 48484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_522
timestamp 1649977179
transform 1 0 49128 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_528
timestamp 1649977179
transform 1 0 49680 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_536
timestamp 1649977179
transform 1 0 50416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_543
timestamp 1649977179
transform 1 0 51060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_550
timestamp 1649977179
transform 1 0 51704 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_557
timestamp 1649977179
transform 1 0 52348 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_564
timestamp 1649977179
transform 1 0 52992 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_571
timestamp 1649977179
transform 1 0 53636 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_577
timestamp 1649977179
transform 1 0 54188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_583
timestamp 1649977179
transform 1 0 54740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1649977179
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_591
timestamp 1649977179
transform 1 0 55476 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_597
timestamp 1649977179
transform 1 0 56028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_609
timestamp 1649977179
transform 1 0 57132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_621
timestamp 1649977179
transform 1 0 58236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_633
timestamp 1649977179
transform 1 0 59340 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_641
timestamp 1649977179
transform 1 0 60076 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_645
timestamp 1649977179
transform 1 0 60444 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_657
timestamp 1649977179
transform 1 0 61548 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_669
timestamp 1649977179
transform 1 0 62652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_681
timestamp 1649977179
transform 1 0 63756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_693
timestamp 1649977179
transform 1 0 64860 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_699
timestamp 1649977179
transform 1 0 65412 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_701
timestamp 1649977179
transform 1 0 65596 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_713
timestamp 1649977179
transform 1 0 66700 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_725
timestamp 1649977179
transform 1 0 67804 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_60
timestamp 1649977179
transform 1 0 6624 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_72
timestamp 1649977179
transform 1 0 7728 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_84
timestamp 1649977179
transform 1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1649977179
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_119
timestamp 1649977179
transform 1 0 12052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_126
timestamp 1649977179
transform 1 0 12696 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_133
timestamp 1649977179
transform 1 0 13340 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_140
timestamp 1649977179
transform 1 0 13984 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_147
timestamp 1649977179
transform 1 0 14628 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_154
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_162
timestamp 1649977179
transform 1 0 16008 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_173
timestamp 1649977179
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_177
timestamp 1649977179
transform 1 0 17388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_184
timestamp 1649977179
transform 1 0 18032 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1649977179
transform 1 0 18676 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_211
timestamp 1649977179
transform 1 0 20516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_228
timestamp 1649977179
transform 1 0 22080 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_235
timestamp 1649977179
transform 1 0 22724 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_248
timestamp 1649977179
transform 1 0 23920 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_304
timestamp 1649977179
transform 1 0 29072 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_316
timestamp 1649977179
transform 1 0 30176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_322
timestamp 1649977179
transform 1 0 30728 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_328
timestamp 1649977179
transform 1 0 31280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_346
timestamp 1649977179
transform 1 0 32936 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_358
timestamp 1649977179
transform 1 0 34040 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_370
timestamp 1649977179
transform 1 0 35144 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_378
timestamp 1649977179
transform 1 0 35880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_382
timestamp 1649977179
transform 1 0 36248 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1649977179
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_402
timestamp 1649977179
transform 1 0 38088 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_409
timestamp 1649977179
transform 1 0 38732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_417
timestamp 1649977179
transform 1 0 39468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_427
timestamp 1649977179
transform 1 0 40388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_440
timestamp 1649977179
transform 1 0 41584 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_455
timestamp 1649977179
transform 1 0 42964 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_461
timestamp 1649977179
transform 1 0 43516 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_467
timestamp 1649977179
transform 1 0 44068 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_481
timestamp 1649977179
transform 1 0 45356 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_488
timestamp 1649977179
transform 1 0 46000 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_495
timestamp 1649977179
transform 1 0 46644 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1649977179
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_508
timestamp 1649977179
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_515
timestamp 1649977179
transform 1 0 48484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_533
timestamp 1649977179
transform 1 0 50140 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_540
timestamp 1649977179
transform 1 0 50784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_547
timestamp 1649977179
transform 1 0 51428 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_554
timestamp 1649977179
transform 1 0 52072 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_564
timestamp 1649977179
transform 1 0 52992 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_570
timestamp 1649977179
transform 1 0 53544 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_582
timestamp 1649977179
transform 1 0 54648 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_594
timestamp 1649977179
transform 1 0 55752 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_606
timestamp 1649977179
transform 1 0 56856 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_614
timestamp 1649977179
transform 1 0 57592 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_629
timestamp 1649977179
transform 1 0 58972 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_641
timestamp 1649977179
transform 1 0 60076 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_653
timestamp 1649977179
transform 1 0 61180 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_665
timestamp 1649977179
transform 1 0 62284 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_671
timestamp 1649977179
transform 1 0 62836 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_673
timestamp 1649977179
transform 1 0 63020 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_685
timestamp 1649977179
transform 1 0 64124 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_697
timestamp 1649977179
transform 1 0 65228 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_709
timestamp 1649977179
transform 1 0 66332 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_721
timestamp 1649977179
transform 1 0 67436 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_727
timestamp 1649977179
transform 1 0 67988 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_729
timestamp 1649977179
transform 1 0 68172 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_49
timestamp 1649977179
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_67
timestamp 1649977179
transform 1 0 7268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_71
timestamp 1649977179
transform 1 0 7636 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_74
timestamp 1649977179
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_92
timestamp 1649977179
transform 1 0 9568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_96
timestamp 1649977179
transform 1 0 9936 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_113
timestamp 1649977179
transform 1 0 11500 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_120
timestamp 1649977179
transform 1 0 12144 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_129
timestamp 1649977179
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_144
timestamp 1649977179
transform 1 0 14352 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_152
timestamp 1649977179
transform 1 0 15088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_166
timestamp 1649977179
transform 1 0 16376 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_174
timestamp 1649977179
transform 1 0 17112 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_178
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_185
timestamp 1649977179
transform 1 0 18124 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_192
timestamp 1649977179
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_207
timestamp 1649977179
transform 1 0 20148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_219
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_229
timestamp 1649977179
transform 1 0 22172 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_242
timestamp 1649977179
transform 1 0 23368 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1649977179
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_256
timestamp 1649977179
transform 1 0 24656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_262
timestamp 1649977179
transform 1 0 25208 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_271
timestamp 1649977179
transform 1 0 26036 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_291
timestamp 1649977179
transform 1 0 27876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_299
timestamp 1649977179
transform 1 0 28612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_302
timestamp 1649977179
transform 1 0 28888 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_318
timestamp 1649977179
transform 1 0 30360 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_324
timestamp 1649977179
transform 1 0 30912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_353
timestamp 1649977179
transform 1 0 33580 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_358
timestamp 1649977179
transform 1 0 34040 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_373
timestamp 1649977179
transform 1 0 35420 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_394
timestamp 1649977179
transform 1 0 37352 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_407
timestamp 1649977179
transform 1 0 38548 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_416
timestamp 1649977179
transform 1 0 39376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_421
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_428
timestamp 1649977179
transform 1 0 40480 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_442
timestamp 1649977179
transform 1 0 41768 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_454
timestamp 1649977179
transform 1 0 42872 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_466
timestamp 1649977179
transform 1 0 43976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1649977179
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_485
timestamp 1649977179
transform 1 0 45724 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_490
timestamp 1649977179
transform 1 0 46184 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_497
timestamp 1649977179
transform 1 0 46828 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_517
timestamp 1649977179
transform 1 0 48668 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_526
timestamp 1649977179
transform 1 0 49496 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_551
timestamp 1649977179
transform 1 0 51796 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_563
timestamp 1649977179
transform 1 0 52900 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_575
timestamp 1649977179
transform 1 0 54004 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1649977179
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_589
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_601
timestamp 1649977179
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_613
timestamp 1649977179
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_625
timestamp 1649977179
transform 1 0 58604 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_637
timestamp 1649977179
transform 1 0 59708 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_643
timestamp 1649977179
transform 1 0 60260 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_645
timestamp 1649977179
transform 1 0 60444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_657
timestamp 1649977179
transform 1 0 61548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_669
timestamp 1649977179
transform 1 0 62652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_681
timestamp 1649977179
transform 1 0 63756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_693
timestamp 1649977179
transform 1 0 64860 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_699
timestamp 1649977179
transform 1 0 65412 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_701
timestamp 1649977179
transform 1 0 65596 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_713
timestamp 1649977179
transform 1 0 66700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_725
timestamp 1649977179
transform 1 0 67804 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_72
timestamp 1649977179
transform 1 0 7728 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_78
timestamp 1649977179
transform 1 0 8280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_95
timestamp 1649977179
transform 1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_129
timestamp 1649977179
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1649977179
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_172
timestamp 1649977179
transform 1 0 16928 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_185
timestamp 1649977179
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1649977179
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_198
timestamp 1649977179
transform 1 0 19320 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_210
timestamp 1649977179
transform 1 0 20424 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_214
timestamp 1649977179
transform 1 0 20792 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_231
timestamp 1649977179
transform 1 0 22356 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_243
timestamp 1649977179
transform 1 0 23460 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_267
timestamp 1649977179
transform 1 0 25668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1649977179
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_301
timestamp 1649977179
transform 1 0 28796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_311
timestamp 1649977179
transform 1 0 29716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_315
timestamp 1649977179
transform 1 0 30084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1649977179
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_345
timestamp 1649977179
transform 1 0 32844 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_367
timestamp 1649977179
transform 1 0 34868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_379
timestamp 1649977179
transform 1 0 35972 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_396
timestamp 1649977179
transform 1 0 37536 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_408
timestamp 1649977179
transform 1 0 38640 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_420
timestamp 1649977179
transform 1 0 39744 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_444
timestamp 1649977179
transform 1 0 41952 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_486
timestamp 1649977179
transform 1 0 45816 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_494
timestamp 1649977179
transform 1 0 46552 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_498
timestamp 1649977179
transform 1 0 46920 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_534
timestamp 1649977179
transform 1 0 50232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_541
timestamp 1649977179
transform 1 0 50876 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_548
timestamp 1649977179
transform 1 0 51520 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_561
timestamp 1649977179
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_573
timestamp 1649977179
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_585
timestamp 1649977179
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_597
timestamp 1649977179
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_609
timestamp 1649977179
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_629
timestamp 1649977179
transform 1 0 58972 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_641
timestamp 1649977179
transform 1 0 60076 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_653
timestamp 1649977179
transform 1 0 61180 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_665
timestamp 1649977179
transform 1 0 62284 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_671
timestamp 1649977179
transform 1 0 62836 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_673
timestamp 1649977179
transform 1 0 63020 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_685
timestamp 1649977179
transform 1 0 64124 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_697
timestamp 1649977179
transform 1 0 65228 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_709
timestamp 1649977179
transform 1 0 66332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_721
timestamp 1649977179
transform 1 0 67436 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_727
timestamp 1649977179
transform 1 0 67988 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_729
timestamp 1649977179
transform 1 0 68172 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_45
timestamp 1649977179
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_62
timestamp 1649977179
transform 1 0 6808 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_75
timestamp 1649977179
transform 1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1649977179
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_98
timestamp 1649977179
transform 1 0 10120 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_105
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_111
timestamp 1649977179
transform 1 0 11316 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1649977179
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_143
timestamp 1649977179
transform 1 0 14260 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_163
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_170
timestamp 1649977179
transform 1 0 16744 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_176
timestamp 1649977179
transform 1 0 17296 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_188
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1649977179
transform 1 0 18768 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_201
timestamp 1649977179
transform 1 0 19596 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_207
timestamp 1649977179
transform 1 0 20148 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_213
timestamp 1649977179
transform 1 0 20700 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_223
timestamp 1649977179
transform 1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_230
timestamp 1649977179
transform 1 0 22264 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_236
timestamp 1649977179
transform 1 0 22816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_240
timestamp 1649977179
transform 1 0 23184 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1649977179
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_258
timestamp 1649977179
transform 1 0 24840 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_280
timestamp 1649977179
transform 1 0 26864 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_286
timestamp 1649977179
transform 1 0 27416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_292
timestamp 1649977179
transform 1 0 27968 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_298
timestamp 1649977179
transform 1 0 28520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_306
timestamp 1649977179
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_314
timestamp 1649977179
transform 1 0 29992 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_320
timestamp 1649977179
transform 1 0 30544 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_332
timestamp 1649977179
transform 1 0 31648 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_344
timestamp 1649977179
transform 1 0 32752 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_349
timestamp 1649977179
transform 1 0 33212 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1649977179
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_368
timestamp 1649977179
transform 1 0 34960 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_380
timestamp 1649977179
transform 1 0 36064 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_392
timestamp 1649977179
transform 1 0 37168 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_404
timestamp 1649977179
transform 1 0 38272 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_416
timestamp 1649977179
transform 1 0 39376 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_428
timestamp 1649977179
transform 1 0 40480 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_440
timestamp 1649977179
transform 1 0 41584 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_452
timestamp 1649977179
transform 1 0 42688 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_460
timestamp 1649977179
transform 1 0 43424 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_471
timestamp 1649977179
transform 1 0 44436 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1649977179
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_480
timestamp 1649977179
transform 1 0 45264 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_487
timestamp 1649977179
transform 1 0 45908 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_499
timestamp 1649977179
transform 1 0 47012 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1649977179
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_528
timestamp 1649977179
transform 1 0 49680 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_536
timestamp 1649977179
transform 1 0 50416 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_542
timestamp 1649977179
transform 1 0 50968 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_554
timestamp 1649977179
transform 1 0 52072 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_566
timestamp 1649977179
transform 1 0 53176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_578
timestamp 1649977179
transform 1 0 54280 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_586
timestamp 1649977179
transform 1 0 55016 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_625
timestamp 1649977179
transform 1 0 58604 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_637
timestamp 1649977179
transform 1 0 59708 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_643
timestamp 1649977179
transform 1 0 60260 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_645
timestamp 1649977179
transform 1 0 60444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_657
timestamp 1649977179
transform 1 0 61548 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_669
timestamp 1649977179
transform 1 0 62652 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_681
timestamp 1649977179
transform 1 0 63756 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_693
timestamp 1649977179
transform 1 0 64860 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_699
timestamp 1649977179
transform 1 0 65412 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_701
timestamp 1649977179
transform 1 0 65596 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_713
timestamp 1649977179
transform 1 0 66700 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_725
timestamp 1649977179
transform 1 0 67804 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_60
timestamp 1649977179
transform 1 0 6624 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_84
timestamp 1649977179
transform 1 0 8832 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_97
timestamp 1649977179
transform 1 0 10028 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_108
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_119
timestamp 1649977179
transform 1 0 12052 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_148
timestamp 1649977179
transform 1 0 14720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_171
timestamp 1649977179
transform 1 0 16836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_183
timestamp 1649977179
transform 1 0 17940 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_191
timestamp 1649977179
transform 1 0 18676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_213
timestamp 1649977179
transform 1 0 20700 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_231
timestamp 1649977179
transform 1 0 22356 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_258
timestamp 1649977179
transform 1 0 24840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_265
timestamp 1649977179
transform 1 0 25484 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_271
timestamp 1649977179
transform 1 0 26036 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1649977179
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_291
timestamp 1649977179
transform 1 0 27876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_297
timestamp 1649977179
transform 1 0 28428 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_303
timestamp 1649977179
transform 1 0 28980 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_315
timestamp 1649977179
transform 1 0 30084 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_323
timestamp 1649977179
transform 1 0 30820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1649977179
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_347
timestamp 1649977179
transform 1 0 33028 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_353
timestamp 1649977179
transform 1 0 33580 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_366
timestamp 1649977179
transform 1 0 34776 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_375
timestamp 1649977179
transform 1 0 35604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_387
timestamp 1649977179
transform 1 0 36708 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_397
timestamp 1649977179
transform 1 0 37628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_403
timestamp 1649977179
transform 1 0 38180 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_429
timestamp 1649977179
transform 1 0 40572 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_436
timestamp 1649977179
transform 1 0 41216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_443
timestamp 1649977179
transform 1 0 41860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1649977179
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_449
timestamp 1649977179
transform 1 0 42412 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_455
timestamp 1649977179
transform 1 0 42964 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_459
timestamp 1649977179
transform 1 0 43332 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_483
timestamp 1649977179
transform 1 0 45540 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_495
timestamp 1649977179
transform 1 0 46644 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1649977179
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_505
timestamp 1649977179
transform 1 0 47564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_509
timestamp 1649977179
transform 1 0 47932 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_516
timestamp 1649977179
transform 1 0 48576 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_532
timestamp 1649977179
transform 1 0 50048 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_544
timestamp 1649977179
transform 1 0 51152 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_556
timestamp 1649977179
transform 1 0 52256 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_561
timestamp 1649977179
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_573
timestamp 1649977179
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_585
timestamp 1649977179
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_597
timestamp 1649977179
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_609
timestamp 1649977179
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_615
timestamp 1649977179
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_629
timestamp 1649977179
transform 1 0 58972 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_641
timestamp 1649977179
transform 1 0 60076 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_653
timestamp 1649977179
transform 1 0 61180 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_665
timestamp 1649977179
transform 1 0 62284 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_671
timestamp 1649977179
transform 1 0 62836 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_673
timestamp 1649977179
transform 1 0 63020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_685
timestamp 1649977179
transform 1 0 64124 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_697
timestamp 1649977179
transform 1 0 65228 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_709
timestamp 1649977179
transform 1 0 66332 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_721
timestamp 1649977179
transform 1 0 67436 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_727
timestamp 1649977179
transform 1 0 67988 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_729
timestamp 1649977179
transform 1 0 68172 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_59
timestamp 1649977179
transform 1 0 6532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_71
timestamp 1649977179
transform 1 0 7636 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 1649977179
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_89
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_96
timestamp 1649977179
transform 1 0 9936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_102
timestamp 1649977179
transform 1 0 10488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_106
timestamp 1649977179
transform 1 0 10856 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_112
timestamp 1649977179
transform 1 0 11408 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_123
timestamp 1649977179
transform 1 0 12420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_130
timestamp 1649977179
transform 1 0 13064 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_144
timestamp 1649977179
transform 1 0 14352 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_157
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_167
timestamp 1649977179
transform 1 0 16468 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_174
timestamp 1649977179
transform 1 0 17112 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_182
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_200
timestamp 1649977179
transform 1 0 19504 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_220
timestamp 1649977179
transform 1 0 21344 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_231
timestamp 1649977179
transform 1 0 22356 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_239
timestamp 1649977179
transform 1 0 23092 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_257
timestamp 1649977179
transform 1 0 24748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_261
timestamp 1649977179
transform 1 0 25116 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_264
timestamp 1649977179
transform 1 0 25392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_270
timestamp 1649977179
transform 1 0 25944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_280
timestamp 1649977179
transform 1 0 26864 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_291
timestamp 1649977179
transform 1 0 27876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_299
timestamp 1649977179
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_311
timestamp 1649977179
transform 1 0 29716 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_317
timestamp 1649977179
transform 1 0 30268 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_343
timestamp 1649977179
transform 1 0 32660 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_349
timestamp 1649977179
transform 1 0 33212 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_359
timestamp 1649977179
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_372
timestamp 1649977179
transform 1 0 35328 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_379
timestamp 1649977179
transform 1 0 35972 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_391
timestamp 1649977179
transform 1 0 37076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_403
timestamp 1649977179
transform 1 0 38180 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_411
timestamp 1649977179
transform 1 0 38916 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1649977179
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_421
timestamp 1649977179
transform 1 0 39836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_425
timestamp 1649977179
transform 1 0 40204 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_431
timestamp 1649977179
transform 1 0 40756 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_437
timestamp 1649977179
transform 1 0 41308 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_446
timestamp 1649977179
transform 1 0 42136 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_458
timestamp 1649977179
transform 1 0 43240 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_462
timestamp 1649977179
transform 1 0 43608 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1649977179
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1649977179
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_480
timestamp 1649977179
transform 1 0 45264 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_492
timestamp 1649977179
transform 1 0 46368 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_504
timestamp 1649977179
transform 1 0 47472 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_512
timestamp 1649977179
transform 1 0 48208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_516
timestamp 1649977179
transform 1 0 48576 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_526
timestamp 1649977179
transform 1 0 49496 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_10_536
timestamp 1649977179
transform 1 0 50416 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_548
timestamp 1649977179
transform 1 0 51520 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_560
timestamp 1649977179
transform 1 0 52624 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_572
timestamp 1649977179
transform 1 0 53728 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_584
timestamp 1649977179
transform 1 0 54832 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_589
timestamp 1649977179
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_601
timestamp 1649977179
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_613
timestamp 1649977179
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_625
timestamp 1649977179
transform 1 0 58604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_637
timestamp 1649977179
transform 1 0 59708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_643
timestamp 1649977179
transform 1 0 60260 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_645
timestamp 1649977179
transform 1 0 60444 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_657
timestamp 1649977179
transform 1 0 61548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_669
timestamp 1649977179
transform 1 0 62652 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_681
timestamp 1649977179
transform 1 0 63756 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_693
timestamp 1649977179
transform 1 0 64860 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_699
timestamp 1649977179
transform 1 0 65412 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_701
timestamp 1649977179
transform 1 0 65596 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_713
timestamp 1649977179
transform 1 0 66700 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_725
timestamp 1649977179
transform 1 0 67804 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_48
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_66
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_72
timestamp 1649977179
transform 1 0 7728 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_80
timestamp 1649977179
transform 1 0 8464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_90
timestamp 1649977179
transform 1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1649977179
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_115
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp 1649977179
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_127
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_135
timestamp 1649977179
transform 1 0 13524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_138
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_147
timestamp 1649977179
transform 1 0 14628 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_158
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_185
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_197
timestamp 1649977179
transform 1 0 19228 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_201
timestamp 1649977179
transform 1 0 19596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_214
timestamp 1649977179
transform 1 0 20792 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1649977179
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_229
timestamp 1649977179
transform 1 0 22172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_233
timestamp 1649977179
transform 1 0 22540 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_244
timestamp 1649977179
transform 1 0 23552 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_250
timestamp 1649977179
transform 1 0 24104 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_253
timestamp 1649977179
transform 1 0 24380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_259
timestamp 1649977179
transform 1 0 24932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_269
timestamp 1649977179
transform 1 0 25852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_276
timestamp 1649977179
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_294
timestamp 1649977179
transform 1 0 28152 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_313
timestamp 1649977179
transform 1 0 29900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_319
timestamp 1649977179
transform 1 0 30452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_332
timestamp 1649977179
transform 1 0 31648 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_342
timestamp 1649977179
transform 1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_357
timestamp 1649977179
transform 1 0 33948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_365
timestamp 1649977179
transform 1 0 34684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_381
timestamp 1649977179
transform 1 0 36156 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_389
timestamp 1649977179
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_420
timestamp 1649977179
transform 1 0 39744 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_428
timestamp 1649977179
transform 1 0 40480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_439
timestamp 1649977179
transform 1 0 41492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1649977179
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_449
timestamp 1649977179
transform 1 0 42412 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_457
timestamp 1649977179
transform 1 0 43148 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_481
timestamp 1649977179
transform 1 0 45356 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_493
timestamp 1649977179
transform 1 0 46460 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_501
timestamp 1649977179
transform 1 0 47196 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1649977179
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_513
timestamp 1649977179
transform 1 0 48300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_519
timestamp 1649977179
transform 1 0 48852 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_529
timestamp 1649977179
transform 1 0 49772 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_538
timestamp 1649977179
transform 1 0 50600 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_550
timestamp 1649977179
transform 1 0 51704 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_558
timestamp 1649977179
transform 1 0 52440 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_561
timestamp 1649977179
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_573
timestamp 1649977179
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_585
timestamp 1649977179
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_597
timestamp 1649977179
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_609
timestamp 1649977179
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_615
timestamp 1649977179
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_617
timestamp 1649977179
transform 1 0 57868 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_629
timestamp 1649977179
transform 1 0 58972 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_641
timestamp 1649977179
transform 1 0 60076 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_653
timestamp 1649977179
transform 1 0 61180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_665
timestamp 1649977179
transform 1 0 62284 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_671
timestamp 1649977179
transform 1 0 62836 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_673
timestamp 1649977179
transform 1 0 63020 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_685
timestamp 1649977179
transform 1 0 64124 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_697
timestamp 1649977179
transform 1 0 65228 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_709
timestamp 1649977179
transform 1 0 66332 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_721
timestamp 1649977179
transform 1 0 67436 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_727
timestamp 1649977179
transform 1 0 67988 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_729
timestamp 1649977179
transform 1 0 68172 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1649977179
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_149
timestamp 1649977179
transform 1 0 14812 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_155
timestamp 1649977179
transform 1 0 15364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_176
timestamp 1649977179
transform 1 0 17296 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_182
timestamp 1649977179
transform 1 0 17848 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1649977179
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_215
timestamp 1649977179
transform 1 0 20884 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1649977179
transform 1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_234
timestamp 1649977179
transform 1 0 22632 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_246
timestamp 1649977179
transform 1 0 23736 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_259
timestamp 1649977179
transform 1 0 24932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_273
timestamp 1649977179
transform 1 0 26220 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_297
timestamp 1649977179
transform 1 0 28428 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1649977179
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_315
timestamp 1649977179
transform 1 0 30084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_335
timestamp 1649977179
transform 1 0 31924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_346
timestamp 1649977179
transform 1 0 32936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_353
timestamp 1649977179
transform 1 0 33580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_359
timestamp 1649977179
transform 1 0 34132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_393
timestamp 1649977179
transform 1 0 37260 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_405
timestamp 1649977179
transform 1 0 38364 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_417
timestamp 1649977179
transform 1 0 39468 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_421
timestamp 1649977179
transform 1 0 39836 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_442
timestamp 1649977179
transform 1 0 41768 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_454
timestamp 1649977179
transform 1 0 42872 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_466
timestamp 1649977179
transform 1 0 43976 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_471
timestamp 1649977179
transform 1 0 44436 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1649977179
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1649977179
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1649977179
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_501
timestamp 1649977179
transform 1 0 47196 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1649977179
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_525
timestamp 1649977179
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_531
timestamp 1649977179
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_539
timestamp 1649977179
transform 1 0 50692 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_548
timestamp 1649977179
transform 1 0 51520 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_560
timestamp 1649977179
transform 1 0 52624 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_572
timestamp 1649977179
transform 1 0 53728 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_584
timestamp 1649977179
transform 1 0 54832 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_589
timestamp 1649977179
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_601
timestamp 1649977179
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_613
timestamp 1649977179
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_625
timestamp 1649977179
transform 1 0 58604 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_637
timestamp 1649977179
transform 1 0 59708 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_643
timestamp 1649977179
transform 1 0 60260 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_645
timestamp 1649977179
transform 1 0 60444 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_657
timestamp 1649977179
transform 1 0 61548 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_669
timestamp 1649977179
transform 1 0 62652 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_681
timestamp 1649977179
transform 1 0 63756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_693
timestamp 1649977179
transform 1 0 64860 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_699
timestamp 1649977179
transform 1 0 65412 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_701
timestamp 1649977179
transform 1 0 65596 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_713
timestamp 1649977179
transform 1 0 66700 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_725
timestamp 1649977179
transform 1 0 67804 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_65
timestamp 1649977179
transform 1 0 7084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_92
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_104
timestamp 1649977179
transform 1 0 10672 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_157
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_176
timestamp 1649977179
transform 1 0 17296 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_188
timestamp 1649977179
transform 1 0 18400 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_200
timestamp 1649977179
transform 1 0 19504 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_208
timestamp 1649977179
transform 1 0 20240 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1649977179
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_231
timestamp 1649977179
transform 1 0 22356 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_243
timestamp 1649977179
transform 1 0 23460 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_255
timestamp 1649977179
transform 1 0 24564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_267
timestamp 1649977179
transform 1 0 25668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1649977179
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_283
timestamp 1649977179
transform 1 0 27140 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_13_299
timestamp 1649977179
transform 1 0 28612 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_308
timestamp 1649977179
transform 1 0 29440 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_314
timestamp 1649977179
transform 1 0 29992 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_327
timestamp 1649977179
transform 1 0 31188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_343
timestamp 1649977179
transform 1 0 32660 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_372
timestamp 1649977179
transform 1 0 35328 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1649977179
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_403
timestamp 1649977179
transform 1 0 38180 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_429
timestamp 1649977179
transform 1 0 40572 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_436
timestamp 1649977179
transform 1 0 41216 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1649977179
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_461
timestamp 1649977179
transform 1 0 43516 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_482
timestamp 1649977179
transform 1 0 45448 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_494
timestamp 1649977179
transform 1 0 46552 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_502
timestamp 1649977179
transform 1 0 47288 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_509
timestamp 1649977179
transform 1 0 47932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_523
timestamp 1649977179
transform 1 0 49220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_535
timestamp 1649977179
transform 1 0 50324 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_546
timestamp 1649977179
transform 1 0 51336 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1649977179
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1649977179
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_561
timestamp 1649977179
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_573
timestamp 1649977179
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_585
timestamp 1649977179
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_597
timestamp 1649977179
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_609
timestamp 1649977179
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_615
timestamp 1649977179
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_617
timestamp 1649977179
transform 1 0 57868 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_629
timestamp 1649977179
transform 1 0 58972 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_641
timestamp 1649977179
transform 1 0 60076 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_653
timestamp 1649977179
transform 1 0 61180 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_665
timestamp 1649977179
transform 1 0 62284 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_671
timestamp 1649977179
transform 1 0 62836 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_673
timestamp 1649977179
transform 1 0 63020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_685
timestamp 1649977179
transform 1 0 64124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_697
timestamp 1649977179
transform 1 0 65228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_709
timestamp 1649977179
transform 1 0 66332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_721
timestamp 1649977179
transform 1 0 67436 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_727
timestamp 1649977179
transform 1 0 67988 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_729
timestamp 1649977179
transform 1 0 68172 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_66
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_92
timestamp 1649977179
transform 1 0 9568 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_104
timestamp 1649977179
transform 1 0 10672 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_116
timestamp 1649977179
transform 1 0 11776 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_120
timestamp 1649977179
transform 1 0 12144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_143
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_155
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_178
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_184
timestamp 1649977179
transform 1 0 18032 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1649977179
transform 1 0 20424 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_220
timestamp 1649977179
transform 1 0 21344 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_238
timestamp 1649977179
transform 1 0 23000 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_244
timestamp 1649977179
transform 1 0 23552 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_260
timestamp 1649977179
transform 1 0 25024 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_266
timestamp 1649977179
transform 1 0 25576 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_273
timestamp 1649977179
transform 1 0 26220 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_285
timestamp 1649977179
transform 1 0 27324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_291
timestamp 1649977179
transform 1 0 27876 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_297
timestamp 1649977179
transform 1 0 28428 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_305
timestamp 1649977179
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_314
timestamp 1649977179
transform 1 0 29992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_322
timestamp 1649977179
transform 1 0 30728 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_326
timestamp 1649977179
transform 1 0 31096 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_329
timestamp 1649977179
transform 1 0 31372 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_346
timestamp 1649977179
transform 1 0 32936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_352
timestamp 1649977179
transform 1 0 33488 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_358
timestamp 1649977179
transform 1 0 34040 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_394
timestamp 1649977179
transform 1 0 37352 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_402
timestamp 1649977179
transform 1 0 38088 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_414
timestamp 1649977179
transform 1 0 39192 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_424
timestamp 1649977179
transform 1 0 40112 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_430
timestamp 1649977179
transform 1 0 40664 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_442
timestamp 1649977179
transform 1 0 41768 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_450
timestamp 1649977179
transform 1 0 42504 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_472
timestamp 1649977179
transform 1 0 44528 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_480
timestamp 1649977179
transform 1 0 45264 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_487
timestamp 1649977179
transform 1 0 45908 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_499
timestamp 1649977179
transform 1 0 47012 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_506
timestamp 1649977179
transform 1 0 47656 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_520
timestamp 1649977179
transform 1 0 48944 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_528
timestamp 1649977179
transform 1 0 49680 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_540
timestamp 1649977179
transform 1 0 50784 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_547
timestamp 1649977179
transform 1 0 51428 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_559
timestamp 1649977179
transform 1 0 52532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_571
timestamp 1649977179
transform 1 0 53636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_583
timestamp 1649977179
transform 1 0 54740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1649977179
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_589
timestamp 1649977179
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_601
timestamp 1649977179
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_613
timestamp 1649977179
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_625
timestamp 1649977179
transform 1 0 58604 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_637
timestamp 1649977179
transform 1 0 59708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_643
timestamp 1649977179
transform 1 0 60260 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_645
timestamp 1649977179
transform 1 0 60444 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_657
timestamp 1649977179
transform 1 0 61548 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_669
timestamp 1649977179
transform 1 0 62652 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_681
timestamp 1649977179
transform 1 0 63756 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_693
timestamp 1649977179
transform 1 0 64860 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_699
timestamp 1649977179
transform 1 0 65412 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_701
timestamp 1649977179
transform 1 0 65596 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_713
timestamp 1649977179
transform 1 0 66700 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_725
timestamp 1649977179
transform 1 0 67804 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_43
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_47
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_66
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_72
timestamp 1649977179
transform 1 0 7728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_80
timestamp 1649977179
transform 1 0 8464 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_86
timestamp 1649977179
transform 1 0 9016 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_98
timestamp 1649977179
transform 1 0 10120 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_133
timestamp 1649977179
transform 1 0 13340 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_144
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_152
timestamp 1649977179
transform 1 0 15088 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_172
timestamp 1649977179
transform 1 0 16928 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_184
timestamp 1649977179
transform 1 0 18032 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_196
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_208
timestamp 1649977179
transform 1 0 20240 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_216
timestamp 1649977179
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_227
timestamp 1649977179
transform 1 0 21988 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_239
timestamp 1649977179
transform 1 0 23092 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_251
timestamp 1649977179
transform 1 0 24196 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_259
timestamp 1649977179
transform 1 0 24932 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_262
timestamp 1649977179
transform 1 0 25208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_266
timestamp 1649977179
transform 1 0 25576 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1649977179
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_301
timestamp 1649977179
transform 1 0 28796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_311
timestamp 1649977179
transform 1 0 29716 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_319
timestamp 1649977179
transform 1 0 30452 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_327
timestamp 1649977179
transform 1 0 31188 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_343
timestamp 1649977179
transform 1 0 32660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_347
timestamp 1649977179
transform 1 0 33028 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_357
timestamp 1649977179
transform 1 0 33948 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_369
timestamp 1649977179
transform 1 0 35052 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_381
timestamp 1649977179
transform 1 0 36156 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_389
timestamp 1649977179
transform 1 0 36892 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_408
timestamp 1649977179
transform 1 0 38640 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_418
timestamp 1649977179
transform 1 0 39560 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_426
timestamp 1649977179
transform 1 0 40296 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_433
timestamp 1649977179
transform 1 0 40940 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_439
timestamp 1649977179
transform 1 0 41492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1649977179
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_453
timestamp 1649977179
transform 1 0 42780 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_459
timestamp 1649977179
transform 1 0 43332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_463
timestamp 1649977179
transform 1 0 43700 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_484
timestamp 1649977179
transform 1 0 45632 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_496
timestamp 1649977179
transform 1 0 46736 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1649977179
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_510
timestamp 1649977179
transform 1 0 48024 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_520
timestamp 1649977179
transform 1 0 48944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_534
timestamp 1649977179
transform 1 0 50232 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_541
timestamp 1649977179
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_553
timestamp 1649977179
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_559
timestamp 1649977179
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_561
timestamp 1649977179
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_573
timestamp 1649977179
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_585
timestamp 1649977179
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_597
timestamp 1649977179
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_609
timestamp 1649977179
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_615
timestamp 1649977179
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_617
timestamp 1649977179
transform 1 0 57868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_629
timestamp 1649977179
transform 1 0 58972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_641
timestamp 1649977179
transform 1 0 60076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_653
timestamp 1649977179
transform 1 0 61180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_665
timestamp 1649977179
transform 1 0 62284 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_671
timestamp 1649977179
transform 1 0 62836 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_673
timestamp 1649977179
transform 1 0 63020 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_685
timestamp 1649977179
transform 1 0 64124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_697
timestamp 1649977179
transform 1 0 65228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_709
timestamp 1649977179
transform 1 0 66332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_721
timestamp 1649977179
transform 1 0 67436 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_727
timestamp 1649977179
transform 1 0 67988 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_729
timestamp 1649977179
transform 1 0 68172 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_37
timestamp 1649977179
transform 1 0 4508 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_16_56
timestamp 1649977179
transform 1 0 6256 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 1649977179
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_79
timestamp 1649977179
transform 1 0 8372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_92
timestamp 1649977179
transform 1 0 9568 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_104
timestamp 1649977179
transform 1 0 10672 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_108
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_111
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_119
timestamp 1649977179
transform 1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_130
timestamp 1649977179
transform 1 0 13064 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_152
timestamp 1649977179
transform 1 0 15088 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_170
timestamp 1649977179
transform 1 0 16744 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_179
timestamp 1649977179
transform 1 0 17572 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_187
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_206
timestamp 1649977179
transform 1 0 20056 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_216
timestamp 1649977179
transform 1 0 20976 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_226
timestamp 1649977179
transform 1 0 21896 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_232
timestamp 1649977179
transform 1 0 22448 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_257
timestamp 1649977179
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_264
timestamp 1649977179
transform 1 0 25392 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_270
timestamp 1649977179
transform 1 0 25944 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_276
timestamp 1649977179
transform 1 0 26496 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_282
timestamp 1649977179
transform 1 0 27048 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_290
timestamp 1649977179
transform 1 0 27784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_298
timestamp 1649977179
transform 1 0 28520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1649977179
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_315
timestamp 1649977179
transform 1 0 30084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_319
timestamp 1649977179
transform 1 0 30452 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_329
timestamp 1649977179
transform 1 0 31372 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_349
timestamp 1649977179
transform 1 0 33212 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_356
timestamp 1649977179
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_383
timestamp 1649977179
transform 1 0 36340 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_396
timestamp 1649977179
transform 1 0 37536 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_402
timestamp 1649977179
transform 1 0 38088 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_416
timestamp 1649977179
transform 1 0 39376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_441
timestamp 1649977179
transform 1 0 41676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_449
timestamp 1649977179
transform 1 0 42412 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_457
timestamp 1649977179
transform 1 0 43148 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_465
timestamp 1649977179
transform 1 0 43884 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_472
timestamp 1649977179
transform 1 0 44528 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_497
timestamp 1649977179
transform 1 0 46828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_504
timestamp 1649977179
transform 1 0 47472 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_513
timestamp 1649977179
transform 1 0 48300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_522
timestamp 1649977179
transform 1 0 49128 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_530
timestamp 1649977179
transform 1 0 49864 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_538
timestamp 1649977179
transform 1 0 50600 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_550
timestamp 1649977179
transform 1 0 51704 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_562
timestamp 1649977179
transform 1 0 52808 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_574
timestamp 1649977179
transform 1 0 53912 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_586
timestamp 1649977179
transform 1 0 55016 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_589
timestamp 1649977179
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_601
timestamp 1649977179
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_613
timestamp 1649977179
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_625
timestamp 1649977179
transform 1 0 58604 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_637
timestamp 1649977179
transform 1 0 59708 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_643
timestamp 1649977179
transform 1 0 60260 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_645
timestamp 1649977179
transform 1 0 60444 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_657
timestamp 1649977179
transform 1 0 61548 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_669
timestamp 1649977179
transform 1 0 62652 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_681
timestamp 1649977179
transform 1 0 63756 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_693
timestamp 1649977179
transform 1 0 64860 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_699
timestamp 1649977179
transform 1 0 65412 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_701
timestamp 1649977179
transform 1 0 65596 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_713
timestamp 1649977179
transform 1 0 66700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_717
timestamp 1649977179
transform 1 0 67068 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_721
timestamp 1649977179
transform 1 0 67436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_727
timestamp 1649977179
transform 1 0 67988 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp 1649977179
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 1649977179
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_68
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_79
timestamp 1649977179
transform 1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_86
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_98
timestamp 1649977179
transform 1 0 10120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_130
timestamp 1649977179
transform 1 0 13064 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_138
timestamp 1649977179
transform 1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_153
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_157
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_175
timestamp 1649977179
transform 1 0 17204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1649977179
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 1649977179
transform 1 0 20056 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_258
timestamp 1649977179
transform 1 0 24840 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_269
timestamp 1649977179
transform 1 0 25852 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1649977179
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_284
timestamp 1649977179
transform 1 0 27232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_290
timestamp 1649977179
transform 1 0 27784 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_298
timestamp 1649977179
transform 1 0 28520 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_307
timestamp 1649977179
transform 1 0 29348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_331
timestamp 1649977179
transform 1 0 31556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_341
timestamp 1649977179
transform 1 0 32476 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_345
timestamp 1649977179
transform 1 0 32844 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_365
timestamp 1649977179
transform 1 0 34684 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_397
timestamp 1649977179
transform 1 0 37628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_421
timestamp 1649977179
transform 1 0 39836 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_428
timestamp 1649977179
transform 1 0 40480 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_440
timestamp 1649977179
transform 1 0 41584 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_451
timestamp 1649977179
transform 1 0 42596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_457
timestamp 1649977179
transform 1 0 43148 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_485
timestamp 1649977179
transform 1 0 45724 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_492
timestamp 1649977179
transform 1 0 46368 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_505
timestamp 1649977179
transform 1 0 47564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_517
timestamp 1649977179
transform 1 0 48668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_526
timestamp 1649977179
transform 1 0 49496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_534
timestamp 1649977179
transform 1 0 50232 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_541
timestamp 1649977179
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_553
timestamp 1649977179
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_559
timestamp 1649977179
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_561
timestamp 1649977179
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_573
timestamp 1649977179
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_585
timestamp 1649977179
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_597
timestamp 1649977179
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_609
timestamp 1649977179
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1649977179
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_617
timestamp 1649977179
transform 1 0 57868 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_629
timestamp 1649977179
transform 1 0 58972 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_641
timestamp 1649977179
transform 1 0 60076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_653
timestamp 1649977179
transform 1 0 61180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_665
timestamp 1649977179
transform 1 0 62284 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_671
timestamp 1649977179
transform 1 0 62836 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_673
timestamp 1649977179
transform 1 0 63020 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_685
timestamp 1649977179
transform 1 0 64124 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_697
timestamp 1649977179
transform 1 0 65228 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_709
timestamp 1649977179
transform 1 0 66332 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_717
timestamp 1649977179
transform 1 0 67068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_724
timestamp 1649977179
transform 1 0 67712 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_729
timestamp 1649977179
transform 1 0 68172 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_57
timestamp 1649977179
transform 1 0 6348 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp 1649977179
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_94
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_106
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_117
timestamp 1649977179
transform 1 0 11868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_125
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_128
timestamp 1649977179
transform 1 0 12880 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_132
timestamp 1649977179
transform 1 0 13248 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1649977179
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_149
timestamp 1649977179
transform 1 0 14812 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_155
timestamp 1649977179
transform 1 0 15364 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_158
timestamp 1649977179
transform 1 0 15640 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_171
timestamp 1649977179
transform 1 0 16836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_183
timestamp 1649977179
transform 1 0 17940 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_200
timestamp 1649977179
transform 1 0 19504 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_204
timestamp 1649977179
transform 1 0 19872 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_211
timestamp 1649977179
transform 1 0 20516 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_218
timestamp 1649977179
transform 1 0 21160 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_224
timestamp 1649977179
transform 1 0 21712 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_227
timestamp 1649977179
transform 1 0 21988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_239
timestamp 1649977179
transform 1 0 23092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_256
timestamp 1649977179
transform 1 0 24656 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_283
timestamp 1649977179
transform 1 0 27140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_295
timestamp 1649977179
transform 1 0 28244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_329
timestamp 1649977179
transform 1 0 31372 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_348
timestamp 1649977179
transform 1 0 33120 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_354
timestamp 1649977179
transform 1 0 33672 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_362
timestamp 1649977179
transform 1 0 34408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_375
timestamp 1649977179
transform 1 0 35604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_386
timestamp 1649977179
transform 1 0 36616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_402
timestamp 1649977179
transform 1 0 38088 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_411
timestamp 1649977179
transform 1 0 38916 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1649977179
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_423
timestamp 1649977179
transform 1 0 40020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_429
timestamp 1649977179
transform 1 0 40572 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_437
timestamp 1649977179
transform 1 0 41308 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_449
timestamp 1649977179
transform 1 0 42412 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_461
timestamp 1649977179
transform 1 0 43516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_473
timestamp 1649977179
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_480
timestamp 1649977179
transform 1 0 45264 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_492
timestamp 1649977179
transform 1 0 46368 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_504
timestamp 1649977179
transform 1 0 47472 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_513
timestamp 1649977179
transform 1 0 48300 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_522
timestamp 1649977179
transform 1 0 49128 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_530
timestamp 1649977179
transform 1 0 49864 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_533
timestamp 1649977179
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_545
timestamp 1649977179
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_557
timestamp 1649977179
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_569
timestamp 1649977179
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1649977179
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1649977179
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_589
timestamp 1649977179
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_601
timestamp 1649977179
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_613
timestamp 1649977179
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_625
timestamp 1649977179
transform 1 0 58604 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_637
timestamp 1649977179
transform 1 0 59708 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_643
timestamp 1649977179
transform 1 0 60260 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_645
timestamp 1649977179
transform 1 0 60444 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_657
timestamp 1649977179
transform 1 0 61548 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_669
timestamp 1649977179
transform 1 0 62652 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_681
timestamp 1649977179
transform 1 0 63756 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_693
timestamp 1649977179
transform 1 0 64860 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_699
timestamp 1649977179
transform 1 0 65412 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_701
timestamp 1649977179
transform 1 0 65596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_713
timestamp 1649977179
transform 1 0 66700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_725
timestamp 1649977179
transform 1 0 67804 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_35
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_38
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_64
timestamp 1649977179
transform 1 0 6992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_75
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_88
timestamp 1649977179
transform 1 0 9200 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_94
timestamp 1649977179
transform 1 0 9752 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_116
timestamp 1649977179
transform 1 0 11776 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_126
timestamp 1649977179
transform 1 0 12696 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_134
timestamp 1649977179
transform 1 0 13432 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_144
timestamp 1649977179
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_148
timestamp 1649977179
transform 1 0 14720 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_156
timestamp 1649977179
transform 1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_160
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_186
timestamp 1649977179
transform 1 0 18216 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_196
timestamp 1649977179
transform 1 0 19136 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_207
timestamp 1649977179
transform 1 0 20148 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_214
timestamp 1649977179
transform 1 0 20792 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_236
timestamp 1649977179
transform 1 0 22816 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_248
timestamp 1649977179
transform 1 0 23920 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_256
timestamp 1649977179
transform 1 0 24656 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_259
timestamp 1649977179
transform 1 0 24932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_270
timestamp 1649977179
transform 1 0 25944 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1649977179
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_290
timestamp 1649977179
transform 1 0 27784 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_301
timestamp 1649977179
transform 1 0 28796 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_313
timestamp 1649977179
transform 1 0 29900 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_325
timestamp 1649977179
transform 1 0 31004 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1649977179
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_341
timestamp 1649977179
transform 1 0 32476 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_344
timestamp 1649977179
transform 1 0 32752 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_357
timestamp 1649977179
transform 1 0 33948 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_369
timestamp 1649977179
transform 1 0 35052 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_377
timestamp 1649977179
transform 1 0 35788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1649977179
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_400
timestamp 1649977179
transform 1 0 37904 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_408
timestamp 1649977179
transform 1 0 38640 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_420
timestamp 1649977179
transform 1 0 39744 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_427
timestamp 1649977179
transform 1 0 40388 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_439
timestamp 1649977179
transform 1 0 41492 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1649977179
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_449
timestamp 1649977179
transform 1 0 42412 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_459
timestamp 1649977179
transform 1 0 43332 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_465
timestamp 1649977179
transform 1 0 43884 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_477
timestamp 1649977179
transform 1 0 44988 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_489
timestamp 1649977179
transform 1 0 46092 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_501
timestamp 1649977179
transform 1 0 47196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1649977179
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1649977179
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_520
timestamp 1649977179
transform 1 0 48944 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_527
timestamp 1649977179
transform 1 0 49588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_539
timestamp 1649977179
transform 1 0 50692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_551
timestamp 1649977179
transform 1 0 51796 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1649977179
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_561
timestamp 1649977179
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_573
timestamp 1649977179
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_585
timestamp 1649977179
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_597
timestamp 1649977179
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1649977179
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1649977179
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_617
timestamp 1649977179
transform 1 0 57868 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_629
timestamp 1649977179
transform 1 0 58972 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_641
timestamp 1649977179
transform 1 0 60076 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_653
timestamp 1649977179
transform 1 0 61180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_665
timestamp 1649977179
transform 1 0 62284 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_671
timestamp 1649977179
transform 1 0 62836 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_673
timestamp 1649977179
transform 1 0 63020 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_685
timestamp 1649977179
transform 1 0 64124 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_697
timestamp 1649977179
transform 1 0 65228 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_709
timestamp 1649977179
transform 1 0 66332 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_721
timestamp 1649977179
transform 1 0 67436 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_727
timestamp 1649977179
transform 1 0 67988 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_729
timestamp 1649977179
transform 1 0 68172 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_37
timestamp 1649977179
transform 1 0 4508 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_55
timestamp 1649977179
transform 1 0 6164 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_101
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_118
timestamp 1649977179
transform 1 0 11960 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_149
timestamp 1649977179
transform 1 0 14812 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_157
timestamp 1649977179
transform 1 0 15548 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_161
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_168
timestamp 1649977179
transform 1 0 16560 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_174
timestamp 1649977179
transform 1 0 17112 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_188
timestamp 1649977179
transform 1 0 18400 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_217
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_238
timestamp 1649977179
transform 1 0 23000 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_244
timestamp 1649977179
transform 1 0 23552 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_268
timestamp 1649977179
transform 1 0 25760 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_288
timestamp 1649977179
transform 1 0 27600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_295
timestamp 1649977179
transform 1 0 28244 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1649977179
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_316
timestamp 1649977179
transform 1 0 30176 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_328
timestamp 1649977179
transform 1 0 31280 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_334
timestamp 1649977179
transform 1 0 31832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_342
timestamp 1649977179
transform 1 0 32568 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_355
timestamp 1649977179
transform 1 0 33764 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_383
timestamp 1649977179
transform 1 0 36340 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_388
timestamp 1649977179
transform 1 0 36800 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_398
timestamp 1649977179
transform 1 0 37720 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_402
timestamp 1649977179
transform 1 0 38088 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_407
timestamp 1649977179
transform 1 0 38548 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_414
timestamp 1649977179
transform 1 0 39192 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_423
timestamp 1649977179
transform 1 0 40020 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_435
timestamp 1649977179
transform 1 0 41124 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_441
timestamp 1649977179
transform 1 0 41676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_452
timestamp 1649977179
transform 1 0 42688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_462
timestamp 1649977179
transform 1 0 43608 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1649977179
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1649977179
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1649977179
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1649977179
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1649977179
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1649977179
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1649977179
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1649977179
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_533
timestamp 1649977179
transform 1 0 50140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_545
timestamp 1649977179
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_557
timestamp 1649977179
transform 1 0 52348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_569
timestamp 1649977179
transform 1 0 53452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_581
timestamp 1649977179
transform 1 0 54556 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_587
timestamp 1649977179
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_589
timestamp 1649977179
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_601
timestamp 1649977179
transform 1 0 56396 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_613
timestamp 1649977179
transform 1 0 57500 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_625
timestamp 1649977179
transform 1 0 58604 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_637
timestamp 1649977179
transform 1 0 59708 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_643
timestamp 1649977179
transform 1 0 60260 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_645
timestamp 1649977179
transform 1 0 60444 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_657
timestamp 1649977179
transform 1 0 61548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_669
timestamp 1649977179
transform 1 0 62652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_681
timestamp 1649977179
transform 1 0 63756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_693
timestamp 1649977179
transform 1 0 64860 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_699
timestamp 1649977179
transform 1 0 65412 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_701
timestamp 1649977179
transform 1 0 65596 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_713
timestamp 1649977179
transform 1 0 66700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_725
timestamp 1649977179
transform 1 0 67804 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_42
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_67
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_73
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_85
timestamp 1649977179
transform 1 0 8924 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1649977179
transform 1 0 10028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_106
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_122
timestamp 1649977179
transform 1 0 12328 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_128
timestamp 1649977179
transform 1 0 12880 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_134
timestamp 1649977179
transform 1 0 13432 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_143
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_156
timestamp 1649977179
transform 1 0 15456 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_171
timestamp 1649977179
transform 1 0 16836 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_183
timestamp 1649977179
transform 1 0 17940 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_188
timestamp 1649977179
transform 1 0 18400 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_194
timestamp 1649977179
transform 1 0 18952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_201
timestamp 1649977179
transform 1 0 19596 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_212
timestamp 1649977179
transform 1 0 20608 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1649977179
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_228
timestamp 1649977179
transform 1 0 22080 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_236
timestamp 1649977179
transform 1 0 22816 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_246
timestamp 1649977179
transform 1 0 23736 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_258
timestamp 1649977179
transform 1 0 24840 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_268
timestamp 1649977179
transform 1 0 25760 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1649977179
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_285
timestamp 1649977179
transform 1 0 27324 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_296
timestamp 1649977179
transform 1 0 28336 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_308
timestamp 1649977179
transform 1 0 29440 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_320
timestamp 1649977179
transform 1 0 30544 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1649977179
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_345
timestamp 1649977179
transform 1 0 32844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_364
timestamp 1649977179
transform 1 0 34592 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_372
timestamp 1649977179
transform 1 0 35328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_377
timestamp 1649977179
transform 1 0 35788 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_384
timestamp 1649977179
transform 1 0 36432 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_400
timestamp 1649977179
transform 1 0 37904 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_21_422
timestamp 1649977179
transform 1 0 39928 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_432
timestamp 1649977179
transform 1 0 40848 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_440
timestamp 1649977179
transform 1 0 41584 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_444
timestamp 1649977179
transform 1 0 41952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_465
timestamp 1649977179
transform 1 0 43884 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_475
timestamp 1649977179
transform 1 0 44804 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_481
timestamp 1649977179
transform 1 0 45356 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_493
timestamp 1649977179
transform 1 0 46460 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_501
timestamp 1649977179
transform 1 0 47196 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1649977179
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_517
timestamp 1649977179
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_529
timestamp 1649977179
transform 1 0 49772 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_541
timestamp 1649977179
transform 1 0 50876 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_553
timestamp 1649977179
transform 1 0 51980 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_559
timestamp 1649977179
transform 1 0 52532 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_561
timestamp 1649977179
transform 1 0 52716 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_573
timestamp 1649977179
transform 1 0 53820 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_585
timestamp 1649977179
transform 1 0 54924 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_597
timestamp 1649977179
transform 1 0 56028 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_609
timestamp 1649977179
transform 1 0 57132 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1649977179
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_617
timestamp 1649977179
transform 1 0 57868 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_629
timestamp 1649977179
transform 1 0 58972 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_641
timestamp 1649977179
transform 1 0 60076 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_653
timestamp 1649977179
transform 1 0 61180 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_665
timestamp 1649977179
transform 1 0 62284 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_671
timestamp 1649977179
transform 1 0 62836 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_673
timestamp 1649977179
transform 1 0 63020 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_685
timestamp 1649977179
transform 1 0 64124 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_697
timestamp 1649977179
transform 1 0 65228 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_709
timestamp 1649977179
transform 1 0 66332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_721
timestamp 1649977179
transform 1 0 67436 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_727
timestamp 1649977179
transform 1 0 67988 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_729
timestamp 1649977179
transform 1 0 68172 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_60
timestamp 1649977179
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_64
timestamp 1649977179
transform 1 0 6992 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_67
timestamp 1649977179
transform 1 0 7268 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_75
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_99
timestamp 1649977179
transform 1 0 10212 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_111
timestamp 1649977179
transform 1 0 11316 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_119
timestamp 1649977179
transform 1 0 12052 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_124
timestamp 1649977179
transform 1 0 12512 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1649977179
transform 1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_160
timestamp 1649977179
transform 1 0 15824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_167
timestamp 1649977179
transform 1 0 16468 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1649977179
transform 1 0 17112 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_181
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1649977179
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_206
timestamp 1649977179
transform 1 0 20056 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_214
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_229
timestamp 1649977179
transform 1 0 22172 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_234
timestamp 1649977179
transform 1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_238
timestamp 1649977179
transform 1 0 23000 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_242
timestamp 1649977179
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1649977179
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_273
timestamp 1649977179
transform 1 0 26220 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_276
timestamp 1649977179
transform 1 0 26496 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_282
timestamp 1649977179
transform 1 0 27048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1649977179
transform 1 0 27600 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_296
timestamp 1649977179
transform 1 0 28336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1649977179
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_313
timestamp 1649977179
transform 1 0 29900 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_325
timestamp 1649977179
transform 1 0 31004 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_341
timestamp 1649977179
transform 1 0 32476 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_347
timestamp 1649977179
transform 1 0 33028 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_351
timestamp 1649977179
transform 1 0 33396 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_394
timestamp 1649977179
transform 1 0 37352 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_407
timestamp 1649977179
transform 1 0 38548 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_416
timestamp 1649977179
transform 1 0 39376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_428
timestamp 1649977179
transform 1 0 40480 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_438
timestamp 1649977179
transform 1 0 41400 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_455
timestamp 1649977179
transform 1 0 42964 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_468
timestamp 1649977179
transform 1 0 44160 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_22_490
timestamp 1649977179
transform 1 0 46184 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_502
timestamp 1649977179
transform 1 0 47288 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_514
timestamp 1649977179
transform 1 0 48392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_526
timestamp 1649977179
transform 1 0 49496 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_533
timestamp 1649977179
transform 1 0 50140 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_545
timestamp 1649977179
transform 1 0 51244 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_557
timestamp 1649977179
transform 1 0 52348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_569
timestamp 1649977179
transform 1 0 53452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_581
timestamp 1649977179
transform 1 0 54556 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_587
timestamp 1649977179
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_589
timestamp 1649977179
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_601
timestamp 1649977179
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_613
timestamp 1649977179
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_625
timestamp 1649977179
transform 1 0 58604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_637
timestamp 1649977179
transform 1 0 59708 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_643
timestamp 1649977179
transform 1 0 60260 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_645
timestamp 1649977179
transform 1 0 60444 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_657
timestamp 1649977179
transform 1 0 61548 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_669
timestamp 1649977179
transform 1 0 62652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_681
timestamp 1649977179
transform 1 0 63756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_693
timestamp 1649977179
transform 1 0 64860 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_699
timestamp 1649977179
transform 1 0 65412 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_701
timestamp 1649977179
transform 1 0 65596 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_713
timestamp 1649977179
transform 1 0 66700 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_725
timestamp 1649977179
transform 1 0 67804 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_75
timestamp 1649977179
transform 1 0 8004 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_87
timestamp 1649977179
transform 1 0 9108 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1649977179
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_115
timestamp 1649977179
transform 1 0 11684 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1649977179
transform 1 0 12236 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_140
timestamp 1649977179
transform 1 0 13984 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_147
timestamp 1649977179
transform 1 0 14628 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1649977179
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_177
timestamp 1649977179
transform 1 0 17388 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_201
timestamp 1649977179
transform 1 0 19596 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_213
timestamp 1649977179
transform 1 0 20700 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1649977179
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_230
timestamp 1649977179
transform 1 0 22264 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_254
timestamp 1649977179
transform 1 0 24472 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1649977179
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_286
timestamp 1649977179
transform 1 0 27416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_299
timestamp 1649977179
transform 1 0 28612 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_313
timestamp 1649977179
transform 1 0 29900 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_324
timestamp 1649977179
transform 1 0 30912 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_341
timestamp 1649977179
transform 1 0 32476 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_354
timestamp 1649977179
transform 1 0 33672 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_362
timestamp 1649977179
transform 1 0 34408 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_374
timestamp 1649977179
transform 1 0 35512 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_388
timestamp 1649977179
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_399
timestamp 1649977179
transform 1 0 37812 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_415
timestamp 1649977179
transform 1 0 39284 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_428
timestamp 1649977179
transform 1 0 40480 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_440
timestamp 1649977179
transform 1 0 41584 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_449
timestamp 1649977179
transform 1 0 42412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_453
timestamp 1649977179
transform 1 0 42780 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_460
timestamp 1649977179
transform 1 0 43424 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_480
timestamp 1649977179
transform 1 0 45264 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_486
timestamp 1649977179
transform 1 0 45816 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_498
timestamp 1649977179
transform 1 0 46920 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1649977179
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_517
timestamp 1649977179
transform 1 0 48668 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_529
timestamp 1649977179
transform 1 0 49772 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_541
timestamp 1649977179
transform 1 0 50876 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_553
timestamp 1649977179
transform 1 0 51980 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_559
timestamp 1649977179
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_561
timestamp 1649977179
transform 1 0 52716 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_573
timestamp 1649977179
transform 1 0 53820 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_585
timestamp 1649977179
transform 1 0 54924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_597
timestamp 1649977179
transform 1 0 56028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_609
timestamp 1649977179
transform 1 0 57132 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_615
timestamp 1649977179
transform 1 0 57684 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_617
timestamp 1649977179
transform 1 0 57868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_629
timestamp 1649977179
transform 1 0 58972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_641
timestamp 1649977179
transform 1 0 60076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_653
timestamp 1649977179
transform 1 0 61180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_665
timestamp 1649977179
transform 1 0 62284 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_671
timestamp 1649977179
transform 1 0 62836 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_673
timestamp 1649977179
transform 1 0 63020 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_685
timestamp 1649977179
transform 1 0 64124 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_697
timestamp 1649977179
transform 1 0 65228 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_709
timestamp 1649977179
transform 1 0 66332 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_721
timestamp 1649977179
transform 1 0 67436 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_727
timestamp 1649977179
transform 1 0 67988 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_729
timestamp 1649977179
transform 1 0 68172 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_47
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_67
timestamp 1649977179
transform 1 0 7268 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 1649977179
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_95
timestamp 1649977179
transform 1 0 9844 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_108
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_128
timestamp 1649977179
transform 1 0 12880 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_144
timestamp 1649977179
transform 1 0 14352 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_164
timestamp 1649977179
transform 1 0 16192 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_168
timestamp 1649977179
transform 1 0 16560 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1649977179
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_184
timestamp 1649977179
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_199
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_211
timestamp 1649977179
transform 1 0 20516 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_223
timestamp 1649977179
transform 1 0 21620 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_226
timestamp 1649977179
transform 1 0 21896 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_239
timestamp 1649977179
transform 1 0 23092 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_248
timestamp 1649977179
transform 1 0 23920 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_258
timestamp 1649977179
transform 1 0 24840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_270
timestamp 1649977179
transform 1 0 25944 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_273
timestamp 1649977179
transform 1 0 26220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_284
timestamp 1649977179
transform 1 0 27232 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_292
timestamp 1649977179
transform 1 0 27968 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_299
timestamp 1649977179
transform 1 0 28612 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_316
timestamp 1649977179
transform 1 0 30176 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_328
timestamp 1649977179
transform 1 0 31280 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_336
timestamp 1649977179
transform 1 0 32016 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_353
timestamp 1649977179
transform 1 0 33580 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_361
timestamp 1649977179
transform 1 0 34316 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_413
timestamp 1649977179
transform 1 0 39100 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_416
timestamp 1649977179
transform 1 0 39376 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_427
timestamp 1649977179
transform 1 0 40388 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_435
timestamp 1649977179
transform 1 0 41124 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_443
timestamp 1649977179
transform 1 0 41860 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_449
timestamp 1649977179
transform 1 0 42412 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_24_459
timestamp 1649977179
transform 1 0 43332 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_472
timestamp 1649977179
transform 1 0 44528 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1649977179
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1649977179
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1649977179
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1649977179
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_525
timestamp 1649977179
transform 1 0 49404 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_531
timestamp 1649977179
transform 1 0 49956 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_533
timestamp 1649977179
transform 1 0 50140 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_545
timestamp 1649977179
transform 1 0 51244 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_557
timestamp 1649977179
transform 1 0 52348 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_569
timestamp 1649977179
transform 1 0 53452 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_581
timestamp 1649977179
transform 1 0 54556 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_587
timestamp 1649977179
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_589
timestamp 1649977179
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_601
timestamp 1649977179
transform 1 0 56396 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_613
timestamp 1649977179
transform 1 0 57500 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_625
timestamp 1649977179
transform 1 0 58604 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_637
timestamp 1649977179
transform 1 0 59708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_643
timestamp 1649977179
transform 1 0 60260 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_645
timestamp 1649977179
transform 1 0 60444 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_657
timestamp 1649977179
transform 1 0 61548 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_669
timestamp 1649977179
transform 1 0 62652 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_681
timestamp 1649977179
transform 1 0 63756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_693
timestamp 1649977179
transform 1 0 64860 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_699
timestamp 1649977179
transform 1 0 65412 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_701
timestamp 1649977179
transform 1 0 65596 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_713
timestamp 1649977179
transform 1 0 66700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_725
timestamp 1649977179
transform 1 0 67804 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_35
timestamp 1649977179
transform 1 0 4324 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1649977179
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_77
timestamp 1649977179
transform 1 0 8188 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_83
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_95
timestamp 1649977179
transform 1 0 9844 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_108
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_128
timestamp 1649977179
transform 1 0 12880 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_134
timestamp 1649977179
transform 1 0 13432 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_144
timestamp 1649977179
transform 1 0 14352 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_150
timestamp 1649977179
transform 1 0 14904 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1649977179
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_175
timestamp 1649977179
transform 1 0 17204 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_187
timestamp 1649977179
transform 1 0 18308 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_230
timestamp 1649977179
transform 1 0 22264 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_236
timestamp 1649977179
transform 1 0 22816 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_244
timestamp 1649977179
transform 1 0 23552 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_252
timestamp 1649977179
transform 1 0 24288 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_262
timestamp 1649977179
transform 1 0 25208 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_268
timestamp 1649977179
transform 1 0 25760 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_290
timestamp 1649977179
transform 1 0 27784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_297
timestamp 1649977179
transform 1 0 28428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_303
timestamp 1649977179
transform 1 0 28980 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_307
timestamp 1649977179
transform 1 0 29348 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1649977179
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_348
timestamp 1649977179
transform 1 0 33120 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_354
timestamp 1649977179
transform 1 0 33672 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_358
timestamp 1649977179
transform 1 0 34040 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_369
timestamp 1649977179
transform 1 0 35052 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_381
timestamp 1649977179
transform 1 0 36156 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_389
timestamp 1649977179
transform 1 0 36892 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1649977179
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1649977179
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1649977179
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1649977179
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_449
timestamp 1649977179
transform 1 0 42412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_454
timestamp 1649977179
transform 1 0 42872 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_461
timestamp 1649977179
transform 1 0 43516 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_481
timestamp 1649977179
transform 1 0 45356 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_493
timestamp 1649977179
transform 1 0 46460 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_501
timestamp 1649977179
transform 1 0 47196 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1649977179
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_517
timestamp 1649977179
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_529
timestamp 1649977179
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_541
timestamp 1649977179
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1649977179
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1649977179
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_561
timestamp 1649977179
transform 1 0 52716 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_573
timestamp 1649977179
transform 1 0 53820 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_585
timestamp 1649977179
transform 1 0 54924 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_597
timestamp 1649977179
transform 1 0 56028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_609
timestamp 1649977179
transform 1 0 57132 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_615
timestamp 1649977179
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_617
timestamp 1649977179
transform 1 0 57868 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_629
timestamp 1649977179
transform 1 0 58972 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_641
timestamp 1649977179
transform 1 0 60076 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_653
timestamp 1649977179
transform 1 0 61180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_665
timestamp 1649977179
transform 1 0 62284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_671
timestamp 1649977179
transform 1 0 62836 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_673
timestamp 1649977179
transform 1 0 63020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_685
timestamp 1649977179
transform 1 0 64124 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_697
timestamp 1649977179
transform 1 0 65228 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_709
timestamp 1649977179
transform 1 0 66332 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_721
timestamp 1649977179
transform 1 0 67436 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_727
timestamp 1649977179
transform 1 0 67988 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_729
timestamp 1649977179
transform 1 0 68172 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_51
timestamp 1649977179
transform 1 0 5796 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_59
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1649977179
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_91
timestamp 1649977179
transform 1 0 9476 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_103
timestamp 1649977179
transform 1 0 10580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_111
timestamp 1649977179
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_120
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_126
timestamp 1649977179
transform 1 0 12696 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_159
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_176
timestamp 1649977179
transform 1 0 17296 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_186
timestamp 1649977179
transform 1 0 18216 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_203
timestamp 1649977179
transform 1 0 19780 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_211
timestamp 1649977179
transform 1 0 20516 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_216
timestamp 1649977179
transform 1 0 20976 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_230
timestamp 1649977179
transform 1 0 22264 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_257
timestamp 1649977179
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_268
timestamp 1649977179
transform 1 0 25760 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_288
timestamp 1649977179
transform 1 0 27600 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_295
timestamp 1649977179
transform 1 0 28244 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1649977179
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_325
timestamp 1649977179
transform 1 0 31004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_335
timestamp 1649977179
transform 1 0 31924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_342
timestamp 1649977179
transform 1 0 32568 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_350
timestamp 1649977179
transform 1 0 33304 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_360
timestamp 1649977179
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_381
timestamp 1649977179
transform 1 0 36156 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_402
timestamp 1649977179
transform 1 0 38088 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_415
timestamp 1649977179
transform 1 0 39284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1649977179
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_428
timestamp 1649977179
transform 1 0 40480 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_439
timestamp 1649977179
transform 1 0 41492 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_450
timestamp 1649977179
transform 1 0 42504 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_467
timestamp 1649977179
transform 1 0 44068 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1649977179
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_484
timestamp 1649977179
transform 1 0 45632 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_492
timestamp 1649977179
transform 1 0 46368 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_504
timestamp 1649977179
transform 1 0 47472 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_516
timestamp 1649977179
transform 1 0 48576 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_528
timestamp 1649977179
transform 1 0 49680 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_533
timestamp 1649977179
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_545
timestamp 1649977179
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_557
timestamp 1649977179
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_569
timestamp 1649977179
transform 1 0 53452 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1649977179
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1649977179
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_589
timestamp 1649977179
transform 1 0 55292 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_601
timestamp 1649977179
transform 1 0 56396 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_613
timestamp 1649977179
transform 1 0 57500 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_625
timestamp 1649977179
transform 1 0 58604 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_637
timestamp 1649977179
transform 1 0 59708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_643
timestamp 1649977179
transform 1 0 60260 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_645
timestamp 1649977179
transform 1 0 60444 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_657
timestamp 1649977179
transform 1 0 61548 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_669
timestamp 1649977179
transform 1 0 62652 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_681
timestamp 1649977179
transform 1 0 63756 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_693
timestamp 1649977179
transform 1 0 64860 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_699
timestamp 1649977179
transform 1 0 65412 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_701
timestamp 1649977179
transform 1 0 65596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_713
timestamp 1649977179
transform 1 0 66700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_725
timestamp 1649977179
transform 1 0 67804 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_34
timestamp 1649977179
transform 1 0 4232 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_47
timestamp 1649977179
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_59
timestamp 1649977179
transform 1 0 6532 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_72
timestamp 1649977179
transform 1 0 7728 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_78
timestamp 1649977179
transform 1 0 8280 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_90
timestamp 1649977179
transform 1 0 9384 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_98
timestamp 1649977179
transform 1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1649977179
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_120
timestamp 1649977179
transform 1 0 12144 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_127
timestamp 1649977179
transform 1 0 12788 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_133
timestamp 1649977179
transform 1 0 13340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_145
timestamp 1649977179
transform 1 0 14444 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_27_156
timestamp 1649977179
transform 1 0 15456 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_172
timestamp 1649977179
transform 1 0 16928 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_186
timestamp 1649977179
transform 1 0 18216 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_200
timestamp 1649977179
transform 1 0 19504 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_208
timestamp 1649977179
transform 1 0 20240 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_219
timestamp 1649977179
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_228
timestamp 1649977179
transform 1 0 22080 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_235
timestamp 1649977179
transform 1 0 22724 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_245
timestamp 1649977179
transform 1 0 23644 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_256
timestamp 1649977179
transform 1 0 24656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1649977179
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_287
timestamp 1649977179
transform 1 0 27508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1649977179
transform 1 0 28152 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_300
timestamp 1649977179
transform 1 0 28704 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_312
timestamp 1649977179
transform 1 0 29808 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_320
timestamp 1649977179
transform 1 0 30544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_325
timestamp 1649977179
transform 1 0 31004 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_333
timestamp 1649977179
transform 1 0 31740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_345
timestamp 1649977179
transform 1 0 32844 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_355
timestamp 1649977179
transform 1 0 33764 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_368
timestamp 1649977179
transform 1 0 34960 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_376
timestamp 1649977179
transform 1 0 35696 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_386
timestamp 1649977179
transform 1 0 36616 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_396
timestamp 1649977179
transform 1 0 37536 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_416
timestamp 1649977179
transform 1 0 39376 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_428
timestamp 1649977179
transform 1 0 40480 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_444
timestamp 1649977179
transform 1 0 41952 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_456
timestamp 1649977179
transform 1 0 43056 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_478
timestamp 1649977179
transform 1 0 45080 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_489
timestamp 1649977179
transform 1 0 46092 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_501
timestamp 1649977179
transform 1 0 47196 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1649977179
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_517
timestamp 1649977179
transform 1 0 48668 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_529
timestamp 1649977179
transform 1 0 49772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_541
timestamp 1649977179
transform 1 0 50876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_553
timestamp 1649977179
transform 1 0 51980 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_559
timestamp 1649977179
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_561
timestamp 1649977179
transform 1 0 52716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_573
timestamp 1649977179
transform 1 0 53820 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_585
timestamp 1649977179
transform 1 0 54924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_597
timestamp 1649977179
transform 1 0 56028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_609
timestamp 1649977179
transform 1 0 57132 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_615
timestamp 1649977179
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_617
timestamp 1649977179
transform 1 0 57868 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_629
timestamp 1649977179
transform 1 0 58972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_641
timestamp 1649977179
transform 1 0 60076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_653
timestamp 1649977179
transform 1 0 61180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_665
timestamp 1649977179
transform 1 0 62284 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_671
timestamp 1649977179
transform 1 0 62836 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_673
timestamp 1649977179
transform 1 0 63020 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_685
timestamp 1649977179
transform 1 0 64124 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_697
timestamp 1649977179
transform 1 0 65228 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_709
timestamp 1649977179
transform 1 0 66332 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_721
timestamp 1649977179
transform 1 0 67436 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_727
timestamp 1649977179
transform 1 0 67988 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_729
timestamp 1649977179
transform 1 0 68172 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_51
timestamp 1649977179
transform 1 0 5796 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_63
timestamp 1649977179
transform 1 0 6900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_75
timestamp 1649977179
transform 1 0 8004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_105
timestamp 1649977179
transform 1 0 10764 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_114
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_127
timestamp 1649977179
transform 1 0 12788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_135
timestamp 1649977179
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_143
timestamp 1649977179
transform 1 0 14260 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_167
timestamp 1649977179
transform 1 0 16468 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_182
timestamp 1649977179
transform 1 0 17848 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_188
timestamp 1649977179
transform 1 0 18400 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_205
timestamp 1649977179
transform 1 0 19964 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_211
timestamp 1649977179
transform 1 0 20516 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1649977179
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_239
timestamp 1649977179
transform 1 0 23092 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1649977179
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_257
timestamp 1649977179
transform 1 0 24748 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1649977179
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_286
timestamp 1649977179
transform 1 0 27416 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_298
timestamp 1649977179
transform 1 0 28520 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1649977179
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_331
timestamp 1649977179
transform 1 0 31556 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_344
timestamp 1649977179
transform 1 0 32752 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_350
timestamp 1649977179
transform 1 0 33304 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_353
timestamp 1649977179
transform 1 0 33580 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1649977179
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_381
timestamp 1649977179
transform 1 0 36156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_385
timestamp 1649977179
transform 1 0 36524 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_390
timestamp 1649977179
transform 1 0 36984 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_412
timestamp 1649977179
transform 1 0 39008 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_424
timestamp 1649977179
transform 1 0 40112 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_436
timestamp 1649977179
transform 1 0 41216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_28_446
timestamp 1649977179
transform 1 0 42136 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_454
timestamp 1649977179
transform 1 0 42872 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_459
timestamp 1649977179
transform 1 0 43332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1649977179
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1649977179
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1649977179
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1649977179
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1649977179
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_525
timestamp 1649977179
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_531
timestamp 1649977179
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_533
timestamp 1649977179
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_545
timestamp 1649977179
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_557
timestamp 1649977179
transform 1 0 52348 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_569
timestamp 1649977179
transform 1 0 53452 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_581
timestamp 1649977179
transform 1 0 54556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1649977179
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_592
timestamp 1649977179
transform 1 0 55568 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_598
timestamp 1649977179
transform 1 0 56120 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_610
timestamp 1649977179
transform 1 0 57224 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_622
timestamp 1649977179
transform 1 0 58328 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_634
timestamp 1649977179
transform 1 0 59432 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_642
timestamp 1649977179
transform 1 0 60168 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_645
timestamp 1649977179
transform 1 0 60444 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_657
timestamp 1649977179
transform 1 0 61548 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_669
timestamp 1649977179
transform 1 0 62652 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_681
timestamp 1649977179
transform 1 0 63756 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_693
timestamp 1649977179
transform 1 0 64860 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_699
timestamp 1649977179
transform 1 0 65412 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_701
timestamp 1649977179
transform 1 0 65596 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_713
timestamp 1649977179
transform 1 0 66700 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_725
timestamp 1649977179
transform 1 0 67804 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_65
timestamp 1649977179
transform 1 0 7084 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_72
timestamp 1649977179
transform 1 0 7728 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_129
timestamp 1649977179
transform 1 0 12972 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_139
timestamp 1649977179
transform 1 0 13892 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_145
timestamp 1649977179
transform 1 0 14444 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_153
timestamp 1649977179
transform 1 0 15180 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1649977179
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_189
timestamp 1649977179
transform 1 0 18492 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_199
timestamp 1649977179
transform 1 0 19412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_203
timestamp 1649977179
transform 1 0 19780 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_206
timestamp 1649977179
transform 1 0 20056 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_220
timestamp 1649977179
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_231
timestamp 1649977179
transform 1 0 22356 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_243
timestamp 1649977179
transform 1 0 23460 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_255
timestamp 1649977179
transform 1 0 24564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_265
timestamp 1649977179
transform 1 0 25484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_271
timestamp 1649977179
transform 1 0 26036 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_283
timestamp 1649977179
transform 1 0 27140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_295
timestamp 1649977179
transform 1 0 28244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_303
timestamp 1649977179
transform 1 0 28980 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_308
timestamp 1649977179
transform 1 0 29440 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_316
timestamp 1649977179
transform 1 0 30176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1649977179
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_346
timestamp 1649977179
transform 1 0 32936 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_352
timestamp 1649977179
transform 1 0 33488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_357
timestamp 1649977179
transform 1 0 33948 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_366
timestamp 1649977179
transform 1 0 34776 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_378
timestamp 1649977179
transform 1 0 35880 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_390
timestamp 1649977179
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_406
timestamp 1649977179
transform 1 0 38456 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_413
timestamp 1649977179
transform 1 0 39100 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_425
timestamp 1649977179
transform 1 0 40204 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_437
timestamp 1649977179
transform 1 0 41308 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_445
timestamp 1649977179
transform 1 0 42044 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1649977179
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_463
timestamp 1649977179
transform 1 0 43700 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_475
timestamp 1649977179
transform 1 0 44804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_487
timestamp 1649977179
transform 1 0 45908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_499
timestamp 1649977179
transform 1 0 47012 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1649977179
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1649977179
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_517
timestamp 1649977179
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_529
timestamp 1649977179
transform 1 0 49772 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_541
timestamp 1649977179
transform 1 0 50876 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_553
timestamp 1649977179
transform 1 0 51980 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_559
timestamp 1649977179
transform 1 0 52532 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_561
timestamp 1649977179
transform 1 0 52716 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_573
timestamp 1649977179
transform 1 0 53820 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_585
timestamp 1649977179
transform 1 0 54924 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_597
timestamp 1649977179
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_609
timestamp 1649977179
transform 1 0 57132 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_615
timestamp 1649977179
transform 1 0 57684 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_617
timestamp 1649977179
transform 1 0 57868 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_629
timestamp 1649977179
transform 1 0 58972 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_641
timestamp 1649977179
transform 1 0 60076 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_653
timestamp 1649977179
transform 1 0 61180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_665
timestamp 1649977179
transform 1 0 62284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_671
timestamp 1649977179
transform 1 0 62836 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_673
timestamp 1649977179
transform 1 0 63020 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_685
timestamp 1649977179
transform 1 0 64124 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_697
timestamp 1649977179
transform 1 0 65228 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_709
timestamp 1649977179
transform 1 0 66332 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_721
timestamp 1649977179
transform 1 0 67436 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_727
timestamp 1649977179
transform 1 0 67988 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_729
timestamp 1649977179
transform 1 0 68172 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_51
timestamp 1649977179
transform 1 0 5796 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_57
timestamp 1649977179
transform 1 0 6348 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_71
timestamp 1649977179
transform 1 0 7636 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_74
timestamp 1649977179
transform 1 0 7912 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_107
timestamp 1649977179
transform 1 0 10948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_113
timestamp 1649977179
transform 1 0 11500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_117
timestamp 1649977179
transform 1 0 11868 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_127
timestamp 1649977179
transform 1 0 12788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_171
timestamp 1649977179
transform 1 0 16836 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_175
timestamp 1649977179
transform 1 0 17204 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_184
timestamp 1649977179
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_204
timestamp 1649977179
transform 1 0 19872 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_210
timestamp 1649977179
transform 1 0 20424 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_214
timestamp 1649977179
transform 1 0 20792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_234
timestamp 1649977179
transform 1 0 22632 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_246
timestamp 1649977179
transform 1 0 23736 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_259
timestamp 1649977179
transform 1 0 24932 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_272
timestamp 1649977179
transform 1 0 26128 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_280
timestamp 1649977179
transform 1 0 26864 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_283
timestamp 1649977179
transform 1 0 27140 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_294
timestamp 1649977179
transform 1 0 28152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1649977179
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_311
timestamp 1649977179
transform 1 0 29716 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_323
timestamp 1649977179
transform 1 0 30820 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_329
timestamp 1649977179
transform 1 0 31372 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_346
timestamp 1649977179
transform 1 0 32936 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_359
timestamp 1649977179
transform 1 0 34132 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_397
timestamp 1649977179
transform 1 0 37628 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_416
timestamp 1649977179
transform 1 0 39376 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_421
timestamp 1649977179
transform 1 0 39836 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_427
timestamp 1649977179
transform 1 0 40388 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_439
timestamp 1649977179
transform 1 0 41492 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_451
timestamp 1649977179
transform 1 0 42596 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_463
timestamp 1649977179
transform 1 0 43700 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_467
timestamp 1649977179
transform 1 0 44068 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1649977179
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1649977179
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_480
timestamp 1649977179
transform 1 0 45264 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_492
timestamp 1649977179
transform 1 0 46368 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_504
timestamp 1649977179
transform 1 0 47472 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_516
timestamp 1649977179
transform 1 0 48576 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_528
timestamp 1649977179
transform 1 0 49680 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_533
timestamp 1649977179
transform 1 0 50140 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_545
timestamp 1649977179
transform 1 0 51244 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_557
timestamp 1649977179
transform 1 0 52348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_569
timestamp 1649977179
transform 1 0 53452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_581
timestamp 1649977179
transform 1 0 54556 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_587
timestamp 1649977179
transform 1 0 55108 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_589
timestamp 1649977179
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_601
timestamp 1649977179
transform 1 0 56396 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_613
timestamp 1649977179
transform 1 0 57500 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_625
timestamp 1649977179
transform 1 0 58604 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_637
timestamp 1649977179
transform 1 0 59708 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_643
timestamp 1649977179
transform 1 0 60260 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_645
timestamp 1649977179
transform 1 0 60444 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_657
timestamp 1649977179
transform 1 0 61548 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_669
timestamp 1649977179
transform 1 0 62652 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_681
timestamp 1649977179
transform 1 0 63756 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_693
timestamp 1649977179
transform 1 0 64860 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_699
timestamp 1649977179
transform 1 0 65412 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_701
timestamp 1649977179
transform 1 0 65596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_713
timestamp 1649977179
transform 1 0 66700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_729
timestamp 1649977179
transform 1 0 68172 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_31
timestamp 1649977179
transform 1 0 3956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_63
timestamp 1649977179
transform 1 0 6900 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_71
timestamp 1649977179
transform 1 0 7636 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_83
timestamp 1649977179
transform 1 0 8740 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1649977179
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1649977179
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_115
timestamp 1649977179
transform 1 0 11684 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_127
timestamp 1649977179
transform 1 0 12788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_139
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1649977179
transform 1 0 15548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1649977179
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_171
timestamp 1649977179
transform 1 0 16836 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_183
timestamp 1649977179
transform 1 0 17940 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_191
timestamp 1649977179
transform 1 0 18676 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_196
timestamp 1649977179
transform 1 0 19136 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_207
timestamp 1649977179
transform 1 0 20148 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1649977179
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_227
timestamp 1649977179
transform 1 0 21988 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_235
timestamp 1649977179
transform 1 0 22724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_269
timestamp 1649977179
transform 1 0 25852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_275
timestamp 1649977179
transform 1 0 26404 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1649977179
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_354
timestamp 1649977179
transform 1 0 33672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_362
timestamp 1649977179
transform 1 0 34408 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_367
timestamp 1649977179
transform 1 0 34868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_379
timestamp 1649977179
transform 1 0 35972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_424
timestamp 1649977179
transform 1 0 40112 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_433
timestamp 1649977179
transform 1 0 40940 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_445
timestamp 1649977179
transform 1 0 42044 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_449
timestamp 1649977179
transform 1 0 42412 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_457
timestamp 1649977179
transform 1 0 43148 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_479
timestamp 1649977179
transform 1 0 45172 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_491
timestamp 1649977179
transform 1 0 46276 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1649977179
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1649977179
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_517
timestamp 1649977179
transform 1 0 48668 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_529
timestamp 1649977179
transform 1 0 49772 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_541
timestamp 1649977179
transform 1 0 50876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_553
timestamp 1649977179
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_559
timestamp 1649977179
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_561
timestamp 1649977179
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_573
timestamp 1649977179
transform 1 0 53820 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_585
timestamp 1649977179
transform 1 0 54924 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_597
timestamp 1649977179
transform 1 0 56028 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_609
timestamp 1649977179
transform 1 0 57132 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_615
timestamp 1649977179
transform 1 0 57684 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_617
timestamp 1649977179
transform 1 0 57868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_629
timestamp 1649977179
transform 1 0 58972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_641
timestamp 1649977179
transform 1 0 60076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_653
timestamp 1649977179
transform 1 0 61180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_665
timestamp 1649977179
transform 1 0 62284 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_671
timestamp 1649977179
transform 1 0 62836 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_673
timestamp 1649977179
transform 1 0 63020 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_685
timestamp 1649977179
transform 1 0 64124 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_697
timestamp 1649977179
transform 1 0 65228 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_709
timestamp 1649977179
transform 1 0 66332 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_721
timestamp 1649977179
transform 1 0 67436 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_727
timestamp 1649977179
transform 1 0 67988 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_729
timestamp 1649977179
transform 1 0 68172 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_37
timestamp 1649977179
transform 1 0 4508 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_47
timestamp 1649977179
transform 1 0 5428 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_60
timestamp 1649977179
transform 1 0 6624 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_66
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_70
timestamp 1649977179
transform 1 0 7544 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_90
timestamp 1649977179
transform 1 0 9384 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1649977179
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_127
timestamp 1649977179
transform 1 0 12788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_143
timestamp 1649977179
transform 1 0 14260 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1649977179
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_170
timestamp 1649977179
transform 1 0 16744 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_176
timestamp 1649977179
transform 1 0 17296 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_182
timestamp 1649977179
transform 1 0 17848 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_185
timestamp 1649977179
transform 1 0 18124 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_207
timestamp 1649977179
transform 1 0 20148 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_214
timestamp 1649977179
transform 1 0 20792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_220
timestamp 1649977179
transform 1 0 21344 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_228
timestamp 1649977179
transform 1 0 22080 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_243
timestamp 1649977179
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_272
timestamp 1649977179
transform 1 0 26128 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_287
timestamp 1649977179
transform 1 0 27508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_299
timestamp 1649977179
transform 1 0 28612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_320
timestamp 1649977179
transform 1 0 30544 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_328
timestamp 1649977179
transform 1 0 31280 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_338
timestamp 1649977179
transform 1 0 32200 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1649977179
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_376
timestamp 1649977179
transform 1 0 35696 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_388
timestamp 1649977179
transform 1 0 36800 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_392
timestamp 1649977179
transform 1 0 37168 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_400
timestamp 1649977179
transform 1 0 37904 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_412
timestamp 1649977179
transform 1 0 39008 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1649977179
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_431
timestamp 1649977179
transform 1 0 40756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_435
timestamp 1649977179
transform 1 0 41124 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_441
timestamp 1649977179
transform 1 0 41676 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_465
timestamp 1649977179
transform 1 0 43884 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_473
timestamp 1649977179
transform 1 0 44620 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_483
timestamp 1649977179
transform 1 0 45540 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_495
timestamp 1649977179
transform 1 0 46644 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_507
timestamp 1649977179
transform 1 0 47748 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_519
timestamp 1649977179
transform 1 0 48852 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_531
timestamp 1649977179
transform 1 0 49956 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_533
timestamp 1649977179
transform 1 0 50140 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_545
timestamp 1649977179
transform 1 0 51244 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_557
timestamp 1649977179
transform 1 0 52348 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_569
timestamp 1649977179
transform 1 0 53452 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_581
timestamp 1649977179
transform 1 0 54556 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1649977179
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_589
timestamp 1649977179
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_601
timestamp 1649977179
transform 1 0 56396 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_613
timestamp 1649977179
transform 1 0 57500 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_625
timestamp 1649977179
transform 1 0 58604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_637
timestamp 1649977179
transform 1 0 59708 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_643
timestamp 1649977179
transform 1 0 60260 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_645
timestamp 1649977179
transform 1 0 60444 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_657
timestamp 1649977179
transform 1 0 61548 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_669
timestamp 1649977179
transform 1 0 62652 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_681
timestamp 1649977179
transform 1 0 63756 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_693
timestamp 1649977179
transform 1 0 64860 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_699
timestamp 1649977179
transform 1 0 65412 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_701
timestamp 1649977179
transform 1 0 65596 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_713
timestamp 1649977179
transform 1 0 66700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_725
timestamp 1649977179
transform 1 0 67804 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_49
timestamp 1649977179
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_60
timestamp 1649977179
transform 1 0 6624 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_66
timestamp 1649977179
transform 1 0 7176 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_74
timestamp 1649977179
transform 1 0 7912 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_82
timestamp 1649977179
transform 1 0 8648 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_91
timestamp 1649977179
transform 1 0 9476 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_101
timestamp 1649977179
transform 1 0 10396 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1649977179
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_115
timestamp 1649977179
transform 1 0 11684 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_121
timestamp 1649977179
transform 1 0 12236 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_133
timestamp 1649977179
transform 1 0 13340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_150
timestamp 1649977179
transform 1 0 14904 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1649977179
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_178
timestamp 1649977179
transform 1 0 17480 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1649977179
transform 1 0 17848 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_186
timestamp 1649977179
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1649977179
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_211
timestamp 1649977179
transform 1 0 20516 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_220
timestamp 1649977179
transform 1 0 21344 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_229
timestamp 1649977179
transform 1 0 22172 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_239
timestamp 1649977179
transform 1 0 23092 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_247
timestamp 1649977179
transform 1 0 23828 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_251
timestamp 1649977179
transform 1 0 24196 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_271
timestamp 1649977179
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_296
timestamp 1649977179
transform 1 0 28336 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_302
timestamp 1649977179
transform 1 0 28888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_306
timestamp 1649977179
transform 1 0 29256 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_315
timestamp 1649977179
transform 1 0 30084 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_327
timestamp 1649977179
transform 1 0 31188 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_346
timestamp 1649977179
transform 1 0 32936 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_354
timestamp 1649977179
transform 1 0 33672 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_358
timestamp 1649977179
transform 1 0 34040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_378
timestamp 1649977179
transform 1 0 35880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_398
timestamp 1649977179
transform 1 0 37720 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_413
timestamp 1649977179
transform 1 0 39100 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_421
timestamp 1649977179
transform 1 0 39836 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_430
timestamp 1649977179
transform 1 0 40664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_444
timestamp 1649977179
transform 1 0 41952 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_455
timestamp 1649977179
transform 1 0 42964 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_461
timestamp 1649977179
transform 1 0 43516 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_482
timestamp 1649977179
transform 1 0 45448 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_498
timestamp 1649977179
transform 1 0 46920 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1649977179
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_517
timestamp 1649977179
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_529
timestamp 1649977179
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_541
timestamp 1649977179
transform 1 0 50876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_553
timestamp 1649977179
transform 1 0 51980 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_559
timestamp 1649977179
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_561
timestamp 1649977179
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_573
timestamp 1649977179
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_585
timestamp 1649977179
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_597
timestamp 1649977179
transform 1 0 56028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_609
timestamp 1649977179
transform 1 0 57132 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1649977179
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_617
timestamp 1649977179
transform 1 0 57868 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_629
timestamp 1649977179
transform 1 0 58972 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_641
timestamp 1649977179
transform 1 0 60076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_653
timestamp 1649977179
transform 1 0 61180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_665
timestamp 1649977179
transform 1 0 62284 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_671
timestamp 1649977179
transform 1 0 62836 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_673
timestamp 1649977179
transform 1 0 63020 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_685
timestamp 1649977179
transform 1 0 64124 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_697
timestamp 1649977179
transform 1 0 65228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_709
timestamp 1649977179
transform 1 0 66332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_721
timestamp 1649977179
transform 1 0 67436 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_727
timestamp 1649977179
transform 1 0 67988 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_729
timestamp 1649977179
transform 1 0 68172 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_60
timestamp 1649977179
transform 1 0 6624 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_73
timestamp 1649977179
transform 1 0 7820 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_81
timestamp 1649977179
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_95
timestamp 1649977179
transform 1 0 9844 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_108
timestamp 1649977179
transform 1 0 11040 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_127
timestamp 1649977179
transform 1 0 12788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_161
timestamp 1649977179
transform 1 0 15916 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_167
timestamp 1649977179
transform 1 0 16468 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_184
timestamp 1649977179
transform 1 0 18032 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 1649977179
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_207
timestamp 1649977179
transform 1 0 20148 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_263
timestamp 1649977179
transform 1 0 25300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_271
timestamp 1649977179
transform 1 0 26036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_285
timestamp 1649977179
transform 1 0 27324 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_292
timestamp 1649977179
transform 1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1649977179
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_315
timestamp 1649977179
transform 1 0 30084 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_324
timestamp 1649977179
transform 1 0 30912 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_339
timestamp 1649977179
transform 1 0 32292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_354
timestamp 1649977179
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1649977179
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_367
timestamp 1649977179
transform 1 0 34868 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_397
timestamp 1649977179
transform 1 0 37628 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_408
timestamp 1649977179
transform 1 0 38640 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_427
timestamp 1649977179
transform 1 0 40388 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_431
timestamp 1649977179
transform 1 0 40756 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_434
timestamp 1649977179
transform 1 0 41032 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_440
timestamp 1649977179
transform 1 0 41584 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_444
timestamp 1649977179
transform 1 0 41952 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_453
timestamp 1649977179
transform 1 0 42780 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1649977179
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1649977179
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_480
timestamp 1649977179
transform 1 0 45264 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_487
timestamp 1649977179
transform 1 0 45908 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_499
timestamp 1649977179
transform 1 0 47012 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_511
timestamp 1649977179
transform 1 0 48116 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_523
timestamp 1649977179
transform 1 0 49220 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_531
timestamp 1649977179
transform 1 0 49956 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_533
timestamp 1649977179
transform 1 0 50140 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_545
timestamp 1649977179
transform 1 0 51244 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_557
timestamp 1649977179
transform 1 0 52348 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_569
timestamp 1649977179
transform 1 0 53452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_581
timestamp 1649977179
transform 1 0 54556 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1649977179
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_589
timestamp 1649977179
transform 1 0 55292 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_601
timestamp 1649977179
transform 1 0 56396 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_613
timestamp 1649977179
transform 1 0 57500 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_625
timestamp 1649977179
transform 1 0 58604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_637
timestamp 1649977179
transform 1 0 59708 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_643
timestamp 1649977179
transform 1 0 60260 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_645
timestamp 1649977179
transform 1 0 60444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_657
timestamp 1649977179
transform 1 0 61548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_669
timestamp 1649977179
transform 1 0 62652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_681
timestamp 1649977179
transform 1 0 63756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_693
timestamp 1649977179
transform 1 0 64860 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_699
timestamp 1649977179
transform 1 0 65412 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_701
timestamp 1649977179
transform 1 0 65596 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_713
timestamp 1649977179
transform 1 0 66700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_725
timestamp 1649977179
transform 1 0 67804 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1649977179
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_59
timestamp 1649977179
transform 1 0 6532 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_70
timestamp 1649977179
transform 1 0 7544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_80
timestamp 1649977179
transform 1 0 8464 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_84
timestamp 1649977179
transform 1 0 8832 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_90
timestamp 1649977179
transform 1 0 9384 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_96
timestamp 1649977179
transform 1 0 9936 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_100
timestamp 1649977179
transform 1 0 10304 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_104
timestamp 1649977179
transform 1 0 10672 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_108
timestamp 1649977179
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_129
timestamp 1649977179
transform 1 0 12972 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_146
timestamp 1649977179
transform 1 0 14536 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_153
timestamp 1649977179
transform 1 0 15180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_165
timestamp 1649977179
transform 1 0 16284 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_172
timestamp 1649977179
transform 1 0 16928 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_198
timestamp 1649977179
transform 1 0 19320 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_202
timestamp 1649977179
transform 1 0 19688 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1649977179
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_227
timestamp 1649977179
transform 1 0 21988 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_239
timestamp 1649977179
transform 1 0 23092 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_247
timestamp 1649977179
transform 1 0 23828 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1649977179
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_262
timestamp 1649977179
transform 1 0 25208 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1649977179
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_289
timestamp 1649977179
transform 1 0 27692 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_292
timestamp 1649977179
transform 1 0 27968 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_302
timestamp 1649977179
transform 1 0 28888 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_35_316
timestamp 1649977179
transform 1 0 30176 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_323
timestamp 1649977179
transform 1 0 30820 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_345
timestamp 1649977179
transform 1 0 32844 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_351
timestamp 1649977179
transform 1 0 33396 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_363
timestamp 1649977179
transform 1 0 34500 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_366
timestamp 1649977179
transform 1 0 34776 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_379
timestamp 1649977179
transform 1 0 35972 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_388
timestamp 1649977179
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_395
timestamp 1649977179
transform 1 0 37444 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_406
timestamp 1649977179
transform 1 0 38456 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_418
timestamp 1649977179
transform 1 0 39560 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_430
timestamp 1649977179
transform 1 0 40664 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_442
timestamp 1649977179
transform 1 0 41768 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1649977179
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_461
timestamp 1649977179
transform 1 0 43516 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_472
timestamp 1649977179
transform 1 0 44528 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_484
timestamp 1649977179
transform 1 0 45632 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_500
timestamp 1649977179
transform 1 0 47104 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_505
timestamp 1649977179
transform 1 0 47564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_517
timestamp 1649977179
transform 1 0 48668 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_529
timestamp 1649977179
transform 1 0 49772 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_541
timestamp 1649977179
transform 1 0 50876 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_553
timestamp 1649977179
transform 1 0 51980 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_559
timestamp 1649977179
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_561
timestamp 1649977179
transform 1 0 52716 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_573
timestamp 1649977179
transform 1 0 53820 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_585
timestamp 1649977179
transform 1 0 54924 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_597
timestamp 1649977179
transform 1 0 56028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_609
timestamp 1649977179
transform 1 0 57132 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_615
timestamp 1649977179
transform 1 0 57684 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_617
timestamp 1649977179
transform 1 0 57868 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_629
timestamp 1649977179
transform 1 0 58972 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_641
timestamp 1649977179
transform 1 0 60076 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_653
timestamp 1649977179
transform 1 0 61180 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_665
timestamp 1649977179
transform 1 0 62284 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_671
timestamp 1649977179
transform 1 0 62836 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_673
timestamp 1649977179
transform 1 0 63020 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_685
timestamp 1649977179
transform 1 0 64124 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_697
timestamp 1649977179
transform 1 0 65228 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_709
timestamp 1649977179
transform 1 0 66332 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_721
timestamp 1649977179
transform 1 0 67436 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_727
timestamp 1649977179
transform 1 0 67988 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_729
timestamp 1649977179
transform 1 0 68172 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_51
timestamp 1649977179
transform 1 0 5796 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_58
timestamp 1649977179
transform 1 0 6440 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_70
timestamp 1649977179
transform 1 0 7544 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1649977179
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_100
timestamp 1649977179
transform 1 0 10304 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_106
timestamp 1649977179
transform 1 0 10856 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_118
timestamp 1649977179
transform 1 0 11960 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_127
timestamp 1649977179
transform 1 0 12788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_143
timestamp 1649977179
transform 1 0 14260 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_155
timestamp 1649977179
transform 1 0 15364 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_158
timestamp 1649977179
transform 1 0 15640 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_171
timestamp 1649977179
transform 1 0 16836 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_179
timestamp 1649977179
transform 1 0 17572 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_186
timestamp 1649977179
transform 1 0 18216 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1649977179
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_205
timestamp 1649977179
transform 1 0 19964 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_216
timestamp 1649977179
transform 1 0 20976 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_223
timestamp 1649977179
transform 1 0 21620 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_231
timestamp 1649977179
transform 1 0 22356 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_238
timestamp 1649977179
transform 1 0 23000 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1649977179
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_257
timestamp 1649977179
transform 1 0 24748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_267
timestamp 1649977179
transform 1 0 25668 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_287
timestamp 1649977179
transform 1 0 27508 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_299
timestamp 1649977179
transform 1 0 28612 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_316
timestamp 1649977179
transform 1 0 30176 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_322
timestamp 1649977179
transform 1 0 30728 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_325
timestamp 1649977179
transform 1 0 31004 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_331
timestamp 1649977179
transform 1 0 31556 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_342
timestamp 1649977179
transform 1 0 32568 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_354
timestamp 1649977179
transform 1 0 33672 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1649977179
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_372
timestamp 1649977179
transform 1 0 35328 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_384
timestamp 1649977179
transform 1 0 36432 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_390
timestamp 1649977179
transform 1 0 36984 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_400
timestamp 1649977179
transform 1 0 37904 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_412
timestamp 1649977179
transform 1 0 39008 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_424
timestamp 1649977179
transform 1 0 40112 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_428
timestamp 1649977179
transform 1 0 40480 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_449
timestamp 1649977179
transform 1 0 42412 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_461
timestamp 1649977179
transform 1 0 43516 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_473
timestamp 1649977179
transform 1 0 44620 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1649977179
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1649977179
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_501
timestamp 1649977179
transform 1 0 47196 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_513
timestamp 1649977179
transform 1 0 48300 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_525
timestamp 1649977179
transform 1 0 49404 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_531
timestamp 1649977179
transform 1 0 49956 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_533
timestamp 1649977179
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_545
timestamp 1649977179
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_557
timestamp 1649977179
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_569
timestamp 1649977179
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1649977179
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1649977179
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_589
timestamp 1649977179
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_601
timestamp 1649977179
transform 1 0 56396 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_613
timestamp 1649977179
transform 1 0 57500 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_625
timestamp 1649977179
transform 1 0 58604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_637
timestamp 1649977179
transform 1 0 59708 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_643
timestamp 1649977179
transform 1 0 60260 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_645
timestamp 1649977179
transform 1 0 60444 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_657
timestamp 1649977179
transform 1 0 61548 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_669
timestamp 1649977179
transform 1 0 62652 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_681
timestamp 1649977179
transform 1 0 63756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_693
timestamp 1649977179
transform 1 0 64860 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_699
timestamp 1649977179
transform 1 0 65412 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_701
timestamp 1649977179
transform 1 0 65596 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_713
timestamp 1649977179
transform 1 0 66700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_725
timestamp 1649977179
transform 1 0 67804 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_40
timestamp 1649977179
transform 1 0 4784 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_49
timestamp 1649977179
transform 1 0 5612 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_60
timestamp 1649977179
transform 1 0 6624 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_72
timestamp 1649977179
transform 1 0 7728 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_84
timestamp 1649977179
transform 1 0 8832 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_96
timestamp 1649977179
transform 1 0 9936 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_102
timestamp 1649977179
transform 1 0 10488 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1649977179
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_119
timestamp 1649977179
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_131
timestamp 1649977179
transform 1 0 13156 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_141
timestamp 1649977179
transform 1 0 14076 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_152
timestamp 1649977179
transform 1 0 15088 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_160
timestamp 1649977179
transform 1 0 15824 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1649977179
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_176
timestamp 1649977179
transform 1 0 17296 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_184
timestamp 1649977179
transform 1 0 18032 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_191
timestamp 1649977179
transform 1 0 18676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_203
timestamp 1649977179
transform 1 0 19780 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_215
timestamp 1649977179
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_248
timestamp 1649977179
transform 1 0 23920 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_256
timestamp 1649977179
transform 1 0 24656 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_262
timestamp 1649977179
transform 1 0 25208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_266
timestamp 1649977179
transform 1 0 25576 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_269
timestamp 1649977179
transform 1 0 25852 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1649977179
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_290
timestamp 1649977179
transform 1 0 27784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_302
timestamp 1649977179
transform 1 0 28888 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_310
timestamp 1649977179
transform 1 0 29624 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_319
timestamp 1649977179
transform 1 0 30452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_325
timestamp 1649977179
transform 1 0 31004 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1649977179
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_343
timestamp 1649977179
transform 1 0 32660 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_347
timestamp 1649977179
transform 1 0 33028 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_354
timestamp 1649977179
transform 1 0 33672 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_366
timestamp 1649977179
transform 1 0 34776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_369
timestamp 1649977179
transform 1 0 35052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_381
timestamp 1649977179
transform 1 0 36156 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_389
timestamp 1649977179
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_416
timestamp 1649977179
transform 1 0 39376 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_424
timestamp 1649977179
transform 1 0 40112 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_437
timestamp 1649977179
transform 1 0 41308 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_445
timestamp 1649977179
transform 1 0 42044 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1649977179
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_461
timestamp 1649977179
transform 1 0 43516 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_485
timestamp 1649977179
transform 1 0 45724 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_492
timestamp 1649977179
transform 1 0 46368 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1649977179
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_517
timestamp 1649977179
transform 1 0 48668 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_529
timestamp 1649977179
transform 1 0 49772 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_541
timestamp 1649977179
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_553
timestamp 1649977179
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_559
timestamp 1649977179
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_561
timestamp 1649977179
transform 1 0 52716 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_573
timestamp 1649977179
transform 1 0 53820 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_585
timestamp 1649977179
transform 1 0 54924 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_597
timestamp 1649977179
transform 1 0 56028 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_609
timestamp 1649977179
transform 1 0 57132 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_615
timestamp 1649977179
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_617
timestamp 1649977179
transform 1 0 57868 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_629
timestamp 1649977179
transform 1 0 58972 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_641
timestamp 1649977179
transform 1 0 60076 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_653
timestamp 1649977179
transform 1 0 61180 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_665
timestamp 1649977179
transform 1 0 62284 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_671
timestamp 1649977179
transform 1 0 62836 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_673
timestamp 1649977179
transform 1 0 63020 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_685
timestamp 1649977179
transform 1 0 64124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_697
timestamp 1649977179
transform 1 0 65228 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_709
timestamp 1649977179
transform 1 0 66332 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_721
timestamp 1649977179
transform 1 0 67436 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_727
timestamp 1649977179
transform 1 0 67988 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_729
timestamp 1649977179
transform 1 0 68172 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_45
timestamp 1649977179
transform 1 0 5244 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_54
timestamp 1649977179
transform 1 0 6072 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_66
timestamp 1649977179
transform 1 0 7176 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1649977179
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_118
timestamp 1649977179
transform 1 0 11960 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1649977179
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_154
timestamp 1649977179
transform 1 0 15272 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_171
timestamp 1649977179
transform 1 0 16836 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_179
timestamp 1649977179
transform 1 0 17572 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_185
timestamp 1649977179
transform 1 0 18124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1649977179
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_202
timestamp 1649977179
transform 1 0 19688 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_213
timestamp 1649977179
transform 1 0 20700 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_242
timestamp 1649977179
transform 1 0 23368 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1649977179
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_253
timestamp 1649977179
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_265
timestamp 1649977179
transform 1 0 25484 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_273
timestamp 1649977179
transform 1 0 26220 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_278
timestamp 1649977179
transform 1 0 26680 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_284
timestamp 1649977179
transform 1 0 27232 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_288
timestamp 1649977179
transform 1 0 27600 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_292
timestamp 1649977179
transform 1 0 27968 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_300
timestamp 1649977179
transform 1 0 28704 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 1649977179
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_317
timestamp 1649977179
transform 1 0 30268 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_325
timestamp 1649977179
transform 1 0 31004 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_335
timestamp 1649977179
transform 1 0 31924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_343
timestamp 1649977179
transform 1 0 32660 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_351
timestamp 1649977179
transform 1 0 33396 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_370
timestamp 1649977179
transform 1 0 35144 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_382
timestamp 1649977179
transform 1 0 36248 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_396
timestamp 1649977179
transform 1 0 37536 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_411
timestamp 1649977179
transform 1 0 38916 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1649977179
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_427
timestamp 1649977179
transform 1 0 40388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_437
timestamp 1649977179
transform 1 0 41308 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_446
timestamp 1649977179
transform 1 0 42136 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_454
timestamp 1649977179
transform 1 0 42872 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_460
timestamp 1649977179
transform 1 0 43424 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_464
timestamp 1649977179
transform 1 0 43792 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_471
timestamp 1649977179
transform 1 0 44436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1649977179
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_489
timestamp 1649977179
transform 1 0 46092 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_499
timestamp 1649977179
transform 1 0 47012 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_506
timestamp 1649977179
transform 1 0 47656 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_518
timestamp 1649977179
transform 1 0 48760 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_530
timestamp 1649977179
transform 1 0 49864 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_533
timestamp 1649977179
transform 1 0 50140 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_545
timestamp 1649977179
transform 1 0 51244 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_557
timestamp 1649977179
transform 1 0 52348 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_569
timestamp 1649977179
transform 1 0 53452 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_581
timestamp 1649977179
transform 1 0 54556 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_587
timestamp 1649977179
transform 1 0 55108 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_589
timestamp 1649977179
transform 1 0 55292 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_601
timestamp 1649977179
transform 1 0 56396 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_613
timestamp 1649977179
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_625
timestamp 1649977179
transform 1 0 58604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_637
timestamp 1649977179
transform 1 0 59708 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_643
timestamp 1649977179
transform 1 0 60260 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_645
timestamp 1649977179
transform 1 0 60444 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_657
timestamp 1649977179
transform 1 0 61548 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_669
timestamp 1649977179
transform 1 0 62652 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_681
timestamp 1649977179
transform 1 0 63756 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_693
timestamp 1649977179
transform 1 0 64860 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_699
timestamp 1649977179
transform 1 0 65412 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_701
timestamp 1649977179
transform 1 0 65596 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_713
timestamp 1649977179
transform 1 0 66700 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_725
timestamp 1649977179
transform 1 0 67804 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_43
timestamp 1649977179
transform 1 0 5060 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1649977179
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_64
timestamp 1649977179
transform 1 0 6992 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_71
timestamp 1649977179
transform 1 0 7636 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_78
timestamp 1649977179
transform 1 0 8280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_85
timestamp 1649977179
transform 1 0 8924 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_97
timestamp 1649977179
transform 1 0 10028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_108
timestamp 1649977179
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_129
timestamp 1649977179
transform 1 0 12972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_136
timestamp 1649977179
transform 1 0 13616 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_142
timestamp 1649977179
transform 1 0 14168 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_154
timestamp 1649977179
transform 1 0 15272 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_164
timestamp 1649977179
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_171
timestamp 1649977179
transform 1 0 16836 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_180
timestamp 1649977179
transform 1 0 17664 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_188
timestamp 1649977179
transform 1 0 18400 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_192
timestamp 1649977179
transform 1 0 18768 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_204
timestamp 1649977179
transform 1 0 19872 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_208
timestamp 1649977179
transform 1 0 20240 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_216
timestamp 1649977179
transform 1 0 20976 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_230
timestamp 1649977179
transform 1 0 22264 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_238
timestamp 1649977179
transform 1 0 23000 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_246
timestamp 1649977179
transform 1 0 23736 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_256
timestamp 1649977179
transform 1 0 24656 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_264
timestamp 1649977179
transform 1 0 25392 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_272
timestamp 1649977179
transform 1 0 26128 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_288
timestamp 1649977179
transform 1 0 27600 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_292
timestamp 1649977179
transform 1 0 27968 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_299
timestamp 1649977179
transform 1 0 28612 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_306
timestamp 1649977179
transform 1 0 29256 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_310
timestamp 1649977179
transform 1 0 29624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_316
timestamp 1649977179
transform 1 0 30176 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_324
timestamp 1649977179
transform 1 0 30912 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_341
timestamp 1649977179
transform 1 0 32476 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_348
timestamp 1649977179
transform 1 0 33120 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_360
timestamp 1649977179
transform 1 0 34224 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_368
timestamp 1649977179
transform 1 0 34960 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_375
timestamp 1649977179
transform 1 0 35604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_386
timestamp 1649977179
transform 1 0 36616 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_400
timestamp 1649977179
transform 1 0 37904 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_416
timestamp 1649977179
transform 1 0 39376 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_432
timestamp 1649977179
transform 1 0 40848 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_439
timestamp 1649977179
transform 1 0 41492 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1649977179
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_452
timestamp 1649977179
transform 1 0 42688 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_461
timestamp 1649977179
transform 1 0 43516 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_485
timestamp 1649977179
transform 1 0 45724 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_495
timestamp 1649977179
transform 1 0 46644 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1649977179
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_518
timestamp 1649977179
transform 1 0 48760 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_530
timestamp 1649977179
transform 1 0 49864 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_542
timestamp 1649977179
transform 1 0 50968 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_554
timestamp 1649977179
transform 1 0 52072 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_561
timestamp 1649977179
transform 1 0 52716 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_573
timestamp 1649977179
transform 1 0 53820 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_585
timestamp 1649977179
transform 1 0 54924 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_597
timestamp 1649977179
transform 1 0 56028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_609
timestamp 1649977179
transform 1 0 57132 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1649977179
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_617
timestamp 1649977179
transform 1 0 57868 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_629
timestamp 1649977179
transform 1 0 58972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_641
timestamp 1649977179
transform 1 0 60076 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_653
timestamp 1649977179
transform 1 0 61180 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_665
timestamp 1649977179
transform 1 0 62284 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_671
timestamp 1649977179
transform 1 0 62836 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_673
timestamp 1649977179
transform 1 0 63020 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_685
timestamp 1649977179
transform 1 0 64124 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_697
timestamp 1649977179
transform 1 0 65228 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_709
timestamp 1649977179
transform 1 0 66332 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_721
timestamp 1649977179
transform 1 0 67436 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_727
timestamp 1649977179
transform 1 0 67988 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_729
timestamp 1649977179
transform 1 0 68172 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_35
timestamp 1649977179
transform 1 0 4324 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_43
timestamp 1649977179
transform 1 0 5060 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_51
timestamp 1649977179
transform 1 0 5796 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_60
timestamp 1649977179
transform 1 0 6624 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_66
timestamp 1649977179
transform 1 0 7176 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_76
timestamp 1649977179
transform 1 0 8096 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1649977179
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_96
timestamp 1649977179
transform 1 0 9936 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_108
timestamp 1649977179
transform 1 0 11040 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_112
timestamp 1649977179
transform 1 0 11408 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1649977179
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_151
timestamp 1649977179
transform 1 0 14996 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_157
timestamp 1649977179
transform 1 0 15548 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_161
timestamp 1649977179
transform 1 0 15916 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_167
timestamp 1649977179
transform 1 0 16468 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_173
timestamp 1649977179
transform 1 0 17020 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_181
timestamp 1649977179
transform 1 0 17756 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_185
timestamp 1649977179
transform 1 0 18124 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1649977179
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_210
timestamp 1649977179
transform 1 0 20424 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_237
timestamp 1649977179
transform 1 0 22908 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_263
timestamp 1649977179
transform 1 0 25300 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_274
timestamp 1649977179
transform 1 0 26312 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_286
timestamp 1649977179
transform 1 0 27416 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_290
timestamp 1649977179
transform 1 0 27784 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_293
timestamp 1649977179
transform 1 0 28060 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1649977179
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_312
timestamp 1649977179
transform 1 0 29808 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_318
timestamp 1649977179
transform 1 0 30360 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_330
timestamp 1649977179
transform 1 0 31464 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_342
timestamp 1649977179
transform 1 0 32568 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1649977179
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_368
timestamp 1649977179
transform 1 0 34960 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_396
timestamp 1649977179
transform 1 0 37536 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_408
timestamp 1649977179
transform 1 0 38640 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_421
timestamp 1649977179
transform 1 0 39836 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_427
timestamp 1649977179
transform 1 0 40388 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_448
timestamp 1649977179
transform 1 0 42320 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_465
timestamp 1649977179
transform 1 0 43884 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_472
timestamp 1649977179
transform 1 0 44528 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_485
timestamp 1649977179
transform 1 0 45724 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_494
timestamp 1649977179
transform 1 0 46552 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_501
timestamp 1649977179
transform 1 0 47196 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_513
timestamp 1649977179
transform 1 0 48300 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_525
timestamp 1649977179
transform 1 0 49404 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_531
timestamp 1649977179
transform 1 0 49956 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_533
timestamp 1649977179
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_545
timestamp 1649977179
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_557
timestamp 1649977179
transform 1 0 52348 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_569
timestamp 1649977179
transform 1 0 53452 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_581
timestamp 1649977179
transform 1 0 54556 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_587
timestamp 1649977179
transform 1 0 55108 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_589
timestamp 1649977179
transform 1 0 55292 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_601
timestamp 1649977179
transform 1 0 56396 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_613
timestamp 1649977179
transform 1 0 57500 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_625
timestamp 1649977179
transform 1 0 58604 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_637
timestamp 1649977179
transform 1 0 59708 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_643
timestamp 1649977179
transform 1 0 60260 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_645
timestamp 1649977179
transform 1 0 60444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_657
timestamp 1649977179
transform 1 0 61548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_669
timestamp 1649977179
transform 1 0 62652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_681
timestamp 1649977179
transform 1 0 63756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_693
timestamp 1649977179
transform 1 0 64860 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_699
timestamp 1649977179
transform 1 0 65412 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_701
timestamp 1649977179
transform 1 0 65596 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_713
timestamp 1649977179
transform 1 0 66700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_725
timestamp 1649977179
transform 1 0 67804 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_35
timestamp 1649977179
transform 1 0 4324 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_44
timestamp 1649977179
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_76
timestamp 1649977179
transform 1 0 8096 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_82
timestamp 1649977179
transform 1 0 8648 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_94
timestamp 1649977179
transform 1 0 9752 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_107
timestamp 1649977179
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_126
timestamp 1649977179
transform 1 0 12696 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_134
timestamp 1649977179
transform 1 0 13432 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_138
timestamp 1649977179
transform 1 0 13800 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_155
timestamp 1649977179
transform 1 0 15364 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1649977179
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_178
timestamp 1649977179
transform 1 0 17480 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_202
timestamp 1649977179
transform 1 0 19688 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_212
timestamp 1649977179
transform 1 0 20608 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_228
timestamp 1649977179
transform 1 0 22080 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_234
timestamp 1649977179
transform 1 0 22632 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_246
timestamp 1649977179
transform 1 0 23736 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_258
timestamp 1649977179
transform 1 0 24840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_266
timestamp 1649977179
transform 1 0 25576 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1649977179
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_289
timestamp 1649977179
transform 1 0 27692 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_300
timestamp 1649977179
transform 1 0 28704 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_307
timestamp 1649977179
transform 1 0 29348 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_313
timestamp 1649977179
transform 1 0 29900 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_325
timestamp 1649977179
transform 1 0 31004 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_333
timestamp 1649977179
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_343
timestamp 1649977179
transform 1 0 32660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_355
timestamp 1649977179
transform 1 0 33764 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_363
timestamp 1649977179
transform 1 0 34500 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_366
timestamp 1649977179
transform 1 0 34776 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_379
timestamp 1649977179
transform 1 0 35972 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_386
timestamp 1649977179
transform 1 0 36616 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1649977179
transform 1 0 38180 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_414
timestamp 1649977179
transform 1 0 39192 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_422
timestamp 1649977179
transform 1 0 39928 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_432
timestamp 1649977179
transform 1 0 40848 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_444
timestamp 1649977179
transform 1 0 41952 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1649977179
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_461
timestamp 1649977179
transform 1 0 43516 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_477
timestamp 1649977179
transform 1 0 44988 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_484
timestamp 1649977179
transform 1 0 45632 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_496
timestamp 1649977179
transform 1 0 46736 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_505
timestamp 1649977179
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_517
timestamp 1649977179
transform 1 0 48668 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_529
timestamp 1649977179
transform 1 0 49772 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_541
timestamp 1649977179
transform 1 0 50876 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_553
timestamp 1649977179
transform 1 0 51980 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_559
timestamp 1649977179
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_561
timestamp 1649977179
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_573
timestamp 1649977179
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_585
timestamp 1649977179
transform 1 0 54924 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_597
timestamp 1649977179
transform 1 0 56028 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_609
timestamp 1649977179
transform 1 0 57132 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_615
timestamp 1649977179
transform 1 0 57684 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_617
timestamp 1649977179
transform 1 0 57868 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_629
timestamp 1649977179
transform 1 0 58972 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_641
timestamp 1649977179
transform 1 0 60076 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_653
timestamp 1649977179
transform 1 0 61180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_665
timestamp 1649977179
transform 1 0 62284 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_671
timestamp 1649977179
transform 1 0 62836 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_673
timestamp 1649977179
transform 1 0 63020 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_685
timestamp 1649977179
transform 1 0 64124 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_697
timestamp 1649977179
transform 1 0 65228 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_709
timestamp 1649977179
transform 1 0 66332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_721
timestamp 1649977179
transform 1 0 67436 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_727
timestamp 1649977179
transform 1 0 67988 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_729
timestamp 1649977179
transform 1 0 68172 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_66
timestamp 1649977179
transform 1 0 7176 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_74
timestamp 1649977179
transform 1 0 7912 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1649977179
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_96
timestamp 1649977179
transform 1 0 9936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_108
timestamp 1649977179
transform 1 0 11040 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_111
timestamp 1649977179
transform 1 0 11316 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_117
timestamp 1649977179
transform 1 0 11868 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_125
timestamp 1649977179
transform 1 0 12604 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_128
timestamp 1649977179
transform 1 0 12880 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1649977179
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_147
timestamp 1649977179
transform 1 0 14628 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_160
timestamp 1649977179
transform 1 0 15824 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_170
timestamp 1649977179
transform 1 0 16744 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_178
timestamp 1649977179
transform 1 0 17480 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_200
timestamp 1649977179
transform 1 0 19504 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_212
timestamp 1649977179
transform 1 0 20608 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_224
timestamp 1649977179
transform 1 0 21712 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_232
timestamp 1649977179
transform 1 0 22448 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_237
timestamp 1649977179
transform 1 0 22908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_244
timestamp 1649977179
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_260
timestamp 1649977179
transform 1 0 25024 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_270
timestamp 1649977179
transform 1 0 25944 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_42_284
timestamp 1649977179
transform 1 0 27232 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_296
timestamp 1649977179
transform 1 0 28336 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_315
timestamp 1649977179
transform 1 0 30084 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_323
timestamp 1649977179
transform 1 0 30820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_329
timestamp 1649977179
transform 1 0 31372 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_342
timestamp 1649977179
transform 1 0 32568 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_352
timestamp 1649977179
transform 1 0 33488 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_391
timestamp 1649977179
transform 1 0 37076 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_413
timestamp 1649977179
transform 1 0 39100 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1649977179
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_421
timestamp 1649977179
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_433
timestamp 1649977179
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_445
timestamp 1649977179
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_457
timestamp 1649977179
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1649977179
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1649977179
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_477
timestamp 1649977179
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_489
timestamp 1649977179
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_501
timestamp 1649977179
transform 1 0 47196 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_513
timestamp 1649977179
transform 1 0 48300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_525
timestamp 1649977179
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_531
timestamp 1649977179
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_533
timestamp 1649977179
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_545
timestamp 1649977179
transform 1 0 51244 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_557
timestamp 1649977179
transform 1 0 52348 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_569
timestamp 1649977179
transform 1 0 53452 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_581
timestamp 1649977179
transform 1 0 54556 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_587
timestamp 1649977179
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_589
timestamp 1649977179
transform 1 0 55292 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_601
timestamp 1649977179
transform 1 0 56396 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_613
timestamp 1649977179
transform 1 0 57500 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_625
timestamp 1649977179
transform 1 0 58604 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_637
timestamp 1649977179
transform 1 0 59708 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_643
timestamp 1649977179
transform 1 0 60260 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_645
timestamp 1649977179
transform 1 0 60444 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_649
timestamp 1649977179
transform 1 0 60812 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_655
timestamp 1649977179
transform 1 0 61364 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_667
timestamp 1649977179
transform 1 0 62468 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_679
timestamp 1649977179
transform 1 0 63572 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_691
timestamp 1649977179
transform 1 0 64676 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_699
timestamp 1649977179
transform 1 0 65412 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_701
timestamp 1649977179
transform 1 0 65596 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_713
timestamp 1649977179
transform 1 0 66700 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_725
timestamp 1649977179
transform 1 0 67804 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_42
timestamp 1649977179
transform 1 0 4968 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_48
timestamp 1649977179
transform 1 0 5520 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_65
timestamp 1649977179
transform 1 0 7084 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_68
timestamp 1649977179
transform 1 0 7360 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_80
timestamp 1649977179
transform 1 0 8464 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_104
timestamp 1649977179
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_121
timestamp 1649977179
transform 1 0 12236 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_134
timestamp 1649977179
transform 1 0 13432 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_142
timestamp 1649977179
transform 1 0 14168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_156
timestamp 1649977179
transform 1 0 15456 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_160
timestamp 1649977179
transform 1 0 15824 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1649977179
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_196
timestamp 1649977179
transform 1 0 19136 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_204
timestamp 1649977179
transform 1 0 19872 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_210
timestamp 1649977179
transform 1 0 20424 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_222
timestamp 1649977179
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_228
timestamp 1649977179
transform 1 0 22080 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_234
timestamp 1649977179
transform 1 0 22632 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_244
timestamp 1649977179
transform 1 0 23552 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_250
timestamp 1649977179
transform 1 0 24104 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_259
timestamp 1649977179
transform 1 0 24932 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_270
timestamp 1649977179
transform 1 0 25944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1649977179
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_321
timestamp 1649977179
transform 1 0 30636 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_332
timestamp 1649977179
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_353
timestamp 1649977179
transform 1 0 33580 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_374
timestamp 1649977179
transform 1 0 35512 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_382
timestamp 1649977179
transform 1 0 36248 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_401
timestamp 1649977179
transform 1 0 37996 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_411
timestamp 1649977179
transform 1 0 38916 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_418
timestamp 1649977179
transform 1 0 39560 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_424
timestamp 1649977179
transform 1 0 40112 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_430
timestamp 1649977179
transform 1 0 40664 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_442
timestamp 1649977179
transform 1 0 41768 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1649977179
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1649977179
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1649977179
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_485
timestamp 1649977179
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1649977179
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1649977179
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1649977179
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_517
timestamp 1649977179
transform 1 0 48668 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_529
timestamp 1649977179
transform 1 0 49772 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_541
timestamp 1649977179
transform 1 0 50876 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_553
timestamp 1649977179
transform 1 0 51980 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_559
timestamp 1649977179
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_561
timestamp 1649977179
transform 1 0 52716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_573
timestamp 1649977179
transform 1 0 53820 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_585
timestamp 1649977179
transform 1 0 54924 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_597
timestamp 1649977179
transform 1 0 56028 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_609
timestamp 1649977179
transform 1 0 57132 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_615
timestamp 1649977179
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_617
timestamp 1649977179
transform 1 0 57868 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_629
timestamp 1649977179
transform 1 0 58972 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_641
timestamp 1649977179
transform 1 0 60076 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_653
timestamp 1649977179
transform 1 0 61180 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_665
timestamp 1649977179
transform 1 0 62284 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_671
timestamp 1649977179
transform 1 0 62836 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_673
timestamp 1649977179
transform 1 0 63020 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_685
timestamp 1649977179
transform 1 0 64124 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_697
timestamp 1649977179
transform 1 0 65228 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_709
timestamp 1649977179
transform 1 0 66332 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_721
timestamp 1649977179
transform 1 0 67436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_727
timestamp 1649977179
transform 1 0 67988 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_729
timestamp 1649977179
transform 1 0 68172 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_37
timestamp 1649977179
transform 1 0 4508 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_49
timestamp 1649977179
transform 1 0 5612 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_56
timestamp 1649977179
transform 1 0 6256 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_69
timestamp 1649977179
transform 1 0 7452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1649977179
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_92
timestamp 1649977179
transform 1 0 9568 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_98
timestamp 1649977179
transform 1 0 10120 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_104
timestamp 1649977179
transform 1 0 10672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_110
timestamp 1649977179
transform 1 0 11224 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_116
timestamp 1649977179
transform 1 0 11776 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_122
timestamp 1649977179
transform 1 0 12328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_129
timestamp 1649977179
transform 1 0 12972 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_137
timestamp 1649977179
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_149
timestamp 1649977179
transform 1 0 14812 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_178
timestamp 1649977179
transform 1 0 17480 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_184
timestamp 1649977179
transform 1 0 18032 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_207
timestamp 1649977179
transform 1 0 20148 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_217
timestamp 1649977179
transform 1 0 21068 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_229
timestamp 1649977179
transform 1 0 22172 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_241
timestamp 1649977179
transform 1 0 23276 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1649977179
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_263
timestamp 1649977179
transform 1 0 25300 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_269
timestamp 1649977179
transform 1 0 25852 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_281
timestamp 1649977179
transform 1 0 26956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_293
timestamp 1649977179
transform 1 0 28060 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1649977179
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_316
timestamp 1649977179
transform 1 0 30176 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_324
timestamp 1649977179
transform 1 0 30912 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_344
timestamp 1649977179
transform 1 0 32752 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1649977179
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_381
timestamp 1649977179
transform 1 0 36156 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_395
timestamp 1649977179
transform 1 0 37444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_399
timestamp 1649977179
transform 1 0 37812 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_404
timestamp 1649977179
transform 1 0 38272 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_416
timestamp 1649977179
transform 1 0 39376 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_427
timestamp 1649977179
transform 1 0 40388 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_436
timestamp 1649977179
transform 1 0 41216 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_456
timestamp 1649977179
transform 1 0 43056 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_468
timestamp 1649977179
transform 1 0 44160 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_480
timestamp 1649977179
transform 1 0 45264 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_492
timestamp 1649977179
transform 1 0 46368 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_504
timestamp 1649977179
transform 1 0 47472 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_516
timestamp 1649977179
transform 1 0 48576 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_528
timestamp 1649977179
transform 1 0 49680 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_533
timestamp 1649977179
transform 1 0 50140 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_545
timestamp 1649977179
transform 1 0 51244 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_557
timestamp 1649977179
transform 1 0 52348 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_569
timestamp 1649977179
transform 1 0 53452 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_581
timestamp 1649977179
transform 1 0 54556 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_587
timestamp 1649977179
transform 1 0 55108 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_589
timestamp 1649977179
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_601
timestamp 1649977179
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_613
timestamp 1649977179
transform 1 0 57500 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_625
timestamp 1649977179
transform 1 0 58604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_637
timestamp 1649977179
transform 1 0 59708 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_643
timestamp 1649977179
transform 1 0 60260 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_645
timestamp 1649977179
transform 1 0 60444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_657
timestamp 1649977179
transform 1 0 61548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_669
timestamp 1649977179
transform 1 0 62652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_681
timestamp 1649977179
transform 1 0 63756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_693
timestamp 1649977179
transform 1 0 64860 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_699
timestamp 1649977179
transform 1 0 65412 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_701
timestamp 1649977179
transform 1 0 65596 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_713
timestamp 1649977179
transform 1 0 66700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_729
timestamp 1649977179
transform 1 0 68172 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_35
timestamp 1649977179
transform 1 0 4324 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1649977179
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_73
timestamp 1649977179
transform 1 0 7820 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_77
timestamp 1649977179
transform 1 0 8188 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_84
timestamp 1649977179
transform 1 0 8832 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_95
timestamp 1649977179
transform 1 0 9844 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_108
timestamp 1649977179
transform 1 0 11040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_117
timestamp 1649977179
transform 1 0 11868 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_126
timestamp 1649977179
transform 1 0 12696 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_145
timestamp 1649977179
transform 1 0 14444 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_151
timestamp 1649977179
transform 1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_155
timestamp 1649977179
transform 1 0 15364 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_158
timestamp 1649977179
transform 1 0 15640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1649977179
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_173
timestamp 1649977179
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_177
timestamp 1649977179
transform 1 0 17388 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_183
timestamp 1649977179
transform 1 0 17940 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_200
timestamp 1649977179
transform 1 0 19504 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_213
timestamp 1649977179
transform 1 0 20700 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1649977179
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_233
timestamp 1649977179
transform 1 0 22540 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_241
timestamp 1649977179
transform 1 0 23276 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_254
timestamp 1649977179
transform 1 0 24472 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_265
timestamp 1649977179
transform 1 0 25484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_271
timestamp 1649977179
transform 1 0 26036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_289
timestamp 1649977179
transform 1 0 27692 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_301
timestamp 1649977179
transform 1 0 28796 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_313
timestamp 1649977179
transform 1 0 29900 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_323
timestamp 1649977179
transform 1 0 30820 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1649977179
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_340
timestamp 1649977179
transform 1 0 32384 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_352
timestamp 1649977179
transform 1 0 33488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_360
timestamp 1649977179
transform 1 0 34224 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_366
timestamp 1649977179
transform 1 0 34776 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_372
timestamp 1649977179
transform 1 0 35328 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_383
timestamp 1649977179
transform 1 0 36340 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_414
timestamp 1649977179
transform 1 0 39192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_426
timestamp 1649977179
transform 1 0 40296 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_436
timestamp 1649977179
transform 1 0 41216 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1649977179
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_461
timestamp 1649977179
transform 1 0 43516 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_482
timestamp 1649977179
transform 1 0 45448 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_489
timestamp 1649977179
transform 1 0 46092 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_501
timestamp 1649977179
transform 1 0 47196 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_505
timestamp 1649977179
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_517
timestamp 1649977179
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_529
timestamp 1649977179
transform 1 0 49772 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_541
timestamp 1649977179
transform 1 0 50876 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_553
timestamp 1649977179
transform 1 0 51980 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_559
timestamp 1649977179
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_561
timestamp 1649977179
transform 1 0 52716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_573
timestamp 1649977179
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_585
timestamp 1649977179
transform 1 0 54924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_597
timestamp 1649977179
transform 1 0 56028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_609
timestamp 1649977179
transform 1 0 57132 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_615
timestamp 1649977179
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_617
timestamp 1649977179
transform 1 0 57868 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_629
timestamp 1649977179
transform 1 0 58972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_641
timestamp 1649977179
transform 1 0 60076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_653
timestamp 1649977179
transform 1 0 61180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_665
timestamp 1649977179
transform 1 0 62284 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_671
timestamp 1649977179
transform 1 0 62836 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_673
timestamp 1649977179
transform 1 0 63020 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_685
timestamp 1649977179
transform 1 0 64124 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_697
timestamp 1649977179
transform 1 0 65228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_709
timestamp 1649977179
transform 1 0 66332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_721
timestamp 1649977179
transform 1 0 67436 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_727
timestamp 1649977179
transform 1 0 67988 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_729
timestamp 1649977179
transform 1 0 68172 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_35
timestamp 1649977179
transform 1 0 4324 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_39
timestamp 1649977179
transform 1 0 4692 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_59
timestamp 1649977179
transform 1 0 6532 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_66
timestamp 1649977179
transform 1 0 7176 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_78
timestamp 1649977179
transform 1 0 8280 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_89
timestamp 1649977179
transform 1 0 9292 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_100
timestamp 1649977179
transform 1 0 10304 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_106
timestamp 1649977179
transform 1 0 10856 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_116
timestamp 1649977179
transform 1 0 11776 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_122
timestamp 1649977179
transform 1 0 12328 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_126
timestamp 1649977179
transform 1 0 12696 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_129
timestamp 1649977179
transform 1 0 12972 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_137
timestamp 1649977179
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_152
timestamp 1649977179
transform 1 0 15088 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_158
timestamp 1649977179
transform 1 0 15640 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_170
timestamp 1649977179
transform 1 0 16744 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_174
timestamp 1649977179
transform 1 0 17112 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 1649977179
transform 1 0 18676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_206
timestamp 1649977179
transform 1 0 20056 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_216
timestamp 1649977179
transform 1 0 20976 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_220
timestamp 1649977179
transform 1 0 21344 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_228
timestamp 1649977179
transform 1 0 22080 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_235
timestamp 1649977179
transform 1 0 22724 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_243
timestamp 1649977179
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_261
timestamp 1649977179
transform 1 0 25116 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_269
timestamp 1649977179
transform 1 0 25852 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_286
timestamp 1649977179
transform 1 0 27416 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_290
timestamp 1649977179
transform 1 0 27784 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_297
timestamp 1649977179
transform 1 0 28428 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_304
timestamp 1649977179
transform 1 0 29072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_316
timestamp 1649977179
transform 1 0 30176 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_324
timestamp 1649977179
transform 1 0 30912 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_379
timestamp 1649977179
transform 1 0 35972 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_385
timestamp 1649977179
transform 1 0 36524 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_395
timestamp 1649977179
transform 1 0 37444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_409
timestamp 1649977179
transform 1 0 38732 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_416
timestamp 1649977179
transform 1 0 39376 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_427
timestamp 1649977179
transform 1 0 40388 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_433
timestamp 1649977179
transform 1 0 40940 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_443
timestamp 1649977179
transform 1 0 41860 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_450
timestamp 1649977179
transform 1 0 42504 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_458
timestamp 1649977179
transform 1 0 43240 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_472
timestamp 1649977179
transform 1 0 44528 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_483
timestamp 1649977179
transform 1 0 45540 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_495
timestamp 1649977179
transform 1 0 46644 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_507
timestamp 1649977179
transform 1 0 47748 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_519
timestamp 1649977179
transform 1 0 48852 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1649977179
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_533
timestamp 1649977179
transform 1 0 50140 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_545
timestamp 1649977179
transform 1 0 51244 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_557
timestamp 1649977179
transform 1 0 52348 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_569
timestamp 1649977179
transform 1 0 53452 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_581
timestamp 1649977179
transform 1 0 54556 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_587
timestamp 1649977179
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_589
timestamp 1649977179
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_601
timestamp 1649977179
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_613
timestamp 1649977179
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_625
timestamp 1649977179
transform 1 0 58604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_637
timestamp 1649977179
transform 1 0 59708 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_643
timestamp 1649977179
transform 1 0 60260 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_645
timestamp 1649977179
transform 1 0 60444 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_657
timestamp 1649977179
transform 1 0 61548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_669
timestamp 1649977179
transform 1 0 62652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_681
timestamp 1649977179
transform 1 0 63756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_693
timestamp 1649977179
transform 1 0 64860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_699
timestamp 1649977179
transform 1 0 65412 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_701
timestamp 1649977179
transform 1 0 65596 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_713
timestamp 1649977179
transform 1 0 66700 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_725
timestamp 1649977179
transform 1 0 67804 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_64
timestamp 1649977179
transform 1 0 6992 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_70
timestamp 1649977179
transform 1 0 7544 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_82
timestamp 1649977179
transform 1 0 8648 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_86
timestamp 1649977179
transform 1 0 9016 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_98
timestamp 1649977179
transform 1 0 10120 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1649977179
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_120
timestamp 1649977179
transform 1 0 12144 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_127
timestamp 1649977179
transform 1 0 12788 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_131
timestamp 1649977179
transform 1 0 13156 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_134
timestamp 1649977179
transform 1 0 13432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1649977179
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_173
timestamp 1649977179
transform 1 0 17020 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_176
timestamp 1649977179
transform 1 0 17296 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_182
timestamp 1649977179
transform 1 0 17848 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_188
timestamp 1649977179
transform 1 0 18400 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_194
timestamp 1649977179
transform 1 0 18952 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_202
timestamp 1649977179
transform 1 0 19688 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_206
timestamp 1649977179
transform 1 0 20056 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_209
timestamp 1649977179
transform 1 0 20332 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1649977179
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_243
timestamp 1649977179
transform 1 0 23460 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_251
timestamp 1649977179
transform 1 0 24196 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_262
timestamp 1649977179
transform 1 0 25208 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_270
timestamp 1649977179
transform 1 0 25944 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1649977179
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_290
timestamp 1649977179
transform 1 0 27784 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_301
timestamp 1649977179
transform 1 0 28796 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_309
timestamp 1649977179
transform 1 0 29532 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_319
timestamp 1649977179
transform 1 0 30452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1649977179
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_344
timestamp 1649977179
transform 1 0 32752 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_354
timestamp 1649977179
transform 1 0 33672 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_366
timestamp 1649977179
transform 1 0 34776 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_47_372
timestamp 1649977179
transform 1 0 35328 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_378
timestamp 1649977179
transform 1 0 35880 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1649977179
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_395
timestamp 1649977179
transform 1 0 37444 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_409
timestamp 1649977179
transform 1 0 38732 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_421
timestamp 1649977179
transform 1 0 39836 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_429
timestamp 1649977179
transform 1 0 40572 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_434
timestamp 1649977179
transform 1 0 41032 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_446
timestamp 1649977179
transform 1 0 42136 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1649977179
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_461
timestamp 1649977179
transform 1 0 43516 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_483
timestamp 1649977179
transform 1 0 45540 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_492
timestamp 1649977179
transform 1 0 46368 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_505
timestamp 1649977179
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_517
timestamp 1649977179
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_529
timestamp 1649977179
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_541
timestamp 1649977179
transform 1 0 50876 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_553
timestamp 1649977179
transform 1 0 51980 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1649977179
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_561
timestamp 1649977179
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_573
timestamp 1649977179
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_585
timestamp 1649977179
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_597
timestamp 1649977179
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_609
timestamp 1649977179
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_615
timestamp 1649977179
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_617
timestamp 1649977179
transform 1 0 57868 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_629
timestamp 1649977179
transform 1 0 58972 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_641
timestamp 1649977179
transform 1 0 60076 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_653
timestamp 1649977179
transform 1 0 61180 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_665
timestamp 1649977179
transform 1 0 62284 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_671
timestamp 1649977179
transform 1 0 62836 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_673
timestamp 1649977179
transform 1 0 63020 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_685
timestamp 1649977179
transform 1 0 64124 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_697
timestamp 1649977179
transform 1 0 65228 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_709
timestamp 1649977179
transform 1 0 66332 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_721
timestamp 1649977179
transform 1 0 67436 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_727
timestamp 1649977179
transform 1 0 67988 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_729
timestamp 1649977179
transform 1 0 68172 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_93
timestamp 1649977179
transform 1 0 9660 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_99
timestamp 1649977179
transform 1 0 10212 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_105
timestamp 1649977179
transform 1 0 10764 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_108
timestamp 1649977179
transform 1 0 11040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_122
timestamp 1649977179
transform 1 0 12328 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_132
timestamp 1649977179
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_148
timestamp 1649977179
transform 1 0 14720 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_154
timestamp 1649977179
transform 1 0 15272 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_160
timestamp 1649977179
transform 1 0 15824 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_163
timestamp 1649977179
transform 1 0 16100 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_174
timestamp 1649977179
transform 1 0 17112 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_182
timestamp 1649977179
transform 1 0 17848 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_186
timestamp 1649977179
transform 1 0 18216 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_206
timestamp 1649977179
transform 1 0 20056 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_212
timestamp 1649977179
transform 1 0 20608 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_220
timestamp 1649977179
transform 1 0 21344 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_240
timestamp 1649977179
transform 1 0 23184 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_269
timestamp 1649977179
transform 1 0 25852 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_281
timestamp 1649977179
transform 1 0 26956 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_296
timestamp 1649977179
transform 1 0 28336 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_319
timestamp 1649977179
transform 1 0 30452 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_332
timestamp 1649977179
transform 1 0 31648 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_336
timestamp 1649977179
transform 1 0 32016 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_344
timestamp 1649977179
transform 1 0 32752 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_356
timestamp 1649977179
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_376
timestamp 1649977179
transform 1 0 35696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_396
timestamp 1649977179
transform 1 0 37536 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_407
timestamp 1649977179
transform 1 0 38548 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_413
timestamp 1649977179
transform 1 0 39100 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1649977179
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_421
timestamp 1649977179
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_433
timestamp 1649977179
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_445
timestamp 1649977179
transform 1 0 42044 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_449
timestamp 1649977179
transform 1 0 42412 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_456
timestamp 1649977179
transform 1 0 43056 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_472
timestamp 1649977179
transform 1 0 44528 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_490
timestamp 1649977179
transform 1 0 46184 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_502
timestamp 1649977179
transform 1 0 47288 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_514
timestamp 1649977179
transform 1 0 48392 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_526
timestamp 1649977179
transform 1 0 49496 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_533
timestamp 1649977179
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_545
timestamp 1649977179
transform 1 0 51244 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_557
timestamp 1649977179
transform 1 0 52348 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_569
timestamp 1649977179
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_581
timestamp 1649977179
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_587
timestamp 1649977179
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_589
timestamp 1649977179
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_601
timestamp 1649977179
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_613
timestamp 1649977179
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_625
timestamp 1649977179
transform 1 0 58604 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_637
timestamp 1649977179
transform 1 0 59708 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_643
timestamp 1649977179
transform 1 0 60260 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_645
timestamp 1649977179
transform 1 0 60444 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_657
timestamp 1649977179
transform 1 0 61548 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_669
timestamp 1649977179
transform 1 0 62652 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_681
timestamp 1649977179
transform 1 0 63756 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_693
timestamp 1649977179
transform 1 0 64860 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_699
timestamp 1649977179
transform 1 0 65412 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_701
timestamp 1649977179
transform 1 0 65596 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_713
timestamp 1649977179
transform 1 0 66700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_725
timestamp 1649977179
transform 1 0 67804 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_48
timestamp 1649977179
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_66
timestamp 1649977179
transform 1 0 7176 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_72
timestamp 1649977179
transform 1 0 7728 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_84
timestamp 1649977179
transform 1 0 8832 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_90
timestamp 1649977179
transform 1 0 9384 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_98
timestamp 1649977179
transform 1 0 10120 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_106
timestamp 1649977179
transform 1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_118
timestamp 1649977179
transform 1 0 11960 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_129
timestamp 1649977179
transform 1 0 12972 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_147
timestamp 1649977179
transform 1 0 14628 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_151
timestamp 1649977179
transform 1 0 14996 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_154
timestamp 1649977179
transform 1 0 15272 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1649977179
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_172
timestamp 1649977179
transform 1 0 16928 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_178
timestamp 1649977179
transform 1 0 17480 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_203
timestamp 1649977179
transform 1 0 19780 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_215
timestamp 1649977179
transform 1 0 20884 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_229
timestamp 1649977179
transform 1 0 22172 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_241
timestamp 1649977179
transform 1 0 23276 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_253
timestamp 1649977179
transform 1 0 24380 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_258
timestamp 1649977179
transform 1 0 24840 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_270
timestamp 1649977179
transform 1 0 25944 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1649977179
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_313
timestamp 1649977179
transform 1 0 29900 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1649977179
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_340
timestamp 1649977179
transform 1 0 32384 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_352
timestamp 1649977179
transform 1 0 33488 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_364
timestamp 1649977179
transform 1 0 34592 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_383
timestamp 1649977179
transform 1 0 36340 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_402
timestamp 1649977179
transform 1 0 38088 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_413
timestamp 1649977179
transform 1 0 39100 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_424
timestamp 1649977179
transform 1 0 40112 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_435
timestamp 1649977179
transform 1 0 41124 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1649977179
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_449
timestamp 1649977179
transform 1 0 42412 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_454
timestamp 1649977179
transform 1 0 42872 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_464
timestamp 1649977179
transform 1 0 43792 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_468
timestamp 1649977179
transform 1 0 44160 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_472
timestamp 1649977179
transform 1 0 44528 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_479
timestamp 1649977179
transform 1 0 45172 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_491
timestamp 1649977179
transform 1 0 46276 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1649977179
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1649977179
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_517
timestamp 1649977179
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_529
timestamp 1649977179
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_541
timestamp 1649977179
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_553
timestamp 1649977179
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1649977179
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_561
timestamp 1649977179
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_573
timestamp 1649977179
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_585
timestamp 1649977179
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_597
timestamp 1649977179
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_609
timestamp 1649977179
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_615
timestamp 1649977179
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_617
timestamp 1649977179
transform 1 0 57868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_629
timestamp 1649977179
transform 1 0 58972 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_641
timestamp 1649977179
transform 1 0 60076 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_653
timestamp 1649977179
transform 1 0 61180 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_665
timestamp 1649977179
transform 1 0 62284 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_671
timestamp 1649977179
transform 1 0 62836 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_673
timestamp 1649977179
transform 1 0 63020 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_685
timestamp 1649977179
transform 1 0 64124 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_697
timestamp 1649977179
transform 1 0 65228 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_709
timestamp 1649977179
transform 1 0 66332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_721
timestamp 1649977179
transform 1 0 67436 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_727
timestamp 1649977179
transform 1 0 67988 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_729
timestamp 1649977179
transform 1 0 68172 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_57
timestamp 1649977179
transform 1 0 6348 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_68
timestamp 1649977179
transform 1 0 7360 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_80
timestamp 1649977179
transform 1 0 8464 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_92
timestamp 1649977179
transform 1 0 9568 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_104
timestamp 1649977179
transform 1 0 10672 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_112
timestamp 1649977179
transform 1 0 11408 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_125
timestamp 1649977179
transform 1 0 12604 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_131
timestamp 1649977179
transform 1 0 13156 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_149
timestamp 1649977179
transform 1 0 14812 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_170
timestamp 1649977179
transform 1 0 16744 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_187
timestamp 1649977179
transform 1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_200
timestamp 1649977179
transform 1 0 19504 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_206
timestamp 1649977179
transform 1 0 20056 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_211
timestamp 1649977179
transform 1 0 20516 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_225
timestamp 1649977179
transform 1 0 21804 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_237
timestamp 1649977179
transform 1 0 22908 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1649977179
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_266
timestamp 1649977179
transform 1 0 25576 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_278
timestamp 1649977179
transform 1 0 26680 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_290
timestamp 1649977179
transform 1 0 27784 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_298
timestamp 1649977179
transform 1 0 28520 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1649977179
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_317
timestamp 1649977179
transform 1 0 30268 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_335
timestamp 1649977179
transform 1 0 31924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_347
timestamp 1649977179
transform 1 0 33028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1649977179
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_371
timestamp 1649977179
transform 1 0 35236 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_375
timestamp 1649977179
transform 1 0 35604 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_395
timestamp 1649977179
transform 1 0 37444 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_413
timestamp 1649977179
transform 1 0 39100 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1649977179
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_421
timestamp 1649977179
transform 1 0 39836 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_429
timestamp 1649977179
transform 1 0 40572 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_432
timestamp 1649977179
transform 1 0 40848 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_443
timestamp 1649977179
transform 1 0 41860 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_455
timestamp 1649977179
transform 1 0 42964 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_458
timestamp 1649977179
transform 1 0 43240 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_470
timestamp 1649977179
transform 1 0 44344 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1649977179
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1649977179
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1649977179
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_513
timestamp 1649977179
transform 1 0 48300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_525
timestamp 1649977179
transform 1 0 49404 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1649977179
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_533
timestamp 1649977179
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_545
timestamp 1649977179
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_557
timestamp 1649977179
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_569
timestamp 1649977179
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_581
timestamp 1649977179
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_587
timestamp 1649977179
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_589
timestamp 1649977179
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_601
timestamp 1649977179
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_613
timestamp 1649977179
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_625
timestamp 1649977179
transform 1 0 58604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_637
timestamp 1649977179
transform 1 0 59708 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_643
timestamp 1649977179
transform 1 0 60260 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_645
timestamp 1649977179
transform 1 0 60444 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_657
timestamp 1649977179
transform 1 0 61548 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_669
timestamp 1649977179
transform 1 0 62652 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_681
timestamp 1649977179
transform 1 0 63756 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_693
timestamp 1649977179
transform 1 0 64860 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_699
timestamp 1649977179
transform 1 0 65412 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_701
timestamp 1649977179
transform 1 0 65596 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_713
timestamp 1649977179
transform 1 0 66700 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_717
timestamp 1649977179
transform 1 0 67068 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_721
timestamp 1649977179
transform 1 0 67436 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_727
timestamp 1649977179
transform 1 0 67988 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_99
timestamp 1649977179
transform 1 0 10212 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_107
timestamp 1649977179
transform 1 0 10948 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_116
timestamp 1649977179
transform 1 0 11776 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_128
timestamp 1649977179
transform 1 0 12880 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_140
timestamp 1649977179
transform 1 0 13984 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_148
timestamp 1649977179
transform 1 0 14720 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_151
timestamp 1649977179
transform 1 0 14996 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1649977179
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_172
timestamp 1649977179
transform 1 0 16928 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_178
timestamp 1649977179
transform 1 0 17480 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_186
timestamp 1649977179
transform 1 0 18216 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_192
timestamp 1649977179
transform 1 0 18768 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_198
timestamp 1649977179
transform 1 0 19320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_201
timestamp 1649977179
transform 1 0 19596 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_207
timestamp 1649977179
transform 1 0 20148 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_215
timestamp 1649977179
transform 1 0 20884 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1649977179
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_234
timestamp 1649977179
transform 1 0 22632 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_246
timestamp 1649977179
transform 1 0 23736 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_265
timestamp 1649977179
transform 1 0 25484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_269
timestamp 1649977179
transform 1 0 25852 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_287
timestamp 1649977179
transform 1 0 27508 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_311
timestamp 1649977179
transform 1 0 29716 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_319
timestamp 1649977179
transform 1 0 30452 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_324
timestamp 1649977179
transform 1 0 30912 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1649977179
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_346
timestamp 1649977179
transform 1 0 32936 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_358
timestamp 1649977179
transform 1 0 34040 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_370
timestamp 1649977179
transform 1 0 35144 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_405
timestamp 1649977179
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_417
timestamp 1649977179
transform 1 0 39468 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_431
timestamp 1649977179
transform 1 0 40756 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_444
timestamp 1649977179
transform 1 0 41952 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_465
timestamp 1649977179
transform 1 0 43884 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_477
timestamp 1649977179
transform 1 0 44988 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_489
timestamp 1649977179
transform 1 0 46092 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_501
timestamp 1649977179
transform 1 0 47196 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1649977179
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_517
timestamp 1649977179
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_529
timestamp 1649977179
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_541
timestamp 1649977179
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_553
timestamp 1649977179
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_559
timestamp 1649977179
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_561
timestamp 1649977179
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_573
timestamp 1649977179
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_585
timestamp 1649977179
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_597
timestamp 1649977179
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_609
timestamp 1649977179
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_615
timestamp 1649977179
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_617
timestamp 1649977179
transform 1 0 57868 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_629
timestamp 1649977179
transform 1 0 58972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_641
timestamp 1649977179
transform 1 0 60076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_653
timestamp 1649977179
transform 1 0 61180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_665
timestamp 1649977179
transform 1 0 62284 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_671
timestamp 1649977179
transform 1 0 62836 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_673
timestamp 1649977179
transform 1 0 63020 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_685
timestamp 1649977179
transform 1 0 64124 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_697
timestamp 1649977179
transform 1 0 65228 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_709
timestamp 1649977179
transform 1 0 66332 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_721
timestamp 1649977179
transform 1 0 67436 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_727
timestamp 1649977179
transform 1 0 67988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_729
timestamp 1649977179
transform 1 0 68172 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_47
timestamp 1649977179
transform 1 0 5428 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_67
timestamp 1649977179
transform 1 0 7268 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_80
timestamp 1649977179
transform 1 0 8464 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_87
timestamp 1649977179
transform 1 0 9108 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_99
timestamp 1649977179
transform 1 0 10212 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_143
timestamp 1649977179
transform 1 0 14260 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_149
timestamp 1649977179
transform 1 0 14812 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_152
timestamp 1649977179
transform 1 0 15088 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_159
timestamp 1649977179
transform 1 0 15732 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_170
timestamp 1649977179
transform 1 0 16744 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_179
timestamp 1649977179
transform 1 0 17572 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_192
timestamp 1649977179
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_205
timestamp 1649977179
transform 1 0 19964 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_211
timestamp 1649977179
transform 1 0 20516 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_228
timestamp 1649977179
transform 1 0 22080 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_234
timestamp 1649977179
transform 1 0 22632 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_240
timestamp 1649977179
transform 1 0 23184 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_257
timestamp 1649977179
transform 1 0 24748 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_263
timestamp 1649977179
transform 1 0 25300 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_283
timestamp 1649977179
transform 1 0 27140 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_296
timestamp 1649977179
transform 1 0 28336 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1649977179
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_318
timestamp 1649977179
transform 1 0 30360 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_326
timestamp 1649977179
transform 1 0 31096 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_331
timestamp 1649977179
transform 1 0 31556 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_351
timestamp 1649977179
transform 1 0 33396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_380
timestamp 1649977179
transform 1 0 36064 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_386
timestamp 1649977179
transform 1 0 36616 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_399
timestamp 1649977179
transform 1 0 37812 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_411
timestamp 1649977179
transform 1 0 38916 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1649977179
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_421
timestamp 1649977179
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_433
timestamp 1649977179
transform 1 0 40940 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_452
timestamp 1649977179
transform 1 0 42688 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_464
timestamp 1649977179
transform 1 0 43792 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1649977179
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1649977179
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1649977179
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1649977179
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_525
timestamp 1649977179
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_531
timestamp 1649977179
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_533
timestamp 1649977179
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_545
timestamp 1649977179
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_557
timestamp 1649977179
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_569
timestamp 1649977179
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_581
timestamp 1649977179
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_587
timestamp 1649977179
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_589
timestamp 1649977179
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_601
timestamp 1649977179
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_613
timestamp 1649977179
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_625
timestamp 1649977179
transform 1 0 58604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_637
timestamp 1649977179
transform 1 0 59708 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_643
timestamp 1649977179
transform 1 0 60260 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_645
timestamp 1649977179
transform 1 0 60444 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_657
timestamp 1649977179
transform 1 0 61548 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_669
timestamp 1649977179
transform 1 0 62652 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_681
timestamp 1649977179
transform 1 0 63756 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_693
timestamp 1649977179
transform 1 0 64860 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_699
timestamp 1649977179
transform 1 0 65412 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_701
timestamp 1649977179
transform 1 0 65596 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_713
timestamp 1649977179
transform 1 0 66700 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_725
timestamp 1649977179
transform 1 0 67804 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_35
timestamp 1649977179
transform 1 0 4324 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_52
timestamp 1649977179
transform 1 0 5888 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_73
timestamp 1649977179
transform 1 0 7820 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_80
timestamp 1649977179
transform 1 0 8464 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_84
timestamp 1649977179
transform 1 0 8832 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_92
timestamp 1649977179
transform 1 0 9568 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_102
timestamp 1649977179
transform 1 0 10488 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_110
timestamp 1649977179
transform 1 0 11224 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_128
timestamp 1649977179
transform 1 0 12880 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_141
timestamp 1649977179
transform 1 0 14076 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_151
timestamp 1649977179
transform 1 0 14996 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1649977179
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_202
timestamp 1649977179
transform 1 0 19688 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_210
timestamp 1649977179
transform 1 0 20424 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_219
timestamp 1649977179
transform 1 0 21252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_234
timestamp 1649977179
transform 1 0 22632 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_253
timestamp 1649977179
transform 1 0 24380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_257
timestamp 1649977179
transform 1 0 24748 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_270
timestamp 1649977179
transform 1 0 25944 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1649977179
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_288
timestamp 1649977179
transform 1 0 27600 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_312
timestamp 1649977179
transform 1 0 29808 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_324
timestamp 1649977179
transform 1 0 30912 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_328
timestamp 1649977179
transform 1 0 31280 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_332
timestamp 1649977179
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_346
timestamp 1649977179
transform 1 0 32936 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_352
timestamp 1649977179
transform 1 0 33488 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_372
timestamp 1649977179
transform 1 0 35328 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_379
timestamp 1649977179
transform 1 0 35972 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1649977179
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_409
timestamp 1649977179
transform 1 0 38732 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_421
timestamp 1649977179
transform 1 0 39836 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_427
timestamp 1649977179
transform 1 0 40388 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_440
timestamp 1649977179
transform 1 0 41584 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_452
timestamp 1649977179
transform 1 0 42688 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_464
timestamp 1649977179
transform 1 0 43792 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_476
timestamp 1649977179
transform 1 0 44896 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_488
timestamp 1649977179
transform 1 0 46000 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_500
timestamp 1649977179
transform 1 0 47104 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_505
timestamp 1649977179
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_517
timestamp 1649977179
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_529
timestamp 1649977179
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_541
timestamp 1649977179
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_553
timestamp 1649977179
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_559
timestamp 1649977179
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_561
timestamp 1649977179
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_573
timestamp 1649977179
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_585
timestamp 1649977179
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_597
timestamp 1649977179
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_609
timestamp 1649977179
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_615
timestamp 1649977179
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_617
timestamp 1649977179
transform 1 0 57868 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_629
timestamp 1649977179
transform 1 0 58972 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_641
timestamp 1649977179
transform 1 0 60076 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_653
timestamp 1649977179
transform 1 0 61180 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_665
timestamp 1649977179
transform 1 0 62284 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_671
timestamp 1649977179
transform 1 0 62836 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_673
timestamp 1649977179
transform 1 0 63020 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_685
timestamp 1649977179
transform 1 0 64124 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_697
timestamp 1649977179
transform 1 0 65228 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_709
timestamp 1649977179
transform 1 0 66332 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_721
timestamp 1649977179
transform 1 0 67436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_727
timestamp 1649977179
transform 1 0 67988 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_729
timestamp 1649977179
transform 1 0 68172 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_61
timestamp 1649977179
transform 1 0 6716 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_74
timestamp 1649977179
transform 1 0 7912 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1649977179
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_117
timestamp 1649977179
transform 1 0 11868 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_134
timestamp 1649977179
transform 1 0 13432 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_54_144
timestamp 1649977179
transform 1 0 14352 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_150
timestamp 1649977179
transform 1 0 14904 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_167
timestamp 1649977179
transform 1 0 16468 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_175
timestamp 1649977179
transform 1 0 17204 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1649977179
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_200
timestamp 1649977179
transform 1 0 19504 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_206
timestamp 1649977179
transform 1 0 20056 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_228
timestamp 1649977179
transform 1 0 22080 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1649977179
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_269
timestamp 1649977179
transform 1 0 25852 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_281
timestamp 1649977179
transform 1 0 26956 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_284
timestamp 1649977179
transform 1 0 27232 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_297
timestamp 1649977179
transform 1 0 28428 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1649977179
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_343
timestamp 1649977179
transform 1 0 32660 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_355
timestamp 1649977179
transform 1 0 33764 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_359
timestamp 1649977179
transform 1 0 34132 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_381
timestamp 1649977179
transform 1 0 36156 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_387
timestamp 1649977179
transform 1 0 36708 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_412
timestamp 1649977179
transform 1 0 39008 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_428
timestamp 1649977179
transform 1 0 40480 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_439
timestamp 1649977179
transform 1 0 41492 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_446
timestamp 1649977179
transform 1 0 42136 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_458
timestamp 1649977179
transform 1 0 43240 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_470
timestamp 1649977179
transform 1 0 44344 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1649977179
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1649977179
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_501
timestamp 1649977179
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_513
timestamp 1649977179
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_525
timestamp 1649977179
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_531
timestamp 1649977179
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_533
timestamp 1649977179
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_545
timestamp 1649977179
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_557
timestamp 1649977179
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_569
timestamp 1649977179
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_581
timestamp 1649977179
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_587
timestamp 1649977179
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_589
timestamp 1649977179
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_601
timestamp 1649977179
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_613
timestamp 1649977179
transform 1 0 57500 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_618
timestamp 1649977179
transform 1 0 57960 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_624
timestamp 1649977179
transform 1 0 58512 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_636
timestamp 1649977179
transform 1 0 59616 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_645
timestamp 1649977179
transform 1 0 60444 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_657
timestamp 1649977179
transform 1 0 61548 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_669
timestamp 1649977179
transform 1 0 62652 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_681
timestamp 1649977179
transform 1 0 63756 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_693
timestamp 1649977179
transform 1 0 64860 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_699
timestamp 1649977179
transform 1 0 65412 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_701
timestamp 1649977179
transform 1 0 65596 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_713
timestamp 1649977179
transform 1 0 66700 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_725
timestamp 1649977179
transform 1 0 67804 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_60
timestamp 1649977179
transform 1 0 6624 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_72
timestamp 1649977179
transform 1 0 7728 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_91
timestamp 1649977179
transform 1 0 9476 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_103
timestamp 1649977179
transform 1 0 10580 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_121
timestamp 1649977179
transform 1 0 12236 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_129
timestamp 1649977179
transform 1 0 12972 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_146
timestamp 1649977179
transform 1 0 14536 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_157
timestamp 1649977179
transform 1 0 15548 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_163
timestamp 1649977179
transform 1 0 16100 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_173
timestamp 1649977179
transform 1 0 17020 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_184
timestamp 1649977179
transform 1 0 18032 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_191
timestamp 1649977179
transform 1 0 18676 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_197
timestamp 1649977179
transform 1 0 19228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_209
timestamp 1649977179
transform 1 0 20332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_221
timestamp 1649977179
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_241
timestamp 1649977179
transform 1 0 23276 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_253
timestamp 1649977179
transform 1 0 24380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_259
timestamp 1649977179
transform 1 0 24932 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_266
timestamp 1649977179
transform 1 0 25576 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1649977179
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_289
timestamp 1649977179
transform 1 0 27692 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_297
timestamp 1649977179
transform 1 0 28428 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_304
timestamp 1649977179
transform 1 0 29072 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_316
timestamp 1649977179
transform 1 0 30176 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_328
timestamp 1649977179
transform 1 0 31280 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_355
timestamp 1649977179
transform 1 0 33764 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_368
timestamp 1649977179
transform 1 0 34960 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_381
timestamp 1649977179
transform 1 0 36156 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_388
timestamp 1649977179
transform 1 0 36800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_399
timestamp 1649977179
transform 1 0 37812 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_413
timestamp 1649977179
transform 1 0 39100 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_426
timestamp 1649977179
transform 1 0 40296 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_438
timestamp 1649977179
transform 1 0 41400 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_446
timestamp 1649977179
transform 1 0 42136 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_449
timestamp 1649977179
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_461
timestamp 1649977179
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_473
timestamp 1649977179
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_485
timestamp 1649977179
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1649977179
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1649977179
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_505
timestamp 1649977179
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_517
timestamp 1649977179
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_529
timestamp 1649977179
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_541
timestamp 1649977179
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_553
timestamp 1649977179
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1649977179
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_561
timestamp 1649977179
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_573
timestamp 1649977179
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_585
timestamp 1649977179
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_597
timestamp 1649977179
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_609
timestamp 1649977179
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_615
timestamp 1649977179
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_617
timestamp 1649977179
transform 1 0 57868 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_629
timestamp 1649977179
transform 1 0 58972 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_641
timestamp 1649977179
transform 1 0 60076 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_653
timestamp 1649977179
transform 1 0 61180 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_665
timestamp 1649977179
transform 1 0 62284 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_671
timestamp 1649977179
transform 1 0 62836 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_673
timestamp 1649977179
transform 1 0 63020 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_685
timestamp 1649977179
transform 1 0 64124 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_697
timestamp 1649977179
transform 1 0 65228 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_709
timestamp 1649977179
transform 1 0 66332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_721
timestamp 1649977179
transform 1 0 67436 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_727
timestamp 1649977179
transform 1 0 67988 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_729
timestamp 1649977179
transform 1 0 68172 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_98
timestamp 1649977179
transform 1 0 10120 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_110
timestamp 1649977179
transform 1 0 11224 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_122
timestamp 1649977179
transform 1 0 12328 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_131
timestamp 1649977179
transform 1 0 13156 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_147
timestamp 1649977179
transform 1 0 14628 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_154
timestamp 1649977179
transform 1 0 15272 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_160
timestamp 1649977179
transform 1 0 15824 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_169
timestamp 1649977179
transform 1 0 16652 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_175
timestamp 1649977179
transform 1 0 17204 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_183
timestamp 1649977179
transform 1 0 17940 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_188
timestamp 1649977179
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_199
timestamp 1649977179
transform 1 0 19412 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_211
timestamp 1649977179
transform 1 0 20516 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_219
timestamp 1649977179
transform 1 0 21252 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_224
timestamp 1649977179
transform 1 0 21712 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_234
timestamp 1649977179
transform 1 0 22632 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_246
timestamp 1649977179
transform 1 0 23736 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_257
timestamp 1649977179
transform 1 0 24748 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_266
timestamp 1649977179
transform 1 0 25576 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_273
timestamp 1649977179
transform 1 0 26220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_280
timestamp 1649977179
transform 1 0 26864 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_291
timestamp 1649977179
transform 1 0 27876 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_302
timestamp 1649977179
transform 1 0 28888 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_312
timestamp 1649977179
transform 1 0 29808 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_324
timestamp 1649977179
transform 1 0 30912 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_336
timestamp 1649977179
transform 1 0 32016 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_343
timestamp 1649977179
transform 1 0 32660 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_355
timestamp 1649977179
transform 1 0 33764 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1649977179
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_374
timestamp 1649977179
transform 1 0 35512 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_378
timestamp 1649977179
transform 1 0 35880 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_386
timestamp 1649977179
transform 1 0 36616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_393
timestamp 1649977179
transform 1 0 37260 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_407
timestamp 1649977179
transform 1 0 38548 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1649977179
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_421
timestamp 1649977179
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_433
timestamp 1649977179
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_445
timestamp 1649977179
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_457
timestamp 1649977179
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1649977179
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1649977179
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1649977179
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1649977179
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1649977179
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_513
timestamp 1649977179
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_525
timestamp 1649977179
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1649977179
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_533
timestamp 1649977179
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_545
timestamp 1649977179
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_557
timestamp 1649977179
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_569
timestamp 1649977179
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1649977179
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1649977179
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_589
timestamp 1649977179
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_601
timestamp 1649977179
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_613
timestamp 1649977179
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_625
timestamp 1649977179
transform 1 0 58604 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_637
timestamp 1649977179
transform 1 0 59708 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_643
timestamp 1649977179
transform 1 0 60260 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_645
timestamp 1649977179
transform 1 0 60444 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_657
timestamp 1649977179
transform 1 0 61548 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_669
timestamp 1649977179
transform 1 0 62652 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_681
timestamp 1649977179
transform 1 0 63756 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_693
timestamp 1649977179
transform 1 0 64860 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_699
timestamp 1649977179
transform 1 0 65412 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_701
timestamp 1649977179
transform 1 0 65596 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_713
timestamp 1649977179
transform 1 0 66700 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_725
timestamp 1649977179
transform 1 0 67804 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_88
timestamp 1649977179
transform 1 0 9200 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_100
timestamp 1649977179
transform 1 0 10304 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_133
timestamp 1649977179
transform 1 0 13340 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_142
timestamp 1649977179
transform 1 0 14168 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_155
timestamp 1649977179
transform 1 0 15364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_245
timestamp 1649977179
transform 1 0 23644 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_250
timestamp 1649977179
transform 1 0 24104 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_267
timestamp 1649977179
transform 1 0 25668 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1649977179
transform 1 0 26404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_286
timestamp 1649977179
transform 1 0 27416 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_298
timestamp 1649977179
transform 1 0 28520 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_308
timestamp 1649977179
transform 1 0 29440 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_320
timestamp 1649977179
transform 1 0 30544 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1649977179
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_366
timestamp 1649977179
transform 1 0 34776 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_379
timestamp 1649977179
transform 1 0 35972 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_395
timestamp 1649977179
transform 1 0 37444 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_407
timestamp 1649977179
transform 1 0 38548 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_419
timestamp 1649977179
transform 1 0 39652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_431
timestamp 1649977179
transform 1 0 40756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_443
timestamp 1649977179
transform 1 0 41860 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1649977179
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1649977179
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1649977179
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1649977179
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1649977179
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1649977179
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1649977179
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1649977179
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_517
timestamp 1649977179
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_529
timestamp 1649977179
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_541
timestamp 1649977179
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_553
timestamp 1649977179
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_559
timestamp 1649977179
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_561
timestamp 1649977179
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_573
timestamp 1649977179
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_585
timestamp 1649977179
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_597
timestamp 1649977179
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_609
timestamp 1649977179
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_615
timestamp 1649977179
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_617
timestamp 1649977179
transform 1 0 57868 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_629
timestamp 1649977179
transform 1 0 58972 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_641
timestamp 1649977179
transform 1 0 60076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_653
timestamp 1649977179
transform 1 0 61180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_665
timestamp 1649977179
transform 1 0 62284 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_671
timestamp 1649977179
transform 1 0 62836 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_673
timestamp 1649977179
transform 1 0 63020 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_685
timestamp 1649977179
transform 1 0 64124 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_697
timestamp 1649977179
transform 1 0 65228 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_709
timestamp 1649977179
transform 1 0 66332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_721
timestamp 1649977179
transform 1 0 67436 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_727
timestamp 1649977179
transform 1 0 67988 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_729
timestamp 1649977179
transform 1 0 68172 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_129
timestamp 1649977179
transform 1 0 12972 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_284
timestamp 1649977179
transform 1 0 27232 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_295
timestamp 1649977179
transform 1 0 28244 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_299
timestamp 1649977179
transform 1 0 28612 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_302
timestamp 1649977179
transform 1 0 28888 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1649977179
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1649977179
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1649977179
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_433
timestamp 1649977179
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_445
timestamp 1649977179
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_457
timestamp 1649977179
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1649977179
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1649977179
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1649977179
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1649977179
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1649977179
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_513
timestamp 1649977179
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_525
timestamp 1649977179
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_531
timestamp 1649977179
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_533
timestamp 1649977179
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_545
timestamp 1649977179
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_557
timestamp 1649977179
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_569
timestamp 1649977179
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_581
timestamp 1649977179
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_587
timestamp 1649977179
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_589
timestamp 1649977179
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_601
timestamp 1649977179
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_613
timestamp 1649977179
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_625
timestamp 1649977179
transform 1 0 58604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_637
timestamp 1649977179
transform 1 0 59708 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_643
timestamp 1649977179
transform 1 0 60260 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_645
timestamp 1649977179
transform 1 0 60444 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_657
timestamp 1649977179
transform 1 0 61548 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_669
timestamp 1649977179
transform 1 0 62652 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_681
timestamp 1649977179
transform 1 0 63756 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_693
timestamp 1649977179
transform 1 0 64860 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_699
timestamp 1649977179
transform 1 0 65412 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_701
timestamp 1649977179
transform 1 0 65596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_713
timestamp 1649977179
transform 1 0 66700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_729
timestamp 1649977179
transform 1 0 68172 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_287
timestamp 1649977179
transform 1 0 27508 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_290
timestamp 1649977179
transform 1 0 27784 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_302
timestamp 1649977179
transform 1 0 28888 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_314
timestamp 1649977179
transform 1 0 29992 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_326
timestamp 1649977179
transform 1 0 31096 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1649977179
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_417
timestamp 1649977179
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_429
timestamp 1649977179
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1649977179
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1649977179
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_449
timestamp 1649977179
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_461
timestamp 1649977179
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_473
timestamp 1649977179
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_485
timestamp 1649977179
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_497
timestamp 1649977179
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_503
timestamp 1649977179
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1649977179
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_517
timestamp 1649977179
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_529
timestamp 1649977179
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_541
timestamp 1649977179
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_553
timestamp 1649977179
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_559
timestamp 1649977179
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_561
timestamp 1649977179
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_573
timestamp 1649977179
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_585
timestamp 1649977179
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_597
timestamp 1649977179
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_609
timestamp 1649977179
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_615
timestamp 1649977179
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_617
timestamp 1649977179
transform 1 0 57868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_629
timestamp 1649977179
transform 1 0 58972 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_641
timestamp 1649977179
transform 1 0 60076 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_653
timestamp 1649977179
transform 1 0 61180 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_665
timestamp 1649977179
transform 1 0 62284 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_671
timestamp 1649977179
transform 1 0 62836 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_673
timestamp 1649977179
transform 1 0 63020 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_685
timestamp 1649977179
transform 1 0 64124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_697
timestamp 1649977179
transform 1 0 65228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_709
timestamp 1649977179
transform 1 0 66332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_721
timestamp 1649977179
transform 1 0 67436 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_727
timestamp 1649977179
transform 1 0 67988 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_729
timestamp 1649977179
transform 1 0 68172 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1649977179
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1649977179
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1649977179
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_433
timestamp 1649977179
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_445
timestamp 1649977179
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_457
timestamp 1649977179
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1649977179
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1649977179
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1649977179
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1649977179
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1649977179
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_513
timestamp 1649977179
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1649977179
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1649977179
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_533
timestamp 1649977179
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_545
timestamp 1649977179
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_557
timestamp 1649977179
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_569
timestamp 1649977179
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_581
timestamp 1649977179
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1649977179
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_589
timestamp 1649977179
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_601
timestamp 1649977179
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_613
timestamp 1649977179
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_625
timestamp 1649977179
transform 1 0 58604 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_637
timestamp 1649977179
transform 1 0 59708 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_643
timestamp 1649977179
transform 1 0 60260 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_645
timestamp 1649977179
transform 1 0 60444 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_657
timestamp 1649977179
transform 1 0 61548 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_669
timestamp 1649977179
transform 1 0 62652 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_681
timestamp 1649977179
transform 1 0 63756 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_693
timestamp 1649977179
transform 1 0 64860 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_699
timestamp 1649977179
transform 1 0 65412 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_701
timestamp 1649977179
transform 1 0 65596 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_713
timestamp 1649977179
transform 1 0 66700 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_725
timestamp 1649977179
transform 1 0 67804 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1649977179
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1649977179
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_417
timestamp 1649977179
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_429
timestamp 1649977179
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1649977179
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1649977179
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_449
timestamp 1649977179
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_461
timestamp 1649977179
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_473
timestamp 1649977179
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_485
timestamp 1649977179
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1649977179
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1649977179
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1649977179
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_517
timestamp 1649977179
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_529
timestamp 1649977179
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_541
timestamp 1649977179
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_553
timestamp 1649977179
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_559
timestamp 1649977179
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_561
timestamp 1649977179
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_573
timestamp 1649977179
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_585
timestamp 1649977179
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_597
timestamp 1649977179
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1649977179
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1649977179
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_617
timestamp 1649977179
transform 1 0 57868 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_629
timestamp 1649977179
transform 1 0 58972 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_641
timestamp 1649977179
transform 1 0 60076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_653
timestamp 1649977179
transform 1 0 61180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_665
timestamp 1649977179
transform 1 0 62284 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_671
timestamp 1649977179
transform 1 0 62836 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_673
timestamp 1649977179
transform 1 0 63020 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_685
timestamp 1649977179
transform 1 0 64124 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_697
timestamp 1649977179
transform 1 0 65228 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_709
timestamp 1649977179
transform 1 0 66332 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_721
timestamp 1649977179
transform 1 0 67436 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_727
timestamp 1649977179
transform 1 0 67988 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_729
timestamp 1649977179
transform 1 0 68172 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_401
timestamp 1649977179
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1649977179
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1649977179
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_421
timestamp 1649977179
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_433
timestamp 1649977179
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_445
timestamp 1649977179
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_457
timestamp 1649977179
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1649977179
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1649977179
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1649977179
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1649977179
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1649977179
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1649977179
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_525
timestamp 1649977179
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1649977179
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_533
timestamp 1649977179
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_545
timestamp 1649977179
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_557
timestamp 1649977179
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_569
timestamp 1649977179
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1649977179
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1649977179
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_589
timestamp 1649977179
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_601
timestamp 1649977179
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_613
timestamp 1649977179
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_625
timestamp 1649977179
transform 1 0 58604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_637
timestamp 1649977179
transform 1 0 59708 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_643
timestamp 1649977179
transform 1 0 60260 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_645
timestamp 1649977179
transform 1 0 60444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_657
timestamp 1649977179
transform 1 0 61548 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_669
timestamp 1649977179
transform 1 0 62652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_681
timestamp 1649977179
transform 1 0 63756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_693
timestamp 1649977179
transform 1 0 64860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_699
timestamp 1649977179
transform 1 0 65412 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_701
timestamp 1649977179
transform 1 0 65596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_713
timestamp 1649977179
transform 1 0 66700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_725
timestamp 1649977179
transform 1 0 67804 0 1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_417
timestamp 1649977179
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_429
timestamp 1649977179
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1649977179
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1649977179
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_449
timestamp 1649977179
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_461
timestamp 1649977179
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_473
timestamp 1649977179
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_485
timestamp 1649977179
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_497
timestamp 1649977179
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_503
timestamp 1649977179
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1649977179
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_517
timestamp 1649977179
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_529
timestamp 1649977179
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_541
timestamp 1649977179
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_553
timestamp 1649977179
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_559
timestamp 1649977179
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_561
timestamp 1649977179
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_573
timestamp 1649977179
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_585
timestamp 1649977179
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_597
timestamp 1649977179
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_609
timestamp 1649977179
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_615
timestamp 1649977179
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_617
timestamp 1649977179
transform 1 0 57868 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_629
timestamp 1649977179
transform 1 0 58972 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_641
timestamp 1649977179
transform 1 0 60076 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_653
timestamp 1649977179
transform 1 0 61180 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_665
timestamp 1649977179
transform 1 0 62284 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_671
timestamp 1649977179
transform 1 0 62836 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_673
timestamp 1649977179
transform 1 0 63020 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_685
timestamp 1649977179
transform 1 0 64124 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_697
timestamp 1649977179
transform 1 0 65228 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_709
timestamp 1649977179
transform 1 0 66332 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_721
timestamp 1649977179
transform 1 0 67436 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_727
timestamp 1649977179
transform 1 0 67988 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_729
timestamp 1649977179
transform 1 0 68172 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1649977179
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1649977179
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1649977179
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_233
timestamp 1649977179
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_245
timestamp 1649977179
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_401
timestamp 1649977179
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1649977179
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1649977179
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_421
timestamp 1649977179
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_433
timestamp 1649977179
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_445
timestamp 1649977179
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_457
timestamp 1649977179
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1649977179
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1649977179
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1649977179
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1649977179
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_501
timestamp 1649977179
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_513
timestamp 1649977179
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1649977179
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1649977179
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_533
timestamp 1649977179
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_545
timestamp 1649977179
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_557
timestamp 1649977179
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_569
timestamp 1649977179
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1649977179
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1649977179
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_589
timestamp 1649977179
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_601
timestamp 1649977179
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_613
timestamp 1649977179
transform 1 0 57500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_625
timestamp 1649977179
transform 1 0 58604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_637
timestamp 1649977179
transform 1 0 59708 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_643
timestamp 1649977179
transform 1 0 60260 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_645
timestamp 1649977179
transform 1 0 60444 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_657
timestamp 1649977179
transform 1 0 61548 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_669
timestamp 1649977179
transform 1 0 62652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_681
timestamp 1649977179
transform 1 0 63756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_693
timestamp 1649977179
transform 1 0 64860 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_699
timestamp 1649977179
transform 1 0 65412 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_701
timestamp 1649977179
transform 1 0 65596 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_713
timestamp 1649977179
transform 1 0 66700 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_725
timestamp 1649977179
transform 1 0 67804 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1649977179
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1649977179
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1649977179
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1649977179
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1649977179
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1649977179
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1649977179
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1649977179
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1649977179
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1649977179
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1649977179
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1649977179
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1649977179
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1649977179
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1649977179
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_405
timestamp 1649977179
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_417
timestamp 1649977179
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_429
timestamp 1649977179
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1649977179
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1649977179
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_449
timestamp 1649977179
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_461
timestamp 1649977179
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_473
timestamp 1649977179
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_485
timestamp 1649977179
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_497
timestamp 1649977179
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_503
timestamp 1649977179
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1649977179
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_517
timestamp 1649977179
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_529
timestamp 1649977179
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_541
timestamp 1649977179
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_553
timestamp 1649977179
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_559
timestamp 1649977179
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_561
timestamp 1649977179
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_573
timestamp 1649977179
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_585
timestamp 1649977179
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_597
timestamp 1649977179
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_609
timestamp 1649977179
transform 1 0 57132 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_615
timestamp 1649977179
transform 1 0 57684 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_617
timestamp 1649977179
transform 1 0 57868 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_629
timestamp 1649977179
transform 1 0 58972 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_641
timestamp 1649977179
transform 1 0 60076 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_653
timestamp 1649977179
transform 1 0 61180 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_665
timestamp 1649977179
transform 1 0 62284 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_671
timestamp 1649977179
transform 1 0 62836 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_673
timestamp 1649977179
transform 1 0 63020 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_685
timestamp 1649977179
transform 1 0 64124 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_697
timestamp 1649977179
transform 1 0 65228 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_709
timestamp 1649977179
transform 1 0 66332 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_721
timestamp 1649977179
transform 1 0 67436 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_727
timestamp 1649977179
transform 1 0 67988 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_729
timestamp 1649977179
transform 1 0 68172 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1649977179
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1649977179
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_233
timestamp 1649977179
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1649977179
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1649977179
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1649977179
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_401
timestamp 1649977179
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1649977179
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1649977179
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_421
timestamp 1649977179
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_433
timestamp 1649977179
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_445
timestamp 1649977179
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_457
timestamp 1649977179
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1649977179
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1649977179
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1649977179
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1649977179
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1649977179
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_513
timestamp 1649977179
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_525
timestamp 1649977179
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_531
timestamp 1649977179
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_533
timestamp 1649977179
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_545
timestamp 1649977179
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_557
timestamp 1649977179
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_569
timestamp 1649977179
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_581
timestamp 1649977179
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_587
timestamp 1649977179
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_589
timestamp 1649977179
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_601
timestamp 1649977179
transform 1 0 56396 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_613
timestamp 1649977179
transform 1 0 57500 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_625
timestamp 1649977179
transform 1 0 58604 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_637
timestamp 1649977179
transform 1 0 59708 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_643
timestamp 1649977179
transform 1 0 60260 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_645
timestamp 1649977179
transform 1 0 60444 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_657
timestamp 1649977179
transform 1 0 61548 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_669
timestamp 1649977179
transform 1 0 62652 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_681
timestamp 1649977179
transform 1 0 63756 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_693
timestamp 1649977179
transform 1 0 64860 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_699
timestamp 1649977179
transform 1 0 65412 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_701
timestamp 1649977179
transform 1 0 65596 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_713
timestamp 1649977179
transform 1 0 66700 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_725
timestamp 1649977179
transform 1 0 67804 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1649977179
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1649977179
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1649977179
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1649977179
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1649977179
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1649977179
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1649977179
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_225
timestamp 1649977179
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_237
timestamp 1649977179
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_249
timestamp 1649977179
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_261
timestamp 1649977179
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_273
timestamp 1649977179
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1649977179
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1649977179
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_393
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_405
timestamp 1649977179
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_417
timestamp 1649977179
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_429
timestamp 1649977179
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1649977179
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1649977179
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1649977179
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1649977179
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1649977179
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1649977179
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1649977179
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1649977179
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1649977179
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_517
timestamp 1649977179
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_529
timestamp 1649977179
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_541
timestamp 1649977179
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_553
timestamp 1649977179
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_559
timestamp 1649977179
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_561
timestamp 1649977179
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_573
timestamp 1649977179
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_585
timestamp 1649977179
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_597
timestamp 1649977179
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_609
timestamp 1649977179
transform 1 0 57132 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_615
timestamp 1649977179
transform 1 0 57684 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_617
timestamp 1649977179
transform 1 0 57868 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_629
timestamp 1649977179
transform 1 0 58972 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_641
timestamp 1649977179
transform 1 0 60076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_653
timestamp 1649977179
transform 1 0 61180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_665
timestamp 1649977179
transform 1 0 62284 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_671
timestamp 1649977179
transform 1 0 62836 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_673
timestamp 1649977179
transform 1 0 63020 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_685
timestamp 1649977179
transform 1 0 64124 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_697
timestamp 1649977179
transform 1 0 65228 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_709
timestamp 1649977179
transform 1 0 66332 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_721
timestamp 1649977179
transform 1 0 67436 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_727
timestamp 1649977179
transform 1 0 67988 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_729
timestamp 1649977179
transform 1 0 68172 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1649977179
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1649977179
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1649977179
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1649977179
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_221
timestamp 1649977179
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_233
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_245
timestamp 1649977179
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1649977179
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1649977179
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1649977179
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1649977179
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1649977179
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_421
timestamp 1649977179
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_433
timestamp 1649977179
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_445
timestamp 1649977179
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_457
timestamp 1649977179
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1649977179
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1649977179
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1649977179
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1649977179
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1649977179
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_513
timestamp 1649977179
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_525
timestamp 1649977179
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_531
timestamp 1649977179
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_533
timestamp 1649977179
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_545
timestamp 1649977179
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_557
timestamp 1649977179
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_569
timestamp 1649977179
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_581
timestamp 1649977179
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_587
timestamp 1649977179
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_589
timestamp 1649977179
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_601
timestamp 1649977179
transform 1 0 56396 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_613
timestamp 1649977179
transform 1 0 57500 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_625
timestamp 1649977179
transform 1 0 58604 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_637
timestamp 1649977179
transform 1 0 59708 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_643
timestamp 1649977179
transform 1 0 60260 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_645
timestamp 1649977179
transform 1 0 60444 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_657
timestamp 1649977179
transform 1 0 61548 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_669
timestamp 1649977179
transform 1 0 62652 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_681
timestamp 1649977179
transform 1 0 63756 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_693
timestamp 1649977179
transform 1 0 64860 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_699
timestamp 1649977179
transform 1 0 65412 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_701
timestamp 1649977179
transform 1 0 65596 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_713
timestamp 1649977179
transform 1 0 66700 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_717
timestamp 1649977179
transform 1 0 67068 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_721
timestamp 1649977179
transform 1 0 67436 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_727
timestamp 1649977179
transform 1 0 67988 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1649977179
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1649977179
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1649977179
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1649977179
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1649977179
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1649977179
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_405
timestamp 1649977179
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_417
timestamp 1649977179
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_429
timestamp 1649977179
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1649977179
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1649977179
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1649977179
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1649977179
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1649977179
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1649977179
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1649977179
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1649977179
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_505
timestamp 1649977179
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_517
timestamp 1649977179
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_529
timestamp 1649977179
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_541
timestamp 1649977179
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_553
timestamp 1649977179
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_559
timestamp 1649977179
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_561
timestamp 1649977179
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_573
timestamp 1649977179
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_585
timestamp 1649977179
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_597
timestamp 1649977179
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_609
timestamp 1649977179
transform 1 0 57132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_615
timestamp 1649977179
transform 1 0 57684 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_617
timestamp 1649977179
transform 1 0 57868 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_629
timestamp 1649977179
transform 1 0 58972 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_641
timestamp 1649977179
transform 1 0 60076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_653
timestamp 1649977179
transform 1 0 61180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_665
timestamp 1649977179
transform 1 0 62284 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_671
timestamp 1649977179
transform 1 0 62836 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_673
timestamp 1649977179
transform 1 0 63020 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_685
timestamp 1649977179
transform 1 0 64124 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_697
timestamp 1649977179
transform 1 0 65228 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_709
timestamp 1649977179
transform 1 0 66332 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_721
timestamp 1649977179
transform 1 0 67436 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_727
timestamp 1649977179
transform 1 0 67988 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_729
timestamp 1649977179
transform 1 0 68172 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1649977179
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1649977179
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_401
timestamp 1649977179
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1649977179
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1649977179
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1649977179
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1649977179
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1649977179
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1649977179
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1649977179
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1649977179
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1649977179
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1649977179
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1649977179
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_513
timestamp 1649977179
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_525
timestamp 1649977179
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_531
timestamp 1649977179
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_533
timestamp 1649977179
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_545
timestamp 1649977179
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_557
timestamp 1649977179
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_569
timestamp 1649977179
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_581
timestamp 1649977179
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_587
timestamp 1649977179
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_589
timestamp 1649977179
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_601
timestamp 1649977179
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_613
timestamp 1649977179
transform 1 0 57500 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_625
timestamp 1649977179
transform 1 0 58604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_637
timestamp 1649977179
transform 1 0 59708 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_643
timestamp 1649977179
transform 1 0 60260 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_645
timestamp 1649977179
transform 1 0 60444 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_657
timestamp 1649977179
transform 1 0 61548 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_669
timestamp 1649977179
transform 1 0 62652 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_681
timestamp 1649977179
transform 1 0 63756 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_693
timestamp 1649977179
transform 1 0 64860 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_699
timestamp 1649977179
transform 1 0 65412 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_701
timestamp 1649977179
transform 1 0 65596 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_713
timestamp 1649977179
transform 1 0 66700 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_725
timestamp 1649977179
transform 1 0 67804 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1649977179
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1649977179
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1649977179
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_39
timestamp 1649977179
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1649977179
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1649977179
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_217
timestamp 1649977179
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1649977179
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1649977179
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_281
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_293
timestamp 1649977179
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_305
timestamp 1649977179
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1649977179
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1649977179
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1649977179
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_405
timestamp 1649977179
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_417
timestamp 1649977179
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_429
timestamp 1649977179
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1649977179
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1649977179
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1649977179
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1649977179
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1649977179
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1649977179
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1649977179
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1649977179
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_505
timestamp 1649977179
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_517
timestamp 1649977179
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_529
timestamp 1649977179
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_541
timestamp 1649977179
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_553
timestamp 1649977179
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_559
timestamp 1649977179
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_561
timestamp 1649977179
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_573
timestamp 1649977179
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_585
timestamp 1649977179
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_597
timestamp 1649977179
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_609
timestamp 1649977179
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_615
timestamp 1649977179
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_617
timestamp 1649977179
transform 1 0 57868 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_629
timestamp 1649977179
transform 1 0 58972 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_641
timestamp 1649977179
transform 1 0 60076 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_653
timestamp 1649977179
transform 1 0 61180 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_665
timestamp 1649977179
transform 1 0 62284 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_671
timestamp 1649977179
transform 1 0 62836 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_673
timestamp 1649977179
transform 1 0 63020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_685
timestamp 1649977179
transform 1 0 64124 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_697
timestamp 1649977179
transform 1 0 65228 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_709
timestamp 1649977179
transform 1 0 66332 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_721
timestamp 1649977179
transform 1 0 67436 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_727
timestamp 1649977179
transform 1 0 67988 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_729
timestamp 1649977179
transform 1 0 68172 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_15
timestamp 1649977179
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_221
timestamp 1649977179
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_233
timestamp 1649977179
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_245
timestamp 1649977179
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1649977179
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_401
timestamp 1649977179
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1649977179
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1649977179
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1649977179
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1649977179
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1649977179
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1649977179
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1649977179
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1649977179
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1649977179
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1649977179
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1649977179
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_513
timestamp 1649977179
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_525
timestamp 1649977179
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_531
timestamp 1649977179
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_533
timestamp 1649977179
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_545
timestamp 1649977179
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_557
timestamp 1649977179
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_569
timestamp 1649977179
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_581
timestamp 1649977179
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_587
timestamp 1649977179
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_589
timestamp 1649977179
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_601
timestamp 1649977179
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_613
timestamp 1649977179
transform 1 0 57500 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_625
timestamp 1649977179
transform 1 0 58604 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_637
timestamp 1649977179
transform 1 0 59708 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_643
timestamp 1649977179
transform 1 0 60260 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_645
timestamp 1649977179
transform 1 0 60444 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_657
timestamp 1649977179
transform 1 0 61548 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_669
timestamp 1649977179
transform 1 0 62652 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_681
timestamp 1649977179
transform 1 0 63756 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_693
timestamp 1649977179
transform 1 0 64860 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_699
timestamp 1649977179
transform 1 0 65412 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_701
timestamp 1649977179
transform 1 0 65596 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_713
timestamp 1649977179
transform 1 0 66700 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_721
timestamp 1649977179
transform 1 0 67436 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_729
timestamp 1649977179
transform 1 0 68172 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1649977179
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1649977179
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1649977179
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1649977179
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1649977179
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_293
timestamp 1649977179
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_305
timestamp 1649977179
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_317
timestamp 1649977179
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1649977179
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1649977179
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_417
timestamp 1649977179
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_429
timestamp 1649977179
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1649977179
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1649977179
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1649977179
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1649977179
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1649977179
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1649977179
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1649977179
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1649977179
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_505
timestamp 1649977179
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_517
timestamp 1649977179
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_529
timestamp 1649977179
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_541
timestamp 1649977179
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_553
timestamp 1649977179
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_559
timestamp 1649977179
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_561
timestamp 1649977179
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_573
timestamp 1649977179
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_585
timestamp 1649977179
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_597
timestamp 1649977179
transform 1 0 56028 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_609
timestamp 1649977179
transform 1 0 57132 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_615
timestamp 1649977179
transform 1 0 57684 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_617
timestamp 1649977179
transform 1 0 57868 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_629
timestamp 1649977179
transform 1 0 58972 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_641
timestamp 1649977179
transform 1 0 60076 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_653
timestamp 1649977179
transform 1 0 61180 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_665
timestamp 1649977179
transform 1 0 62284 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_671
timestamp 1649977179
transform 1 0 62836 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_673
timestamp 1649977179
transform 1 0 63020 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_685
timestamp 1649977179
transform 1 0 64124 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_697
timestamp 1649977179
transform 1 0 65228 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_709
timestamp 1649977179
transform 1 0 66332 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_721
timestamp 1649977179
transform 1 0 67436 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_727
timestamp 1649977179
transform 1 0 67988 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_729
timestamp 1649977179
transform 1 0 68172 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1649977179
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1649977179
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1649977179
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1649977179
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1649977179
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1649977179
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1649977179
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1649977179
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_289
timestamp 1649977179
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1649977179
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_401
timestamp 1649977179
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1649977179
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1649977179
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_421
timestamp 1649977179
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_433
timestamp 1649977179
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_445
timestamp 1649977179
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_457
timestamp 1649977179
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1649977179
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1649977179
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1649977179
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1649977179
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1649977179
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_513
timestamp 1649977179
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_525
timestamp 1649977179
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_531
timestamp 1649977179
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_533
timestamp 1649977179
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_545
timestamp 1649977179
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_557
timestamp 1649977179
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_569
timestamp 1649977179
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_581
timestamp 1649977179
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_587
timestamp 1649977179
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_589
timestamp 1649977179
transform 1 0 55292 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_601
timestamp 1649977179
transform 1 0 56396 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_613
timestamp 1649977179
transform 1 0 57500 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_625
timestamp 1649977179
transform 1 0 58604 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_637
timestamp 1649977179
transform 1 0 59708 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_643
timestamp 1649977179
transform 1 0 60260 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_645
timestamp 1649977179
transform 1 0 60444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_657
timestamp 1649977179
transform 1 0 61548 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_669
timestamp 1649977179
transform 1 0 62652 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_681
timestamp 1649977179
transform 1 0 63756 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1649977179
transform 1 0 64860 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1649977179
transform 1 0 65412 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_701
timestamp 1649977179
transform 1 0 65596 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_713
timestamp 1649977179
transform 1 0 66700 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_725
timestamp 1649977179
transform 1 0 67804 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_3
timestamp 1649977179
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_15
timestamp 1649977179
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_27
timestamp 1649977179
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_39
timestamp 1649977179
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1649977179
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_293
timestamp 1649977179
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_305
timestamp 1649977179
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_317
timestamp 1649977179
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1649977179
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1649977179
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1649977179
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_417
timestamp 1649977179
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_429
timestamp 1649977179
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1649977179
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1649977179
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1649977179
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1649977179
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1649977179
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1649977179
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1649977179
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1649977179
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_505
timestamp 1649977179
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_517
timestamp 1649977179
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_529
timestamp 1649977179
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_541
timestamp 1649977179
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_553
timestamp 1649977179
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_559
timestamp 1649977179
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_561
timestamp 1649977179
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_573
timestamp 1649977179
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_585
timestamp 1649977179
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_597
timestamp 1649977179
transform 1 0 56028 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_609
timestamp 1649977179
transform 1 0 57132 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_615
timestamp 1649977179
transform 1 0 57684 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_617
timestamp 1649977179
transform 1 0 57868 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_629
timestamp 1649977179
transform 1 0 58972 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_641
timestamp 1649977179
transform 1 0 60076 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_653
timestamp 1649977179
transform 1 0 61180 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_665
timestamp 1649977179
transform 1 0 62284 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_671
timestamp 1649977179
transform 1 0 62836 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_673
timestamp 1649977179
transform 1 0 63020 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_685
timestamp 1649977179
transform 1 0 64124 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_697
timestamp 1649977179
transform 1 0 65228 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_709
timestamp 1649977179
transform 1 0 66332 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_721
timestamp 1649977179
transform 1 0 67436 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_727
timestamp 1649977179
transform 1 0 67988 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_729
timestamp 1649977179
transform 1 0 68172 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_3
timestamp 1649977179
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_15
timestamp 1649977179
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1649977179
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_289
timestamp 1649977179
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_301
timestamp 1649977179
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_307
timestamp 1649977179
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1649977179
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1649977179
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_401
timestamp 1649977179
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1649977179
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1649977179
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1649977179
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1649977179
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1649977179
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1649977179
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1649977179
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1649977179
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1649977179
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1649977179
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1649977179
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_513
timestamp 1649977179
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_525
timestamp 1649977179
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_531
timestamp 1649977179
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_533
timestamp 1649977179
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_545
timestamp 1649977179
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_557
timestamp 1649977179
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_569
timestamp 1649977179
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_581
timestamp 1649977179
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_587
timestamp 1649977179
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_589
timestamp 1649977179
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_601
timestamp 1649977179
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_613
timestamp 1649977179
transform 1 0 57500 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_625
timestamp 1649977179
transform 1 0 58604 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_637
timestamp 1649977179
transform 1 0 59708 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_643
timestamp 1649977179
transform 1 0 60260 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_645
timestamp 1649977179
transform 1 0 60444 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_657
timestamp 1649977179
transform 1 0 61548 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_669
timestamp 1649977179
transform 1 0 62652 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_681
timestamp 1649977179
transform 1 0 63756 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_693
timestamp 1649977179
transform 1 0 64860 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_699
timestamp 1649977179
transform 1 0 65412 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_701
timestamp 1649977179
transform 1 0 65596 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_713
timestamp 1649977179
transform 1 0 66700 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_725
timestamp 1649977179
transform 1 0 67804 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1649977179
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1649977179
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1649977179
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1649977179
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1649977179
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1649977179
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1649977179
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1649977179
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1649977179
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1649977179
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1649977179
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1649977179
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_373
timestamp 1649977179
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1649977179
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1649977179
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1649977179
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_405
timestamp 1649977179
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_417
timestamp 1649977179
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_429
timestamp 1649977179
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1649977179
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1649977179
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1649977179
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1649977179
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1649977179
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1649977179
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1649977179
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1649977179
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1649977179
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_517
timestamp 1649977179
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_529
timestamp 1649977179
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_541
timestamp 1649977179
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_553
timestamp 1649977179
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_559
timestamp 1649977179
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_561
timestamp 1649977179
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_573
timestamp 1649977179
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_585
timestamp 1649977179
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_597
timestamp 1649977179
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_609
timestamp 1649977179
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_615
timestamp 1649977179
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_617
timestamp 1649977179
transform 1 0 57868 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_629
timestamp 1649977179
transform 1 0 58972 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_641
timestamp 1649977179
transform 1 0 60076 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_653
timestamp 1649977179
transform 1 0 61180 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_665
timestamp 1649977179
transform 1 0 62284 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_671
timestamp 1649977179
transform 1 0 62836 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_673
timestamp 1649977179
transform 1 0 63020 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_685
timestamp 1649977179
transform 1 0 64124 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_697
timestamp 1649977179
transform 1 0 65228 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_709
timestamp 1649977179
transform 1 0 66332 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_721
timestamp 1649977179
transform 1 0 67436 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_727
timestamp 1649977179
transform 1 0 67988 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_729
timestamp 1649977179
transform 1 0 68172 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1649977179
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1649977179
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1649977179
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1649977179
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1649977179
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1649977179
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1649977179
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1649977179
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1649977179
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1649977179
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1649977179
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1649977179
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_377
timestamp 1649977179
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_389
timestamp 1649977179
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_401
timestamp 1649977179
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1649977179
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1649977179
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1649977179
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1649977179
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1649977179
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1649977179
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1649977179
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1649977179
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1649977179
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1649977179
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1649977179
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_513
timestamp 1649977179
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_525
timestamp 1649977179
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_531
timestamp 1649977179
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_533
timestamp 1649977179
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_545
timestamp 1649977179
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_557
timestamp 1649977179
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_569
timestamp 1649977179
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_581
timestamp 1649977179
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_587
timestamp 1649977179
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_589
timestamp 1649977179
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_601
timestamp 1649977179
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_613
timestamp 1649977179
transform 1 0 57500 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_625
timestamp 1649977179
transform 1 0 58604 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_637
timestamp 1649977179
transform 1 0 59708 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_643
timestamp 1649977179
transform 1 0 60260 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_645
timestamp 1649977179
transform 1 0 60444 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_657
timestamp 1649977179
transform 1 0 61548 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_669
timestamp 1649977179
transform 1 0 62652 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_681
timestamp 1649977179
transform 1 0 63756 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_693
timestamp 1649977179
transform 1 0 64860 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_699
timestamp 1649977179
transform 1 0 65412 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_701
timestamp 1649977179
transform 1 0 65596 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_713
timestamp 1649977179
transform 1 0 66700 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_725
timestamp 1649977179
transform 1 0 67804 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1649977179
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1649977179
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1649977179
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1649977179
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1649977179
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_149
timestamp 1649977179
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1649977179
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1649977179
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1649977179
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1649977179
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1649977179
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1649977179
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1649977179
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1649977179
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1649977179
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1649977179
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1649977179
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1649977179
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1649977179
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1649977179
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1649977179
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1649977179
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1649977179
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1649977179
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1649977179
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1649977179
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1649977179
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_505
timestamp 1649977179
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_517
timestamp 1649977179
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_529
timestamp 1649977179
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_541
timestamp 1649977179
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_553
timestamp 1649977179
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_559
timestamp 1649977179
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_561
timestamp 1649977179
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_573
timestamp 1649977179
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_585
timestamp 1649977179
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_597
timestamp 1649977179
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_609
timestamp 1649977179
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_615
timestamp 1649977179
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_617
timestamp 1649977179
transform 1 0 57868 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_629
timestamp 1649977179
transform 1 0 58972 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_641
timestamp 1649977179
transform 1 0 60076 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_653
timestamp 1649977179
transform 1 0 61180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_665
timestamp 1649977179
transform 1 0 62284 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_671
timestamp 1649977179
transform 1 0 62836 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_673
timestamp 1649977179
transform 1 0 63020 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_685
timestamp 1649977179
transform 1 0 64124 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_697
timestamp 1649977179
transform 1 0 65228 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_709
timestamp 1649977179
transform 1 0 66332 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_714
timestamp 1649977179
transform 1 0 66792 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_721
timestamp 1649977179
transform 1 0 67436 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_727
timestamp 1649977179
transform 1 0 67988 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_729
timestamp 1649977179
transform 1 0 68172 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_80_3
timestamp 1649977179
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1649977179
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1649977179
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1649977179
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1649977179
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1649977179
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1649977179
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1649977179
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1649977179
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1649977179
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1649977179
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1649977179
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_197
timestamp 1649977179
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_209
timestamp 1649977179
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_221
timestamp 1649977179
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_233
timestamp 1649977179
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1649977179
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1649977179
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1649977179
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_277
timestamp 1649977179
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_289
timestamp 1649977179
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1649977179
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1649977179
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1649977179
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1649977179
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1649977179
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1649977179
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1649977179
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1649977179
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1649977179
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1649977179
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1649977179
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1649977179
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1649977179
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1649977179
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1649977179
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1649977179
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1649977179
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_501
timestamp 1649977179
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_513
timestamp 1649977179
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_525
timestamp 1649977179
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_531
timestamp 1649977179
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_533
timestamp 1649977179
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_545
timestamp 1649977179
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_557
timestamp 1649977179
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_569
timestamp 1649977179
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_581
timestamp 1649977179
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_587
timestamp 1649977179
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_589
timestamp 1649977179
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_601
timestamp 1649977179
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_613
timestamp 1649977179
transform 1 0 57500 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_625
timestamp 1649977179
transform 1 0 58604 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_637
timestamp 1649977179
transform 1 0 59708 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_643
timestamp 1649977179
transform 1 0 60260 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_645
timestamp 1649977179
transform 1 0 60444 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_657
timestamp 1649977179
transform 1 0 61548 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_669
timestamp 1649977179
transform 1 0 62652 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_681
timestamp 1649977179
transform 1 0 63756 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_693
timestamp 1649977179
transform 1 0 64860 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_699
timestamp 1649977179
transform 1 0 65412 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_701
timestamp 1649977179
transform 1 0 65596 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_713
timestamp 1649977179
transform 1 0 66700 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_725
timestamp 1649977179
transform 1 0 67804 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1649977179
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1649977179
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1649977179
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1649977179
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1649977179
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1649977179
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1649977179
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1649977179
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1649977179
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1649977179
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1649977179
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1649977179
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1649977179
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1649977179
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1649977179
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1649977179
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1649977179
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1649977179
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1649977179
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1649977179
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1649977179
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1649977179
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1649977179
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1649977179
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1649977179
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1649977179
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1649977179
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1649977179
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1649977179
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1649977179
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1649977179
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1649977179
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1649977179
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1649977179
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1649977179
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1649977179
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1649977179
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1649977179
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1649977179
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1649977179
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1649977179
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1649977179
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1649977179
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1649977179
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1649977179
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1649977179
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_517
timestamp 1649977179
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_529
timestamp 1649977179
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_541
timestamp 1649977179
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_553
timestamp 1649977179
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_559
timestamp 1649977179
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_561
timestamp 1649977179
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_573
timestamp 1649977179
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_585
timestamp 1649977179
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_597
timestamp 1649977179
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_609
timestamp 1649977179
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_615
timestamp 1649977179
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_617
timestamp 1649977179
transform 1 0 57868 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_629
timestamp 1649977179
transform 1 0 58972 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_641
timestamp 1649977179
transform 1 0 60076 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_653
timestamp 1649977179
transform 1 0 61180 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_665
timestamp 1649977179
transform 1 0 62284 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_671
timestamp 1649977179
transform 1 0 62836 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_673
timestamp 1649977179
transform 1 0 63020 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_685
timestamp 1649977179
transform 1 0 64124 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_697
timestamp 1649977179
transform 1 0 65228 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_709
timestamp 1649977179
transform 1 0 66332 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_721
timestamp 1649977179
transform 1 0 67436 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_727
timestamp 1649977179
transform 1 0 67988 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_729
timestamp 1649977179
transform 1 0 68172 0 -1 46784
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1649977179
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1649977179
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1649977179
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1649977179
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1649977179
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1649977179
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1649977179
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1649977179
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1649977179
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1649977179
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1649977179
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1649977179
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1649977179
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1649977179
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1649977179
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1649977179
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1649977179
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1649977179
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1649977179
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1649977179
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1649977179
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1649977179
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1649977179
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1649977179
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1649977179
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1649977179
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1649977179
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1649977179
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1649977179
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1649977179
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1649977179
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1649977179
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1649977179
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1649977179
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1649977179
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_501
timestamp 1649977179
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_513
timestamp 1649977179
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_525
timestamp 1649977179
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_531
timestamp 1649977179
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_533
timestamp 1649977179
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_545
timestamp 1649977179
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_557
timestamp 1649977179
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_569
timestamp 1649977179
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_581
timestamp 1649977179
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_587
timestamp 1649977179
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_589
timestamp 1649977179
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_601
timestamp 1649977179
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_613
timestamp 1649977179
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_625
timestamp 1649977179
transform 1 0 58604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_637
timestamp 1649977179
transform 1 0 59708 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_643
timestamp 1649977179
transform 1 0 60260 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_645
timestamp 1649977179
transform 1 0 60444 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_657
timestamp 1649977179
transform 1 0 61548 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_669
timestamp 1649977179
transform 1 0 62652 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_681
timestamp 1649977179
transform 1 0 63756 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_693
timestamp 1649977179
transform 1 0 64860 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_699
timestamp 1649977179
transform 1 0 65412 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_701
timestamp 1649977179
transform 1 0 65596 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_713
timestamp 1649977179
transform 1 0 66700 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_725
timestamp 1649977179
transform 1 0 67804 0 1 46784
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1649977179
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1649977179
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1649977179
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1649977179
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1649977179
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1649977179
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1649977179
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1649977179
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1649977179
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1649977179
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1649977179
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1649977179
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1649977179
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1649977179
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1649977179
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1649977179
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1649977179
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1649977179
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1649977179
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1649977179
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1649977179
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1649977179
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1649977179
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1649977179
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1649977179
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1649977179
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_249
timestamp 1649977179
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_261
timestamp 1649977179
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_273
timestamp 1649977179
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1649977179
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1649977179
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1649977179
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1649977179
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1649977179
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1649977179
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1649977179
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1649977179
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1649977179
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1649977179
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1649977179
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1649977179
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1649977179
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1649977179
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1649977179
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1649977179
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1649977179
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1649977179
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1649977179
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1649977179
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1649977179
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1649977179
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1649977179
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1649977179
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1649977179
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1649977179
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_517
timestamp 1649977179
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_529
timestamp 1649977179
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_541
timestamp 1649977179
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_553
timestamp 1649977179
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_559
timestamp 1649977179
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_561
timestamp 1649977179
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_573
timestamp 1649977179
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_585
timestamp 1649977179
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_597
timestamp 1649977179
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_609
timestamp 1649977179
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_615
timestamp 1649977179
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_617
timestamp 1649977179
transform 1 0 57868 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_629
timestamp 1649977179
transform 1 0 58972 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_641
timestamp 1649977179
transform 1 0 60076 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_653
timestamp 1649977179
transform 1 0 61180 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_665
timestamp 1649977179
transform 1 0 62284 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_671
timestamp 1649977179
transform 1 0 62836 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_673
timestamp 1649977179
transform 1 0 63020 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_685
timestamp 1649977179
transform 1 0 64124 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_697
timestamp 1649977179
transform 1 0 65228 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_709
timestamp 1649977179
transform 1 0 66332 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_721
timestamp 1649977179
transform 1 0 67436 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_727
timestamp 1649977179
transform 1 0 67988 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_729
timestamp 1649977179
transform 1 0 68172 0 -1 47872
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_84_3
timestamp 1649977179
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_15
timestamp 1649977179
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1649977179
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1649977179
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1649977179
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1649977179
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1649977179
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1649977179
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1649977179
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1649977179
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_97
timestamp 1649977179
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_109
timestamp 1649977179
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1649977179
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1649977179
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1649977179
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1649977179
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1649977179
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1649977179
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1649977179
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1649977179
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1649977179
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1649977179
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1649977179
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1649977179
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1649977179
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1649977179
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1649977179
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1649977179
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1649977179
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1649977179
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1649977179
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1649977179
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1649977179
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1649977179
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1649977179
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1649977179
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1649977179
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1649977179
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1649977179
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1649977179
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1649977179
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1649977179
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1649977179
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1649977179
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1649977179
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1649977179
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1649977179
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1649977179
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1649977179
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1649977179
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1649977179
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1649977179
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1649977179
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_501
timestamp 1649977179
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_513
timestamp 1649977179
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_525
timestamp 1649977179
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_531
timestamp 1649977179
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_533
timestamp 1649977179
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_545
timestamp 1649977179
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_557
timestamp 1649977179
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_569
timestamp 1649977179
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_581
timestamp 1649977179
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_587
timestamp 1649977179
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_589
timestamp 1649977179
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_601
timestamp 1649977179
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_613
timestamp 1649977179
transform 1 0 57500 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_625
timestamp 1649977179
transform 1 0 58604 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_637
timestamp 1649977179
transform 1 0 59708 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_643
timestamp 1649977179
transform 1 0 60260 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_645
timestamp 1649977179
transform 1 0 60444 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_657
timestamp 1649977179
transform 1 0 61548 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_669
timestamp 1649977179
transform 1 0 62652 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_681
timestamp 1649977179
transform 1 0 63756 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_693
timestamp 1649977179
transform 1 0 64860 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_699
timestamp 1649977179
transform 1 0 65412 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_701
timestamp 1649977179
transform 1 0 65596 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_713
timestamp 1649977179
transform 1 0 66700 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_725
timestamp 1649977179
transform 1 0 67804 0 1 47872
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1649977179
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1649977179
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1649977179
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1649977179
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1649977179
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1649977179
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1649977179
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1649977179
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1649977179
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1649977179
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1649977179
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1649977179
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1649977179
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1649977179
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1649977179
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1649977179
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1649977179
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1649977179
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1649977179
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1649977179
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1649977179
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1649977179
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1649977179
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1649977179
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1649977179
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1649977179
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1649977179
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1649977179
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1649977179
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1649977179
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1649977179
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1649977179
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1649977179
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1649977179
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1649977179
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1649977179
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1649977179
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1649977179
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1649977179
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1649977179
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1649977179
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1649977179
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1649977179
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1649977179
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1649977179
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1649977179
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1649977179
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1649977179
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1649977179
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1649977179
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1649977179
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1649977179
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1649977179
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1649977179
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1649977179
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_517
timestamp 1649977179
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_529
timestamp 1649977179
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_541
timestamp 1649977179
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_553
timestamp 1649977179
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_559
timestamp 1649977179
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_561
timestamp 1649977179
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_573
timestamp 1649977179
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_585
timestamp 1649977179
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_597
timestamp 1649977179
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_609
timestamp 1649977179
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_615
timestamp 1649977179
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_617
timestamp 1649977179
transform 1 0 57868 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_629
timestamp 1649977179
transform 1 0 58972 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_641
timestamp 1649977179
transform 1 0 60076 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_653
timestamp 1649977179
transform 1 0 61180 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_665
timestamp 1649977179
transform 1 0 62284 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_671
timestamp 1649977179
transform 1 0 62836 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_673
timestamp 1649977179
transform 1 0 63020 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_685
timestamp 1649977179
transform 1 0 64124 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_697
timestamp 1649977179
transform 1 0 65228 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_709
timestamp 1649977179
transform 1 0 66332 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_717
timestamp 1649977179
transform 1 0 67068 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_724
timestamp 1649977179
transform 1 0 67712 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_729
timestamp 1649977179
transform 1 0 68172 0 -1 48960
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1649977179
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1649977179
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1649977179
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1649977179
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1649977179
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1649977179
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1649977179
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1649977179
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1649977179
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1649977179
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1649977179
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1649977179
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1649977179
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1649977179
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1649977179
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1649977179
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1649977179
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1649977179
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_177
timestamp 1649977179
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_189
timestamp 1649977179
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_195
timestamp 1649977179
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_197
timestamp 1649977179
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_209
timestamp 1649977179
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_221
timestamp 1649977179
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_233
timestamp 1649977179
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_245
timestamp 1649977179
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1649977179
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1649977179
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1649977179
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1649977179
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1649977179
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1649977179
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1649977179
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1649977179
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1649977179
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1649977179
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1649977179
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1649977179
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1649977179
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1649977179
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1649977179
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1649977179
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1649977179
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1649977179
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1649977179
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1649977179
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1649977179
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1649977179
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1649977179
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1649977179
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1649977179
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1649977179
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1649977179
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1649977179
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_513
timestamp 1649977179
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_525
timestamp 1649977179
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_531
timestamp 1649977179
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_533
timestamp 1649977179
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_545
timestamp 1649977179
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_557
timestamp 1649977179
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_569
timestamp 1649977179
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_581
timestamp 1649977179
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_587
timestamp 1649977179
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_589
timestamp 1649977179
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_601
timestamp 1649977179
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_613
timestamp 1649977179
transform 1 0 57500 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_625
timestamp 1649977179
transform 1 0 58604 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_637
timestamp 1649977179
transform 1 0 59708 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_643
timestamp 1649977179
transform 1 0 60260 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_645
timestamp 1649977179
transform 1 0 60444 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_657
timestamp 1649977179
transform 1 0 61548 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_669
timestamp 1649977179
transform 1 0 62652 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_681
timestamp 1649977179
transform 1 0 63756 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_693
timestamp 1649977179
transform 1 0 64860 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_699
timestamp 1649977179
transform 1 0 65412 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_701
timestamp 1649977179
transform 1 0 65596 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_713
timestamp 1649977179
transform 1 0 66700 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_725
timestamp 1649977179
transform 1 0 67804 0 1 48960
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1649977179
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1649977179
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1649977179
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1649977179
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1649977179
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1649977179
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1649977179
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1649977179
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1649977179
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1649977179
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1649977179
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1649977179
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_113
timestamp 1649977179
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_125
timestamp 1649977179
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_137
timestamp 1649977179
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_149
timestamp 1649977179
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_161
timestamp 1649977179
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_167
timestamp 1649977179
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1649977179
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1649977179
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1649977179
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1649977179
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1649977179
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1649977179
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1649977179
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1649977179
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1649977179
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1649977179
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1649977179
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1649977179
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1649977179
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1649977179
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1649977179
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1649977179
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1649977179
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1649977179
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1649977179
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1649977179
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1649977179
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1649977179
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1649977179
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1649977179
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1649977179
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1649977179
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1649977179
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1649977179
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1649977179
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1649977179
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1649977179
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1649977179
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1649977179
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1649977179
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1649977179
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1649977179
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1649977179
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_517
timestamp 1649977179
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_529
timestamp 1649977179
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_541
timestamp 1649977179
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_553
timestamp 1649977179
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_559
timestamp 1649977179
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_561
timestamp 1649977179
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_573
timestamp 1649977179
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_585
timestamp 1649977179
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_597
timestamp 1649977179
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_609
timestamp 1649977179
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_615
timestamp 1649977179
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_617
timestamp 1649977179
transform 1 0 57868 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_629
timestamp 1649977179
transform 1 0 58972 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_641
timestamp 1649977179
transform 1 0 60076 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_653
timestamp 1649977179
transform 1 0 61180 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_665
timestamp 1649977179
transform 1 0 62284 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_671
timestamp 1649977179
transform 1 0 62836 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_673
timestamp 1649977179
transform 1 0 63020 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_685
timestamp 1649977179
transform 1 0 64124 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_697
timestamp 1649977179
transform 1 0 65228 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_709
timestamp 1649977179
transform 1 0 66332 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_721
timestamp 1649977179
transform 1 0 67436 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_727
timestamp 1649977179
transform 1 0 67988 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_87_729
timestamp 1649977179
transform 1 0 68172 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1649977179
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1649977179
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1649977179
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1649977179
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1649977179
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1649977179
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1649977179
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1649977179
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1649977179
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1649977179
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1649977179
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1649977179
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1649977179
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1649977179
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1649977179
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1649977179
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1649977179
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1649977179
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1649977179
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1649977179
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1649977179
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_197
timestamp 1649977179
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_209
timestamp 1649977179
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_221
timestamp 1649977179
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_233
timestamp 1649977179
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_245
timestamp 1649977179
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_251
timestamp 1649977179
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1649977179
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1649977179
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1649977179
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1649977179
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1649977179
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1649977179
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1649977179
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1649977179
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1649977179
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1649977179
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1649977179
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1649977179
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1649977179
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1649977179
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1649977179
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1649977179
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1649977179
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1649977179
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1649977179
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1649977179
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1649977179
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1649977179
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1649977179
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1649977179
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1649977179
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1649977179
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1649977179
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_513
timestamp 1649977179
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_525
timestamp 1649977179
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_531
timestamp 1649977179
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_533
timestamp 1649977179
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_545
timestamp 1649977179
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_557
timestamp 1649977179
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_569
timestamp 1649977179
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_581
timestamp 1649977179
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_587
timestamp 1649977179
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_589
timestamp 1649977179
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_601
timestamp 1649977179
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_613
timestamp 1649977179
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_625
timestamp 1649977179
transform 1 0 58604 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_637
timestamp 1649977179
transform 1 0 59708 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_643
timestamp 1649977179
transform 1 0 60260 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_645
timestamp 1649977179
transform 1 0 60444 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_657
timestamp 1649977179
transform 1 0 61548 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_669
timestamp 1649977179
transform 1 0 62652 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_681
timestamp 1649977179
transform 1 0 63756 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_693
timestamp 1649977179
transform 1 0 64860 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_699
timestamp 1649977179
transform 1 0 65412 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_701
timestamp 1649977179
transform 1 0 65596 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_713
timestamp 1649977179
transform 1 0 66700 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_725
timestamp 1649977179
transform 1 0 67804 0 1 50048
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_89_3
timestamp 1649977179
transform 1 0 1380 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_15
timestamp 1649977179
transform 1 0 2484 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_27
timestamp 1649977179
transform 1 0 3588 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_39
timestamp 1649977179
transform 1 0 4692 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_51
timestamp 1649977179
transform 1 0 5796 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_89_55
timestamp 1649977179
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1649977179
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1649977179
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1649977179
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1649977179
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1649977179
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1649977179
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1649977179
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1649977179
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1649977179
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1649977179
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1649977179
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1649977179
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1649977179
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1649977179
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1649977179
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1649977179
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1649977179
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1649977179
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_225
timestamp 1649977179
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_237
timestamp 1649977179
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_249
timestamp 1649977179
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_261
timestamp 1649977179
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_273
timestamp 1649977179
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_279
timestamp 1649977179
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1649977179
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1649977179
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1649977179
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1649977179
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1649977179
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1649977179
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1649977179
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1649977179
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1649977179
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1649977179
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1649977179
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1649977179
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1649977179
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1649977179
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1649977179
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1649977179
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1649977179
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1649977179
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1649977179
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1649977179
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1649977179
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1649977179
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1649977179
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1649977179
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1649977179
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_517
timestamp 1649977179
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_529
timestamp 1649977179
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_541
timestamp 1649977179
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_553
timestamp 1649977179
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_559
timestamp 1649977179
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_561
timestamp 1649977179
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_573
timestamp 1649977179
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_585
timestamp 1649977179
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_597
timestamp 1649977179
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_609
timestamp 1649977179
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_615
timestamp 1649977179
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_617
timestamp 1649977179
transform 1 0 57868 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_629
timestamp 1649977179
transform 1 0 58972 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_641
timestamp 1649977179
transform 1 0 60076 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_653
timestamp 1649977179
transform 1 0 61180 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_665
timestamp 1649977179
transform 1 0 62284 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_671
timestamp 1649977179
transform 1 0 62836 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_673
timestamp 1649977179
transform 1 0 63020 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_685
timestamp 1649977179
transform 1 0 64124 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_697
timestamp 1649977179
transform 1 0 65228 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_709
timestamp 1649977179
transform 1 0 66332 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_721
timestamp 1649977179
transform 1 0 67436 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_727
timestamp 1649977179
transform 1 0 67988 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_729
timestamp 1649977179
transform 1 0 68172 0 -1 51136
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1649977179
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1649977179
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1649977179
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1649977179
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1649977179
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1649977179
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1649977179
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1649977179
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1649977179
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1649977179
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1649977179
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1649977179
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_121
timestamp 1649977179
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_133
timestamp 1649977179
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_139
timestamp 1649977179
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_141
timestamp 1649977179
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_153
timestamp 1649977179
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_165
timestamp 1649977179
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_177
timestamp 1649977179
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_189
timestamp 1649977179
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1649977179
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1649977179
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1649977179
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1649977179
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1649977179
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1649977179
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1649977179
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_253
timestamp 1649977179
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_265
timestamp 1649977179
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_277
timestamp 1649977179
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_289
timestamp 1649977179
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_301
timestamp 1649977179
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1649977179
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1649977179
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1649977179
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1649977179
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1649977179
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1649977179
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1649977179
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1649977179
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1649977179
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1649977179
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1649977179
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1649977179
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1649977179
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1649977179
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1649977179
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1649977179
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1649977179
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1649977179
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1649977179
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1649977179
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1649977179
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1649977179
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_513
timestamp 1649977179
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_525
timestamp 1649977179
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_531
timestamp 1649977179
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_533
timestamp 1649977179
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_545
timestamp 1649977179
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_557
timestamp 1649977179
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_569
timestamp 1649977179
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_581
timestamp 1649977179
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_587
timestamp 1649977179
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_589
timestamp 1649977179
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_601
timestamp 1649977179
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_613
timestamp 1649977179
transform 1 0 57500 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_625
timestamp 1649977179
transform 1 0 58604 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_637
timestamp 1649977179
transform 1 0 59708 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_643
timestamp 1649977179
transform 1 0 60260 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_645
timestamp 1649977179
transform 1 0 60444 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_657
timestamp 1649977179
transform 1 0 61548 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_669
timestamp 1649977179
transform 1 0 62652 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_681
timestamp 1649977179
transform 1 0 63756 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_693
timestamp 1649977179
transform 1 0 64860 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_699
timestamp 1649977179
transform 1 0 65412 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_701
timestamp 1649977179
transform 1 0 65596 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_713
timestamp 1649977179
transform 1 0 66700 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_725
timestamp 1649977179
transform 1 0 67804 0 1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_91_3
timestamp 1649977179
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_15
timestamp 1649977179
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_27
timestamp 1649977179
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_39
timestamp 1649977179
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_51
timestamp 1649977179
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_55
timestamp 1649977179
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1649977179
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1649977179
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1649977179
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1649977179
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1649977179
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1649977179
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1649977179
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1649977179
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1649977179
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1649977179
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1649977179
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1649977179
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1649977179
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1649977179
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1649977179
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1649977179
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1649977179
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1649977179
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1649977179
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_237
timestamp 1649977179
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_249
timestamp 1649977179
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_261
timestamp 1649977179
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_273
timestamp 1649977179
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1649977179
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1649977179
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1649977179
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1649977179
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1649977179
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1649977179
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1649977179
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1649977179
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1649977179
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1649977179
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1649977179
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1649977179
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1649977179
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1649977179
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1649977179
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1649977179
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1649977179
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1649977179
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1649977179
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1649977179
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1649977179
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1649977179
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1649977179
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1649977179
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1649977179
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1649977179
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_517
timestamp 1649977179
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_529
timestamp 1649977179
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_541
timestamp 1649977179
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_553
timestamp 1649977179
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_559
timestamp 1649977179
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_561
timestamp 1649977179
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_573
timestamp 1649977179
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_585
timestamp 1649977179
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_597
timestamp 1649977179
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_609
timestamp 1649977179
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_615
timestamp 1649977179
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_617
timestamp 1649977179
transform 1 0 57868 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_629
timestamp 1649977179
transform 1 0 58972 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_641
timestamp 1649977179
transform 1 0 60076 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_653
timestamp 1649977179
transform 1 0 61180 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_665
timestamp 1649977179
transform 1 0 62284 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_671
timestamp 1649977179
transform 1 0 62836 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_673
timestamp 1649977179
transform 1 0 63020 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_685
timestamp 1649977179
transform 1 0 64124 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_697
timestamp 1649977179
transform 1 0 65228 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_709
timestamp 1649977179
transform 1 0 66332 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_721
timestamp 1649977179
transform 1 0 67436 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_727
timestamp 1649977179
transform 1 0 67988 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_729
timestamp 1649977179
transform 1 0 68172 0 -1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_3
timestamp 1649977179
transform 1 0 1380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_15
timestamp 1649977179
transform 1 0 2484 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1649977179
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_29
timestamp 1649977179
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_41
timestamp 1649977179
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_53
timestamp 1649977179
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_65
timestamp 1649977179
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_77
timestamp 1649977179
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_83
timestamp 1649977179
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_85
timestamp 1649977179
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_97
timestamp 1649977179
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_109
timestamp 1649977179
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_121
timestamp 1649977179
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_133
timestamp 1649977179
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_139
timestamp 1649977179
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_141
timestamp 1649977179
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_153
timestamp 1649977179
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_165
timestamp 1649977179
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_177
timestamp 1649977179
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_189
timestamp 1649977179
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_195
timestamp 1649977179
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1649977179
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1649977179
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1649977179
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1649977179
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1649977179
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1649977179
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1649977179
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1649977179
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1649977179
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1649977179
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1649977179
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1649977179
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1649977179
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1649977179
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1649977179
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1649977179
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1649977179
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1649977179
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1649977179
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1649977179
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1649977179
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1649977179
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1649977179
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1649977179
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1649977179
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1649977179
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1649977179
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1649977179
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1649977179
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1649977179
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1649977179
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1649977179
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1649977179
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_513
timestamp 1649977179
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_525
timestamp 1649977179
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_531
timestamp 1649977179
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_533
timestamp 1649977179
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_545
timestamp 1649977179
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_557
timestamp 1649977179
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_569
timestamp 1649977179
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_581
timestamp 1649977179
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_587
timestamp 1649977179
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_589
timestamp 1649977179
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_601
timestamp 1649977179
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_613
timestamp 1649977179
transform 1 0 57500 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_625
timestamp 1649977179
transform 1 0 58604 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_637
timestamp 1649977179
transform 1 0 59708 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_643
timestamp 1649977179
transform 1 0 60260 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_645
timestamp 1649977179
transform 1 0 60444 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_657
timestamp 1649977179
transform 1 0 61548 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_669
timestamp 1649977179
transform 1 0 62652 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_681
timestamp 1649977179
transform 1 0 63756 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_693
timestamp 1649977179
transform 1 0 64860 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_699
timestamp 1649977179
transform 1 0 65412 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_701
timestamp 1649977179
transform 1 0 65596 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_713
timestamp 1649977179
transform 1 0 66700 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_725
timestamp 1649977179
transform 1 0 67804 0 1 52224
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_93_3
timestamp 1649977179
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_15
timestamp 1649977179
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_27
timestamp 1649977179
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_39
timestamp 1649977179
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_51
timestamp 1649977179
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_55
timestamp 1649977179
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1649977179
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_69
timestamp 1649977179
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_81
timestamp 1649977179
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_93
timestamp 1649977179
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_105
timestamp 1649977179
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_111
timestamp 1649977179
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1649977179
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_125
timestamp 1649977179
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_137
timestamp 1649977179
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_149
timestamp 1649977179
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_161
timestamp 1649977179
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_167
timestamp 1649977179
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_169
timestamp 1649977179
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_181
timestamp 1649977179
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_193
timestamp 1649977179
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_205
timestamp 1649977179
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1649977179
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1649977179
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1649977179
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1649977179
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1649977179
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1649977179
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1649977179
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1649977179
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1649977179
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1649977179
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1649977179
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1649977179
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1649977179
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1649977179
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1649977179
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1649977179
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1649977179
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1649977179
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1649977179
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1649977179
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1649977179
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1649977179
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1649977179
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1649977179
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1649977179
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1649977179
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1649977179
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1649977179
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1649977179
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_485
timestamp 1649977179
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_497
timestamp 1649977179
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_503
timestamp 1649977179
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_505
timestamp 1649977179
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_517
timestamp 1649977179
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_529
timestamp 1649977179
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_541
timestamp 1649977179
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_553
timestamp 1649977179
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_559
timestamp 1649977179
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_561
timestamp 1649977179
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_573
timestamp 1649977179
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_585
timestamp 1649977179
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_597
timestamp 1649977179
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_609
timestamp 1649977179
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_615
timestamp 1649977179
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_617
timestamp 1649977179
transform 1 0 57868 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_629
timestamp 1649977179
transform 1 0 58972 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_641
timestamp 1649977179
transform 1 0 60076 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_653
timestamp 1649977179
transform 1 0 61180 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_665
timestamp 1649977179
transform 1 0 62284 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_671
timestamp 1649977179
transform 1 0 62836 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_673
timestamp 1649977179
transform 1 0 63020 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_685
timestamp 1649977179
transform 1 0 64124 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_697
timestamp 1649977179
transform 1 0 65228 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_709
timestamp 1649977179
transform 1 0 66332 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_721
timestamp 1649977179
transform 1 0 67436 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_727
timestamp 1649977179
transform 1 0 67988 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_729
timestamp 1649977179
transform 1 0 68172 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_3
timestamp 1649977179
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_15
timestamp 1649977179
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_27
timestamp 1649977179
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1649977179
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_41
timestamp 1649977179
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_53
timestamp 1649977179
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_65
timestamp 1649977179
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_77
timestamp 1649977179
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_83
timestamp 1649977179
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1649977179
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_97
timestamp 1649977179
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_109
timestamp 1649977179
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_121
timestamp 1649977179
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_133
timestamp 1649977179
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_139
timestamp 1649977179
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1649977179
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_153
timestamp 1649977179
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_165
timestamp 1649977179
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_177
timestamp 1649977179
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_189
timestamp 1649977179
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_195
timestamp 1649977179
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_197
timestamp 1649977179
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_209
timestamp 1649977179
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_221
timestamp 1649977179
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_233
timestamp 1649977179
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_245
timestamp 1649977179
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_251
timestamp 1649977179
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_253
timestamp 1649977179
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_265
timestamp 1649977179
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_277
timestamp 1649977179
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_289
timestamp 1649977179
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_301
timestamp 1649977179
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1649977179
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_309
timestamp 1649977179
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_321
timestamp 1649977179
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_333
timestamp 1649977179
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_345
timestamp 1649977179
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_357
timestamp 1649977179
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_363
timestamp 1649977179
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_365
timestamp 1649977179
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_377
timestamp 1649977179
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_389
timestamp 1649977179
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_401
timestamp 1649977179
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_413
timestamp 1649977179
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_419
timestamp 1649977179
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1649977179
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_433
timestamp 1649977179
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_445
timestamp 1649977179
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_457
timestamp 1649977179
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_469
timestamp 1649977179
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_475
timestamp 1649977179
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1649977179
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_489
timestamp 1649977179
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_501
timestamp 1649977179
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_513
timestamp 1649977179
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_525
timestamp 1649977179
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_531
timestamp 1649977179
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_533
timestamp 1649977179
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_545
timestamp 1649977179
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_557
timestamp 1649977179
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_569
timestamp 1649977179
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_581
timestamp 1649977179
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_587
timestamp 1649977179
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_589
timestamp 1649977179
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_601
timestamp 1649977179
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_613
timestamp 1649977179
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_625
timestamp 1649977179
transform 1 0 58604 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_637
timestamp 1649977179
transform 1 0 59708 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_643
timestamp 1649977179
transform 1 0 60260 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_645
timestamp 1649977179
transform 1 0 60444 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_657
timestamp 1649977179
transform 1 0 61548 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_669
timestamp 1649977179
transform 1 0 62652 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_681
timestamp 1649977179
transform 1 0 63756 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_94_693
timestamp 1649977179
transform 1 0 64860 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_94_699
timestamp 1649977179
transform 1 0 65412 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_701
timestamp 1649977179
transform 1 0 65596 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_713
timestamp 1649977179
transform 1 0 66700 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_725
timestamp 1649977179
transform 1 0 67804 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_95_3
timestamp 1649977179
transform 1 0 1380 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_15
timestamp 1649977179
transform 1 0 2484 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_27
timestamp 1649977179
transform 1 0 3588 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_39
timestamp 1649977179
transform 1 0 4692 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_51
timestamp 1649977179
transform 1 0 5796 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_55
timestamp 1649977179
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_57
timestamp 1649977179
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_69
timestamp 1649977179
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_81
timestamp 1649977179
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_93
timestamp 1649977179
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_105
timestamp 1649977179
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_111
timestamp 1649977179
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_113
timestamp 1649977179
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_125
timestamp 1649977179
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_137
timestamp 1649977179
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_149
timestamp 1649977179
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_161
timestamp 1649977179
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_167
timestamp 1649977179
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_169
timestamp 1649977179
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_181
timestamp 1649977179
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_193
timestamp 1649977179
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_205
timestamp 1649977179
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_217
timestamp 1649977179
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_223
timestamp 1649977179
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_225
timestamp 1649977179
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_237
timestamp 1649977179
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_249
timestamp 1649977179
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_261
timestamp 1649977179
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_273
timestamp 1649977179
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_279
timestamp 1649977179
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_281
timestamp 1649977179
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_293
timestamp 1649977179
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_305
timestamp 1649977179
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_317
timestamp 1649977179
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_329
timestamp 1649977179
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_335
timestamp 1649977179
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_337
timestamp 1649977179
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_349
timestamp 1649977179
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_361
timestamp 1649977179
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_373
timestamp 1649977179
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_385
timestamp 1649977179
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_391
timestamp 1649977179
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_393
timestamp 1649977179
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_405
timestamp 1649977179
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_417
timestamp 1649977179
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_429
timestamp 1649977179
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_441
timestamp 1649977179
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_447
timestamp 1649977179
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_449
timestamp 1649977179
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_461
timestamp 1649977179
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_473
timestamp 1649977179
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_485
timestamp 1649977179
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_497
timestamp 1649977179
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_503
timestamp 1649977179
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_505
timestamp 1649977179
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_517
timestamp 1649977179
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_529
timestamp 1649977179
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_541
timestamp 1649977179
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_553
timestamp 1649977179
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_559
timestamp 1649977179
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_561
timestamp 1649977179
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_573
timestamp 1649977179
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_585
timestamp 1649977179
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_597
timestamp 1649977179
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_609
timestamp 1649977179
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_615
timestamp 1649977179
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_617
timestamp 1649977179
transform 1 0 57868 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_629
timestamp 1649977179
transform 1 0 58972 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_641
timestamp 1649977179
transform 1 0 60076 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_653
timestamp 1649977179
transform 1 0 61180 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_665
timestamp 1649977179
transform 1 0 62284 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_671
timestamp 1649977179
transform 1 0 62836 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_95_673
timestamp 1649977179
transform 1 0 63020 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_685
timestamp 1649977179
transform 1 0 64124 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_697
timestamp 1649977179
transform 1 0 65228 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_95_709
timestamp 1649977179
transform 1 0 66332 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_95_721
timestamp 1649977179
transform 1 0 67436 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_727
timestamp 1649977179
transform 1 0 67988 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_729
timestamp 1649977179
transform 1 0 68172 0 -1 54400
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_96_3
timestamp 1649977179
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_15
timestamp 1649977179
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_27
timestamp 1649977179
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_29
timestamp 1649977179
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_41
timestamp 1649977179
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_53
timestamp 1649977179
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_65
timestamp 1649977179
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_77
timestamp 1649977179
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_83
timestamp 1649977179
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_85
timestamp 1649977179
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_97
timestamp 1649977179
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_109
timestamp 1649977179
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_121
timestamp 1649977179
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_133
timestamp 1649977179
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_139
timestamp 1649977179
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_141
timestamp 1649977179
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_153
timestamp 1649977179
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_165
timestamp 1649977179
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_177
timestamp 1649977179
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_189
timestamp 1649977179
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_195
timestamp 1649977179
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_197
timestamp 1649977179
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_209
timestamp 1649977179
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_221
timestamp 1649977179
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_233
timestamp 1649977179
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_245
timestamp 1649977179
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_251
timestamp 1649977179
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_253
timestamp 1649977179
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_265
timestamp 1649977179
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_277
timestamp 1649977179
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_289
timestamp 1649977179
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_301
timestamp 1649977179
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_307
timestamp 1649977179
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_309
timestamp 1649977179
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_321
timestamp 1649977179
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_333
timestamp 1649977179
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_345
timestamp 1649977179
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_357
timestamp 1649977179
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_363
timestamp 1649977179
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_365
timestamp 1649977179
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_377
timestamp 1649977179
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_389
timestamp 1649977179
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_401
timestamp 1649977179
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_413
timestamp 1649977179
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_419
timestamp 1649977179
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_421
timestamp 1649977179
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_433
timestamp 1649977179
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_445
timestamp 1649977179
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_457
timestamp 1649977179
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_469
timestamp 1649977179
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_475
timestamp 1649977179
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_477
timestamp 1649977179
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_489
timestamp 1649977179
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_501
timestamp 1649977179
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_513
timestamp 1649977179
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_525
timestamp 1649977179
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_531
timestamp 1649977179
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_533
timestamp 1649977179
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_545
timestamp 1649977179
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_557
timestamp 1649977179
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_569
timestamp 1649977179
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_581
timestamp 1649977179
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_587
timestamp 1649977179
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_589
timestamp 1649977179
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_601
timestamp 1649977179
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_613
timestamp 1649977179
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_625
timestamp 1649977179
transform 1 0 58604 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_637
timestamp 1649977179
transform 1 0 59708 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_643
timestamp 1649977179
transform 1 0 60260 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_645
timestamp 1649977179
transform 1 0 60444 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_657
timestamp 1649977179
transform 1 0 61548 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_669
timestamp 1649977179
transform 1 0 62652 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_681
timestamp 1649977179
transform 1 0 63756 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_693
timestamp 1649977179
transform 1 0 64860 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_96_699
timestamp 1649977179
transform 1 0 65412 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_96_701
timestamp 1649977179
transform 1 0 65596 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_96_713
timestamp 1649977179
transform 1 0 66700 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_725
timestamp 1649977179
transform 1 0 67804 0 1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_97_3
timestamp 1649977179
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_15
timestamp 1649977179
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_27
timestamp 1649977179
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_39
timestamp 1649977179
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_51
timestamp 1649977179
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_97_55
timestamp 1649977179
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_57
timestamp 1649977179
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_69
timestamp 1649977179
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_81
timestamp 1649977179
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_93
timestamp 1649977179
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_105
timestamp 1649977179
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_111
timestamp 1649977179
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_113
timestamp 1649977179
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_125
timestamp 1649977179
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_137
timestamp 1649977179
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_149
timestamp 1649977179
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_161
timestamp 1649977179
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_167
timestamp 1649977179
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_169
timestamp 1649977179
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_181
timestamp 1649977179
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_193
timestamp 1649977179
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_205
timestamp 1649977179
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_217
timestamp 1649977179
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_223
timestamp 1649977179
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_225
timestamp 1649977179
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_237
timestamp 1649977179
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_249
timestamp 1649977179
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_261
timestamp 1649977179
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_273
timestamp 1649977179
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_279
timestamp 1649977179
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_281
timestamp 1649977179
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_293
timestamp 1649977179
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_305
timestamp 1649977179
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_317
timestamp 1649977179
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_329
timestamp 1649977179
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_335
timestamp 1649977179
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_337
timestamp 1649977179
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_349
timestamp 1649977179
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_361
timestamp 1649977179
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_373
timestamp 1649977179
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_385
timestamp 1649977179
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_391
timestamp 1649977179
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_393
timestamp 1649977179
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_405
timestamp 1649977179
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_417
timestamp 1649977179
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_429
timestamp 1649977179
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_441
timestamp 1649977179
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_447
timestamp 1649977179
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_449
timestamp 1649977179
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_461
timestamp 1649977179
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_473
timestamp 1649977179
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_485
timestamp 1649977179
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_497
timestamp 1649977179
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_503
timestamp 1649977179
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_505
timestamp 1649977179
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_517
timestamp 1649977179
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_529
timestamp 1649977179
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_541
timestamp 1649977179
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_553
timestamp 1649977179
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_559
timestamp 1649977179
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_561
timestamp 1649977179
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_573
timestamp 1649977179
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_585
timestamp 1649977179
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_597
timestamp 1649977179
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_609
timestamp 1649977179
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_615
timestamp 1649977179
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_617
timestamp 1649977179
transform 1 0 57868 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_629
timestamp 1649977179
transform 1 0 58972 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_641
timestamp 1649977179
transform 1 0 60076 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_653
timestamp 1649977179
transform 1 0 61180 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_665
timestamp 1649977179
transform 1 0 62284 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_671
timestamp 1649977179
transform 1 0 62836 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_97_673
timestamp 1649977179
transform 1 0 63020 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_685
timestamp 1649977179
transform 1 0 64124 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_697
timestamp 1649977179
transform 1 0 65228 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_97_709
timestamp 1649977179
transform 1 0 66332 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_97_721
timestamp 1649977179
transform 1 0 67436 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_97_727
timestamp 1649977179
transform 1 0 67988 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_97_729
timestamp 1649977179
transform 1 0 68172 0 -1 55488
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_98_3
timestamp 1649977179
transform 1 0 1380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_15
timestamp 1649977179
transform 1 0 2484 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_27
timestamp 1649977179
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_29
timestamp 1649977179
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_41
timestamp 1649977179
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_53
timestamp 1649977179
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_65
timestamp 1649977179
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_77
timestamp 1649977179
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_83
timestamp 1649977179
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_85
timestamp 1649977179
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_97
timestamp 1649977179
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_109
timestamp 1649977179
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_121
timestamp 1649977179
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_133
timestamp 1649977179
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_139
timestamp 1649977179
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_141
timestamp 1649977179
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_153
timestamp 1649977179
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_165
timestamp 1649977179
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_177
timestamp 1649977179
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_189
timestamp 1649977179
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_195
timestamp 1649977179
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_197
timestamp 1649977179
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_209
timestamp 1649977179
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_221
timestamp 1649977179
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_233
timestamp 1649977179
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_245
timestamp 1649977179
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_251
timestamp 1649977179
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_253
timestamp 1649977179
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_265
timestamp 1649977179
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_277
timestamp 1649977179
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_289
timestamp 1649977179
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_301
timestamp 1649977179
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_307
timestamp 1649977179
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_309
timestamp 1649977179
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_321
timestamp 1649977179
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_333
timestamp 1649977179
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_345
timestamp 1649977179
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_357
timestamp 1649977179
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_363
timestamp 1649977179
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_365
timestamp 1649977179
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_377
timestamp 1649977179
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_389
timestamp 1649977179
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_401
timestamp 1649977179
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_413
timestamp 1649977179
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_419
timestamp 1649977179
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_421
timestamp 1649977179
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_433
timestamp 1649977179
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_445
timestamp 1649977179
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_457
timestamp 1649977179
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_469
timestamp 1649977179
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_475
timestamp 1649977179
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_477
timestamp 1649977179
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_489
timestamp 1649977179
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_501
timestamp 1649977179
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_513
timestamp 1649977179
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_525
timestamp 1649977179
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_531
timestamp 1649977179
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_533
timestamp 1649977179
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_545
timestamp 1649977179
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_557
timestamp 1649977179
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_569
timestamp 1649977179
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_581
timestamp 1649977179
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_587
timestamp 1649977179
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_589
timestamp 1649977179
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_601
timestamp 1649977179
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_613
timestamp 1649977179
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_625
timestamp 1649977179
transform 1 0 58604 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_637
timestamp 1649977179
transform 1 0 59708 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_643
timestamp 1649977179
transform 1 0 60260 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_645
timestamp 1649977179
transform 1 0 60444 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_657
timestamp 1649977179
transform 1 0 61548 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_669
timestamp 1649977179
transform 1 0 62652 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_681
timestamp 1649977179
transform 1 0 63756 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_98_693
timestamp 1649977179
transform 1 0 64860 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_699
timestamp 1649977179
transform 1 0 65412 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_98_701
timestamp 1649977179
transform 1 0 65596 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_98_713
timestamp 1649977179
transform 1 0 66700 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_725
timestamp 1649977179
transform 1 0 67804 0 1 55488
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_99_3
timestamp 1649977179
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_15
timestamp 1649977179
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_27
timestamp 1649977179
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_39
timestamp 1649977179
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_51
timestamp 1649977179
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_99_55
timestamp 1649977179
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_57
timestamp 1649977179
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_69
timestamp 1649977179
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_81
timestamp 1649977179
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_93
timestamp 1649977179
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_105
timestamp 1649977179
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_111
timestamp 1649977179
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_113
timestamp 1649977179
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_125
timestamp 1649977179
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_137
timestamp 1649977179
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_149
timestamp 1649977179
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_161
timestamp 1649977179
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_167
timestamp 1649977179
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_169
timestamp 1649977179
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_181
timestamp 1649977179
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_193
timestamp 1649977179
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_205
timestamp 1649977179
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_217
timestamp 1649977179
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_223
timestamp 1649977179
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_225
timestamp 1649977179
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_237
timestamp 1649977179
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_249
timestamp 1649977179
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_261
timestamp 1649977179
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_273
timestamp 1649977179
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_279
timestamp 1649977179
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_281
timestamp 1649977179
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_293
timestamp 1649977179
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_305
timestamp 1649977179
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_317
timestamp 1649977179
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_329
timestamp 1649977179
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_335
timestamp 1649977179
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_337
timestamp 1649977179
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_349
timestamp 1649977179
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_361
timestamp 1649977179
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_373
timestamp 1649977179
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_385
timestamp 1649977179
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_391
timestamp 1649977179
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_393
timestamp 1649977179
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_405
timestamp 1649977179
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_417
timestamp 1649977179
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_429
timestamp 1649977179
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_441
timestamp 1649977179
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_447
timestamp 1649977179
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_449
timestamp 1649977179
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_461
timestamp 1649977179
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_473
timestamp 1649977179
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_485
timestamp 1649977179
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_497
timestamp 1649977179
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_503
timestamp 1649977179
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_505
timestamp 1649977179
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_517
timestamp 1649977179
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_529
timestamp 1649977179
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_541
timestamp 1649977179
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_553
timestamp 1649977179
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_559
timestamp 1649977179
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_561
timestamp 1649977179
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_573
timestamp 1649977179
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_585
timestamp 1649977179
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_597
timestamp 1649977179
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_609
timestamp 1649977179
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_615
timestamp 1649977179
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_617
timestamp 1649977179
transform 1 0 57868 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_629
timestamp 1649977179
transform 1 0 58972 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_641
timestamp 1649977179
transform 1 0 60076 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_653
timestamp 1649977179
transform 1 0 61180 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_99_665
timestamp 1649977179
transform 1 0 62284 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_99_671
timestamp 1649977179
transform 1 0 62836 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_99_673
timestamp 1649977179
transform 1 0 63020 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_685
timestamp 1649977179
transform 1 0 64124 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_99_697
timestamp 1649977179
transform 1 0 65228 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_99_709
timestamp 1649977179
transform 1 0 66332 0 -1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_99_717
timestamp 1649977179
transform 1 0 67068 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_99_724
timestamp 1649977179
transform 1 0 67712 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_99_729
timestamp 1649977179
transform 1 0 68172 0 -1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_3
timestamp 1649977179
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_15
timestamp 1649977179
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_27
timestamp 1649977179
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_29
timestamp 1649977179
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_41
timestamp 1649977179
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_53
timestamp 1649977179
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_65
timestamp 1649977179
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_77
timestamp 1649977179
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_83
timestamp 1649977179
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_85
timestamp 1649977179
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_97
timestamp 1649977179
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_109
timestamp 1649977179
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_121
timestamp 1649977179
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_133
timestamp 1649977179
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_139
timestamp 1649977179
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_141
timestamp 1649977179
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_153
timestamp 1649977179
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_165
timestamp 1649977179
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_177
timestamp 1649977179
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_189
timestamp 1649977179
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_195
timestamp 1649977179
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_197
timestamp 1649977179
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_209
timestamp 1649977179
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_221
timestamp 1649977179
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_233
timestamp 1649977179
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_245
timestamp 1649977179
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_251
timestamp 1649977179
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_256
timestamp 1649977179
transform 1 0 24656 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_268
timestamp 1649977179
transform 1 0 25760 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_280
timestamp 1649977179
transform 1 0 26864 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_292
timestamp 1649977179
transform 1 0 27968 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_304
timestamp 1649977179
transform 1 0 29072 0 1 56576
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_100_309
timestamp 1649977179
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_321
timestamp 1649977179
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_333
timestamp 1649977179
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_345
timestamp 1649977179
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_357
timestamp 1649977179
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_363
timestamp 1649977179
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_365
timestamp 1649977179
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_377
timestamp 1649977179
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_389
timestamp 1649977179
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_401
timestamp 1649977179
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_413
timestamp 1649977179
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_419
timestamp 1649977179
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_421
timestamp 1649977179
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_433
timestamp 1649977179
transform 1 0 40940 0 1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_100_437
timestamp 1649977179
transform 1 0 41308 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_441
timestamp 1649977179
transform 1 0 41676 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_453
timestamp 1649977179
transform 1 0 42780 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_465
timestamp 1649977179
transform 1 0 43884 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_100_473
timestamp 1649977179
transform 1 0 44620 0 1 56576
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_100_477
timestamp 1649977179
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_489
timestamp 1649977179
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_501
timestamp 1649977179
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_513
timestamp 1649977179
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_525
timestamp 1649977179
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_531
timestamp 1649977179
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_533
timestamp 1649977179
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_545
timestamp 1649977179
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_557
timestamp 1649977179
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_569
timestamp 1649977179
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_581
timestamp 1649977179
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_587
timestamp 1649977179
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_589
timestamp 1649977179
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_601
timestamp 1649977179
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_613
timestamp 1649977179
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_625
timestamp 1649977179
transform 1 0 58604 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_637
timestamp 1649977179
transform 1 0 59708 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_643
timestamp 1649977179
transform 1 0 60260 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_645
timestamp 1649977179
transform 1 0 60444 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_657
timestamp 1649977179
transform 1 0 61548 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_669
timestamp 1649977179
transform 1 0 62652 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_681
timestamp 1649977179
transform 1 0 63756 0 1 56576
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_689
timestamp 1649977179
transform 1 0 64492 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_693
timestamp 1649977179
transform 1 0 64860 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_699
timestamp 1649977179
transform 1 0 65412 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_100_701
timestamp 1649977179
transform 1 0 65596 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_100_713
timestamp 1649977179
transform 1 0 66700 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_725
timestamp 1649977179
transform 1 0 67804 0 1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_101_3
timestamp 1649977179
transform 1 0 1380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_101_15
timestamp 1649977179
transform 1 0 2484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_101_27
timestamp 1649977179
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_29
timestamp 1649977179
transform 1 0 3772 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_38
timestamp 1649977179
transform 1 0 4600 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_45
timestamp 1649977179
transform 1 0 5244 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_52
timestamp 1649977179
transform 1 0 5888 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_101_57
timestamp 1649977179
transform 1 0 6348 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_63
timestamp 1649977179
transform 1 0 6900 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_69
timestamp 1649977179
transform 1 0 7452 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_73
timestamp 1649977179
transform 1 0 7820 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_80
timestamp 1649977179
transform 1 0 8464 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_85
timestamp 1649977179
transform 1 0 8924 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_92
timestamp 1649977179
transform 1 0 9568 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_99
timestamp 1649977179
transform 1 0 10212 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_108
timestamp 1649977179
transform 1 0 11040 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_113
timestamp 1649977179
transform 1 0 11500 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_117
timestamp 1649977179
transform 1 0 11868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_128
timestamp 1649977179
transform 1 0 12880 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_135
timestamp 1649977179
transform 1 0 13524 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_139
timestamp 1649977179
transform 1 0 13892 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_141
timestamp 1649977179
transform 1 0 14076 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_146
timestamp 1649977179
transform 1 0 14536 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_153
timestamp 1649977179
transform 1 0 15180 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_164
timestamp 1649977179
transform 1 0 16192 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_172
timestamp 1649977179
transform 1 0 16928 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_178
timestamp 1649977179
transform 1 0 17480 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_182
timestamp 1649977179
transform 1 0 17848 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_189
timestamp 1649977179
transform 1 0 18492 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_195
timestamp 1649977179
transform 1 0 19044 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_200
timestamp 1649977179
transform 1 0 19504 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_207
timestamp 1649977179
transform 1 0 20148 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_215
timestamp 1649977179
transform 1 0 20884 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_219
timestamp 1649977179
transform 1 0 21252 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_223
timestamp 1649977179
transform 1 0 21620 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_228
timestamp 1649977179
transform 1 0 22080 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_232
timestamp 1649977179
transform 1 0 22448 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_236
timestamp 1649977179
transform 1 0 22816 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_243
timestamp 1649977179
transform 1 0 23460 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_251
timestamp 1649977179
transform 1 0 24196 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_253
timestamp 1649977179
transform 1 0 24380 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_257
timestamp 1649977179
transform 1 0 24748 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_261
timestamp 1649977179
transform 1 0 25116 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_265
timestamp 1649977179
transform 1 0 25484 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_269
timestamp 1649977179
transform 1 0 25852 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_276
timestamp 1649977179
transform 1 0 26496 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_281
timestamp 1649977179
transform 1 0 26956 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_290
timestamp 1649977179
transform 1 0 27784 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_297
timestamp 1649977179
transform 1 0 28428 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_304
timestamp 1649977179
transform 1 0 29072 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_101_309
timestamp 1649977179
transform 1 0 29532 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_101_315
timestamp 1649977179
transform 1 0 30084 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_321
timestamp 1649977179
transform 1 0 30636 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_325
timestamp 1649977179
transform 1 0 31004 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_332
timestamp 1649977179
transform 1 0 31648 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_337
timestamp 1649977179
transform 1 0 32108 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_344
timestamp 1649977179
transform 1 0 32752 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_351
timestamp 1649977179
transform 1 0 33396 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_360
timestamp 1649977179
transform 1 0 34224 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_365
timestamp 1649977179
transform 1 0 34684 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_369
timestamp 1649977179
transform 1 0 35052 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_377
timestamp 1649977179
transform 1 0 35788 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_381
timestamp 1649977179
transform 1 0 36156 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_388
timestamp 1649977179
transform 1 0 36800 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_101_393
timestamp 1649977179
transform 1 0 37260 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_101_399
timestamp 1649977179
transform 1 0 37812 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_406
timestamp 1649977179
transform 1 0 38456 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_101_418
timestamp 1649977179
transform 1 0 39560 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_424
timestamp 1649977179
transform 1 0 40112 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_431
timestamp 1649977179
transform 1 0 40756 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_438
timestamp 1649977179
transform 1 0 41400 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_446
timestamp 1649977179
transform 1 0 42136 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_449
timestamp 1649977179
transform 1 0 42412 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_453
timestamp 1649977179
transform 1 0 42780 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_460
timestamp 1649977179
transform 1 0 43424 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_471
timestamp 1649977179
transform 1 0 44436 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_475
timestamp 1649977179
transform 1 0 44804 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_480
timestamp 1649977179
transform 1 0 45264 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_101_489
timestamp 1649977179
transform 1 0 46092 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_496
timestamp 1649977179
transform 1 0 46736 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_101_508
timestamp 1649977179
transform 1 0 47840 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_101_515
timestamp 1649977179
transform 1 0 48484 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_521
timestamp 1649977179
transform 1 0 49036 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_525
timestamp 1649977179
transform 1 0 49404 0 -1 57664
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_101_531
timestamp 1649977179
transform 1 0 49956 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_536
timestamp 1649977179
transform 1 0 50416 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_543
timestamp 1649977179
transform 1 0 51060 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_550
timestamp 1649977179
transform 1 0 51704 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_558
timestamp 1649977179
transform 1 0 52440 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_564
timestamp 1649977179
transform 1 0 52992 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_571
timestamp 1649977179
transform 1 0 53636 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_575
timestamp 1649977179
transform 1 0 54004 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_579
timestamp 1649977179
transform 1 0 54372 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_101_587
timestamp 1649977179
transform 1 0 55108 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_592
timestamp 1649977179
transform 1 0 55568 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_599
timestamp 1649977179
transform 1 0 56212 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_606
timestamp 1649977179
transform 1 0 56856 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_614
timestamp 1649977179
transform 1 0 57592 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_620
timestamp 1649977179
transform 1 0 58144 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_627
timestamp 1649977179
transform 1 0 58788 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_634
timestamp 1649977179
transform 1 0 59432 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_642
timestamp 1649977179
transform 1 0 60168 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_648
timestamp 1649977179
transform 1 0 60720 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_655
timestamp 1649977179
transform 1 0 61364 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_662
timestamp 1649977179
transform 1 0 62008 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_670
timestamp 1649977179
transform 1 0 62744 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_676
timestamp 1649977179
transform 1 0 63296 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_683
timestamp 1649977179
transform 1 0 63940 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_101_690
timestamp 1649977179
transform 1 0 64584 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_698
timestamp 1649977179
transform 1 0 65320 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_701
timestamp 1649977179
transform 1 0 65596 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_101_705
timestamp 1649977179
transform 1 0 65964 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_101_712
timestamp 1649977179
transform 1 0 66608 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_724
timestamp 1649977179
transform 1 0 67712 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_101_729
timestamp 1649977179
transform 1 0 68172 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 68816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 68816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 68816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 68816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 68816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 68816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 68816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 68816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 68816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 68816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 68816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 68816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 68816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 68816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 68816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 68816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 68816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 68816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 68816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 68816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 68816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 68816 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 68816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 68816 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 68816 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 68816 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 68816 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 68816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 68816 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 68816 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 68816 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 68816 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 68816 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 68816 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 68816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 68816 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 68816 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 68816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 68816 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 68816 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 68816 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 68816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 68816 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 68816 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 68816 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 68816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 68816 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 68816 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 68816 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 68816 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 68816 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 68816 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 68816 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 68816 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 68816 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 68816 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 68816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 68816 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 68816 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 68816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 68816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 68816 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 68816 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 68816 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 68816 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 68816 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 68816 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 68816 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 68816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 68816 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 68816 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 68816 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 68816 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 68816 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 68816 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 68816 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 68816 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 68816 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 68816 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 68816 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 68816 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 68816 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 68816 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1649977179
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1649977179
transform -1 0 68816 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1649977179
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1649977179
transform -1 0 68816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1649977179
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1649977179
transform -1 0 68816 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1649977179
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1649977179
transform -1 0 68816 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1649977179
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1649977179
transform -1 0 68816 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1649977179
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1649977179
transform -1 0 68816 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1649977179
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1649977179
transform -1 0 68816 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1649977179
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1649977179
transform -1 0 68816 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1649977179
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1649977179
transform -1 0 68816 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1649977179
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1649977179
transform -1 0 68816 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1649977179
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1649977179
transform -1 0 68816 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1649977179
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1649977179
transform -1 0 68816 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1649977179
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1649977179
transform -1 0 68816 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1649977179
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1649977179
transform -1 0 68816 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1649977179
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1649977179
transform -1 0 68816 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1649977179
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1649977179
transform -1 0 68816 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1649977179
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1649977179
transform -1 0 68816 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1649977179
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1649977179
transform -1 0 68816 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1649977179
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1649977179
transform -1 0 68816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 60352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 62928 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 65504 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 68080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 62928 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 68080 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 60352 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 65504 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 62928 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 68080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 60352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 65504 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 62928 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 68080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 60352 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 65504 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 62928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 68080 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 60352 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 65504 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 62928 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 68080 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 60352 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 65504 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 62928 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 68080 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 60352 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 65504 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 62928 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 68080 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 60352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 65504 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 62928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 68080 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 60352 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 65504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 62928 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 68080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 60352 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 65504 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 62928 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 68080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 60352 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 65504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 62928 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 68080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 60352 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 65504 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 62928 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 68080 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 60352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 65504 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 62928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 68080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 60352 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 65504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 62928 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 68080 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 60352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 65504 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 62928 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 68080 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 60352 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 65504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 62928 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 68080 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 60352 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 65504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 62928 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 68080 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 60352 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 65504 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 62928 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 68080 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 60352 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 65504 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 62928 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 68080 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 60352 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 65504 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 62928 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 68080 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 60352 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 65504 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1649977179
transform 1 0 62928 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1649977179
transform 1 0 68080 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1649977179
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1649977179
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1649977179
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1649977179
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1649977179
transform 1 0 60352 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1649977179
transform 1 0 65504 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1649977179
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1649977179
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1649977179
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1649977179
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1649977179
transform 1 0 62928 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1649977179
transform 1 0 68080 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1649977179
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1649977179
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1649977179
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1649977179
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1649977179
transform 1 0 60352 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1649977179
transform 1 0 65504 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1649977179
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1649977179
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1649977179
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1649977179
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1649977179
transform 1 0 62928 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1649977179
transform 1 0 68080 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1649977179
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1649977179
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1649977179
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1649977179
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1649977179
transform 1 0 60352 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1649977179
transform 1 0 65504 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1649977179
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1649977179
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1649977179
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1649977179
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1649977179
transform 1 0 62928 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1649977179
transform 1 0 68080 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1649977179
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1649977179
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1649977179
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1649977179
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1649977179
transform 1 0 60352 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1649977179
transform 1 0 65504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1649977179
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1649977179
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1649977179
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1649977179
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1649977179
transform 1 0 62928 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1649977179
transform 1 0 68080 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1649977179
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1649977179
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1649977179
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1649977179
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1649977179
transform 1 0 60352 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1649977179
transform 1 0 65504 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1649977179
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1649977179
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1649977179
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1649977179
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1649977179
transform 1 0 62928 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1649977179
transform 1 0 68080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1649977179
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1649977179
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1649977179
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1649977179
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1649977179
transform 1 0 60352 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1649977179
transform 1 0 65504 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1649977179
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1649977179
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1649977179
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1649977179
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1649977179
transform 1 0 62928 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1649977179
transform 1 0 68080 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1649977179
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1649977179
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1649977179
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1649977179
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1649977179
transform 1 0 60352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1649977179
transform 1 0 65504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1649977179
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1649977179
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1649977179
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1649977179
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1649977179
transform 1 0 62928 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1649977179
transform 1 0 68080 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1649977179
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1649977179
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1649977179
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1649977179
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1649977179
transform 1 0 60352 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1649977179
transform 1 0 65504 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1649977179
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1649977179
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1649977179
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1649977179
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1649977179
transform 1 0 62928 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1649977179
transform 1 0 68080 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1649977179
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1649977179
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1649977179
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1649977179
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1649977179
transform 1 0 60352 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1649977179
transform 1 0 65504 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1649977179
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1649977179
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1649977179
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1649977179
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1649977179
transform 1 0 62928 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1649977179
transform 1 0 68080 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1649977179
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1649977179
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1649977179
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1649977179
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1649977179
transform 1 0 60352 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1649977179
transform 1 0 65504 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1649977179
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1649977179
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1649977179
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1649977179
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1649977179
transform 1 0 62928 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1649977179
transform 1 0 68080 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1649977179
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1649977179
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1649977179
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1649977179
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1649977179
transform 1 0 60352 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1649977179
transform 1 0 65504 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1649977179
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1649977179
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1649977179
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1649977179
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1649977179
transform 1 0 62928 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1649977179
transform 1 0 68080 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1649977179
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1649977179
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1649977179
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1649977179
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1649977179
transform 1 0 60352 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1649977179
transform 1 0 65504 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1649977179
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1649977179
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1649977179
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1649977179
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1649977179
transform 1 0 62928 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1649977179
transform 1 0 68080 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1649977179
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1649977179
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1649977179
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1649977179
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1649977179
transform 1 0 60352 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1649977179
transform 1 0 65504 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1649977179
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1649977179
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1649977179
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1649977179
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1649977179
transform 1 0 62928 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1649977179
transform 1 0 68080 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1649977179
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1649977179
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1649977179
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1649977179
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1649977179
transform 1 0 60352 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1649977179
transform 1 0 65504 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1649977179
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1649977179
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1649977179
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1649977179
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1649977179
transform 1 0 62928 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1649977179
transform 1 0 68080 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1649977179
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1649977179
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1649977179
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1649977179
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1649977179
transform 1 0 60352 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1649977179
transform 1 0 65504 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1649977179
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1649977179
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1649977179
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1649977179
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1649977179
transform 1 0 62928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1649977179
transform 1 0 68080 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1649977179
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1649977179
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1649977179
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1649977179
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1649977179
transform 1 0 60352 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1649977179
transform 1 0 65504 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1649977179
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1649977179
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1649977179
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1649977179
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1649977179
transform 1 0 62928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1649977179
transform 1 0 68080 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1649977179
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1649977179
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1649977179
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1649977179
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1649977179
transform 1 0 60352 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1649977179
transform 1 0 65504 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1649977179
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1649977179
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1649977179
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1649977179
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1649977179
transform 1 0 62928 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1649977179
transform 1 0 68080 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1649977179
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1649977179
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1649977179
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1649977179
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1649977179
transform 1 0 60352 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1649977179
transform 1 0 65504 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1649977179
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1649977179
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1649977179
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1649977179
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1649977179
transform 1 0 62928 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1649977179
transform 1 0 68080 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1649977179
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1649977179
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1649977179
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1649977179
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1649977179
transform 1 0 60352 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1649977179
transform 1 0 65504 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1649977179
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1649977179
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1649977179
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1649977179
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1649977179
transform 1 0 62928 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1649977179
transform 1 0 68080 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1649977179
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1649977179
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1649977179
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1649977179
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1649977179
transform 1 0 60352 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1649977179
transform 1 0 65504 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1649977179
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1649977179
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1649977179
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1649977179
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1649977179
transform 1 0 62928 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1649977179
transform 1 0 68080 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1649977179
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1649977179
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1649977179
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1649977179
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1649977179
transform 1 0 60352 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1649977179
transform 1 0 65504 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1649977179
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1649977179
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1649977179
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1649977179
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1649977179
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1649977179
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1649977179
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1649977179
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1649977179
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1649977179
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1649977179
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1649977179
transform 1 0 62928 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1649977179
transform 1 0 68080 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1649977179
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1649977179
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1649977179
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1649977179
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1649977179
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1649977179
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1649977179
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1649977179
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1649977179
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1649977179
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1649977179
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1649977179
transform 1 0 60352 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1649977179
transform 1 0 65504 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1649977179
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1649977179
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1649977179
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1649977179
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1649977179
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1649977179
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1649977179
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1649977179
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1649977179
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1649977179
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1649977179
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1649977179
transform 1 0 62928 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1649977179
transform 1 0 68080 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1649977179
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1649977179
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1649977179
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1649977179
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1649977179
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1649977179
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1649977179
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1649977179
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1649977179
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1649977179
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1649977179
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1649977179
transform 1 0 60352 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1649977179
transform 1 0 65504 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1348
timestamp 1649977179
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1349
timestamp 1649977179
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1350
timestamp 1649977179
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1351
timestamp 1649977179
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1352
timestamp 1649977179
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1353
timestamp 1649977179
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1354
timestamp 1649977179
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1355
timestamp 1649977179
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1356
timestamp 1649977179
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1357
timestamp 1649977179
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1358
timestamp 1649977179
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1359
timestamp 1649977179
transform 1 0 62928 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1360
timestamp 1649977179
transform 1 0 68080 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1361
timestamp 1649977179
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1362
timestamp 1649977179
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1363
timestamp 1649977179
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1364
timestamp 1649977179
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1365
timestamp 1649977179
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1366
timestamp 1649977179
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1367
timestamp 1649977179
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1368
timestamp 1649977179
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1369
timestamp 1649977179
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1370
timestamp 1649977179
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1371
timestamp 1649977179
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1372
timestamp 1649977179
transform 1 0 60352 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1373
timestamp 1649977179
transform 1 0 65504 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1374
timestamp 1649977179
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1375
timestamp 1649977179
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1376
timestamp 1649977179
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1377
timestamp 1649977179
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1378
timestamp 1649977179
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1379
timestamp 1649977179
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1380
timestamp 1649977179
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1381
timestamp 1649977179
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1382
timestamp 1649977179
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1383
timestamp 1649977179
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1384
timestamp 1649977179
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1385
timestamp 1649977179
transform 1 0 62928 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1386
timestamp 1649977179
transform 1 0 68080 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1387
timestamp 1649977179
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1388
timestamp 1649977179
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1389
timestamp 1649977179
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1390
timestamp 1649977179
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1391
timestamp 1649977179
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1392
timestamp 1649977179
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1393
timestamp 1649977179
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1394
timestamp 1649977179
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1395
timestamp 1649977179
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1396
timestamp 1649977179
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1397
timestamp 1649977179
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1398
timestamp 1649977179
transform 1 0 60352 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1399
timestamp 1649977179
transform 1 0 65504 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1400
timestamp 1649977179
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1401
timestamp 1649977179
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1402
timestamp 1649977179
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1403
timestamp 1649977179
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1404
timestamp 1649977179
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1405
timestamp 1649977179
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1406
timestamp 1649977179
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1407
timestamp 1649977179
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1408
timestamp 1649977179
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1409
timestamp 1649977179
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1410
timestamp 1649977179
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1411
timestamp 1649977179
transform 1 0 62928 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1412
timestamp 1649977179
transform 1 0 68080 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1413
timestamp 1649977179
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1414
timestamp 1649977179
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1415
timestamp 1649977179
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1416
timestamp 1649977179
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1417
timestamp 1649977179
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1418
timestamp 1649977179
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1419
timestamp 1649977179
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1420
timestamp 1649977179
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1421
timestamp 1649977179
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1422
timestamp 1649977179
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1423
timestamp 1649977179
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1424
timestamp 1649977179
transform 1 0 60352 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1425
timestamp 1649977179
transform 1 0 65504 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1426
timestamp 1649977179
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1427
timestamp 1649977179
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1428
timestamp 1649977179
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1429
timestamp 1649977179
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1430
timestamp 1649977179
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1431
timestamp 1649977179
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1432
timestamp 1649977179
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1433
timestamp 1649977179
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1434
timestamp 1649977179
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1435
timestamp 1649977179
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1436
timestamp 1649977179
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1437
timestamp 1649977179
transform 1 0 62928 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1438
timestamp 1649977179
transform 1 0 68080 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1439
timestamp 1649977179
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1440
timestamp 1649977179
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1441
timestamp 1649977179
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1442
timestamp 1649977179
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1443
timestamp 1649977179
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1444
timestamp 1649977179
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1445
timestamp 1649977179
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1446
timestamp 1649977179
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1447
timestamp 1649977179
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1448
timestamp 1649977179
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1449
timestamp 1649977179
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1450
timestamp 1649977179
transform 1 0 60352 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1451
timestamp 1649977179
transform 1 0 65504 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1452
timestamp 1649977179
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1453
timestamp 1649977179
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1454
timestamp 1649977179
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1455
timestamp 1649977179
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1456
timestamp 1649977179
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1457
timestamp 1649977179
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1458
timestamp 1649977179
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1459
timestamp 1649977179
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1460
timestamp 1649977179
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1461
timestamp 1649977179
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1462
timestamp 1649977179
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1463
timestamp 1649977179
transform 1 0 62928 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1464
timestamp 1649977179
transform 1 0 68080 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1465
timestamp 1649977179
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1466
timestamp 1649977179
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1467
timestamp 1649977179
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1468
timestamp 1649977179
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1469
timestamp 1649977179
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1470
timestamp 1649977179
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1471
timestamp 1649977179
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1472
timestamp 1649977179
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1473
timestamp 1649977179
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1474
timestamp 1649977179
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1475
timestamp 1649977179
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1476
timestamp 1649977179
transform 1 0 60352 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1477
timestamp 1649977179
transform 1 0 65504 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1478
timestamp 1649977179
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1479
timestamp 1649977179
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1480
timestamp 1649977179
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1481
timestamp 1649977179
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1482
timestamp 1649977179
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1483
timestamp 1649977179
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1484
timestamp 1649977179
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1485
timestamp 1649977179
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1486
timestamp 1649977179
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1487
timestamp 1649977179
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1488
timestamp 1649977179
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1489
timestamp 1649977179
transform 1 0 62928 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1490
timestamp 1649977179
transform 1 0 68080 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1491
timestamp 1649977179
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1492
timestamp 1649977179
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1493
timestamp 1649977179
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1494
timestamp 1649977179
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1495
timestamp 1649977179
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1496
timestamp 1649977179
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1497
timestamp 1649977179
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1498
timestamp 1649977179
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1499
timestamp 1649977179
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1500
timestamp 1649977179
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1501
timestamp 1649977179
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1502
timestamp 1649977179
transform 1 0 60352 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1503
timestamp 1649977179
transform 1 0 65504 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1504
timestamp 1649977179
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1505
timestamp 1649977179
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1506
timestamp 1649977179
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1507
timestamp 1649977179
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1508
timestamp 1649977179
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1509
timestamp 1649977179
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1510
timestamp 1649977179
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1511
timestamp 1649977179
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1512
timestamp 1649977179
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1513
timestamp 1649977179
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1514
timestamp 1649977179
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1515
timestamp 1649977179
transform 1 0 62928 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1516
timestamp 1649977179
transform 1 0 68080 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1517
timestamp 1649977179
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1518
timestamp 1649977179
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1519
timestamp 1649977179
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1520
timestamp 1649977179
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1521
timestamp 1649977179
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1522
timestamp 1649977179
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1523
timestamp 1649977179
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1524
timestamp 1649977179
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1525
timestamp 1649977179
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1526
timestamp 1649977179
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1527
timestamp 1649977179
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1528
timestamp 1649977179
transform 1 0 60352 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1529
timestamp 1649977179
transform 1 0 65504 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1530
timestamp 1649977179
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1531
timestamp 1649977179
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1532
timestamp 1649977179
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1533
timestamp 1649977179
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1534
timestamp 1649977179
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1535
timestamp 1649977179
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1536
timestamp 1649977179
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1537
timestamp 1649977179
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1538
timestamp 1649977179
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1539
timestamp 1649977179
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1540
timestamp 1649977179
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1541
timestamp 1649977179
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1542
timestamp 1649977179
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1543
timestamp 1649977179
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1544
timestamp 1649977179
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1545
timestamp 1649977179
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1546
timestamp 1649977179
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1547
timestamp 1649977179
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1548
timestamp 1649977179
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1549
timestamp 1649977179
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1550
timestamp 1649977179
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1551
timestamp 1649977179
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1552
timestamp 1649977179
transform 1 0 60352 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1553
timestamp 1649977179
transform 1 0 62928 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1554
timestamp 1649977179
transform 1 0 65504 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1555
timestamp 1649977179
transform 1 0 68080 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__or3b_2  _1022_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 46644 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1023_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 42872 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1024_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 42780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1025_
timestamp 1649977179
transform 1 0 44988 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1026_
timestamp 1649977179
transform 1 0 44988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1027_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 42964 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1029_
timestamp 1649977179
transform 1 0 35972 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1030_
timestamp 1649977179
transform 1 0 37720 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1031_
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1032_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 49128 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1033_
timestamp 1649977179
transform -1 0 51704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1034_
timestamp 1649977179
transform 1 0 41124 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1035_
timestamp 1649977179
transform 1 0 40204 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1036_
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1037_
timestamp 1649977179
transform 1 0 30084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1038_
timestamp 1649977179
transform 1 0 32660 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1039_
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1040_
timestamp 1649977179
transform 1 0 49128 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1041_
timestamp 1649977179
transform 1 0 51704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1042_
timestamp 1649977179
transform 1 0 48576 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1043_
timestamp 1649977179
transform 1 0 48208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1044_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20792 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1045_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20148 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1046_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23092 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1047_
timestamp 1649977179
transform 1 0 18400 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1048_
timestamp 1649977179
transform 1 0 22080 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1049_
timestamp 1649977179
transform 1 0 27324 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1050_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18032 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1051_
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1052_
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1053_
timestamp 1649977179
transform -1 0 23736 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1054_
timestamp 1649977179
transform 1 0 20516 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1055_
timestamp 1649977179
transform -1 0 17848 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1056_
timestamp 1649977179
transform 1 0 23092 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1057_
timestamp 1649977179
transform 1 0 20424 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1058_
timestamp 1649977179
transform 1 0 27048 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1059_
timestamp 1649977179
transform -1 0 22264 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1060_
timestamp 1649977179
transform 1 0 36432 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1061_
timestamp 1649977179
transform 1 0 26128 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1062_
timestamp 1649977179
transform 1 0 22080 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1063_
timestamp 1649977179
transform 1 0 27692 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _1064_
timestamp 1649977179
transform -1 0 27876 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1065_
timestamp 1649977179
transform 1 0 18124 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1066_
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1067_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 24840 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1068_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23644 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1069_
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1070_
timestamp 1649977179
transform -1 0 21252 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1071_
timestamp 1649977179
transform 1 0 20240 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1072_
timestamp 1649977179
transform -1 0 19688 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1073_
timestamp 1649977179
transform 1 0 17756 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1074_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18124 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1075_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18032 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1076_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17848 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1077_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17664 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1078_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17480 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1079_
timestamp 1649977179
transform -1 0 17020 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1080_
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1081_
timestamp 1649977179
transform -1 0 18768 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1082_
timestamp 1649977179
transform 1 0 18492 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1083_
timestamp 1649977179
transform -1 0 20884 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1084_
timestamp 1649977179
transform -1 0 20976 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1085_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19320 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1086_
timestamp 1649977179
transform 1 0 17112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1087_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20332 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1088_
timestamp 1649977179
transform -1 0 22080 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1089_
timestamp 1649977179
transform -1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1090_
timestamp 1649977179
transform -1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1091_
timestamp 1649977179
transform -1 0 22540 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1093_
timestamp 1649977179
transform -1 0 23644 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1094_
timestamp 1649977179
transform 1 0 23276 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1095_
timestamp 1649977179
transform -1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1096_
timestamp 1649977179
transform 1 0 40940 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1097_
timestamp 1649977179
transform 1 0 23552 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1098_
timestamp 1649977179
transform -1 0 23184 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1099_
timestamp 1649977179
transform 1 0 29716 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1649977179
transform -1 0 45264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1101_
timestamp 1649977179
transform 1 0 40848 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or4b_1  _1102_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 42136 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1103_
timestamp 1649977179
transform -1 0 41216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1104_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43700 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1105_
timestamp 1649977179
transform -1 0 43332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1106_
timestamp 1649977179
transform 1 0 40388 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1107_
timestamp 1649977179
transform 1 0 40756 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1108_
timestamp 1649977179
transform -1 0 40388 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1109_
timestamp 1649977179
transform 1 0 41584 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1110_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 40020 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1111_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43792 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1112_
timestamp 1649977179
transform 1 0 41124 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1113_
timestamp 1649977179
transform 1 0 38180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1114_
timestamp 1649977179
transform 1 0 40296 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1115_
timestamp 1649977179
transform 1 0 41584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1116_
timestamp 1649977179
transform 1 0 42504 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1117_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 40848 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1118_
timestamp 1649977179
transform -1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1119_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 40112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1120_
timestamp 1649977179
transform 1 0 39836 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1121_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 50140 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1122_
timestamp 1649977179
transform -1 0 51428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1123_
timestamp 1649977179
transform -1 0 49220 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _1124_
timestamp 1649977179
transform -1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1125_
timestamp 1649977179
transform 1 0 48576 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1126_
timestamp 1649977179
transform -1 0 49496 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1127_
timestamp 1649977179
transform 1 0 46828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1128_
timestamp 1649977179
transform 1 0 48024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1129_
timestamp 1649977179
transform -1 0 49128 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1130_
timestamp 1649977179
transform 1 0 47748 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1131_
timestamp 1649977179
transform 1 0 48300 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1132_
timestamp 1649977179
transform 1 0 46092 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1133_
timestamp 1649977179
transform -1 0 47656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1134_
timestamp 1649977179
transform 1 0 49312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1135_
timestamp 1649977179
transform 1 0 50140 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1136_
timestamp 1649977179
transform -1 0 50876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1137_
timestamp 1649977179
transform 1 0 48024 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1138_
timestamp 1649977179
transform 1 0 51704 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1139_
timestamp 1649977179
transform -1 0 50876 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1140_
timestamp 1649977179
transform -1 0 50600 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1141_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 48944 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1142_
timestamp 1649977179
transform 1 0 50692 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1143_
timestamp 1649977179
transform -1 0 51520 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1144_
timestamp 1649977179
transform 1 0 50140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1649977179
transform 1 0 51152 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a2111oi_1  _1146_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 49588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1649977179
transform -1 0 34960 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1148_
timestamp 1649977179
transform 1 0 34868 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1149_
timestamp 1649977179
transform 1 0 35052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1150_
timestamp 1649977179
transform 1 0 44988 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1151_
timestamp 1649977179
transform -1 0 45908 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1152_
timestamp 1649977179
transform -1 0 37904 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1153_
timestamp 1649977179
transform -1 0 37536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1154_
timestamp 1649977179
transform -1 0 45540 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1155_
timestamp 1649977179
transform -1 0 45172 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1156_
timestamp 1649977179
transform 1 0 40756 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1157_
timestamp 1649977179
transform -1 0 41492 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1158_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 49220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1159_
timestamp 1649977179
transform 1 0 46828 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1160_
timestamp 1649977179
transform -1 0 50232 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _1161_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 47196 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1162_
timestamp 1649977179
transform -1 0 47932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1163_
timestamp 1649977179
transform 1 0 50140 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1164_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 49404 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1165_
timestamp 1649977179
transform -1 0 49680 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1166_
timestamp 1649977179
transform 1 0 48392 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1649977179
transform 1 0 48668 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1168_
timestamp 1649977179
transform -1 0 50232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1169_
timestamp 1649977179
transform 1 0 48116 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1170_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 50140 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1171_
timestamp 1649977179
transform -1 0 48024 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1172_
timestamp 1649977179
transform 1 0 47196 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1173_
timestamp 1649977179
transform -1 0 48208 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1174_
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1175_
timestamp 1649977179
transform -1 0 49496 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1176_
timestamp 1649977179
transform 1 0 51244 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1177_
timestamp 1649977179
transform -1 0 22080 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1178_
timestamp 1649977179
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1179_
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1180_
timestamp 1649977179
transform -1 0 20976 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1181_
timestamp 1649977179
transform -1 0 22356 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _1182_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20424 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1649977179
transform 1 0 17756 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1184_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19412 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1185_
timestamp 1649977179
transform 1 0 20516 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1186_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20148 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1187_
timestamp 1649977179
transform -1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1188_
timestamp 1649977179
transform 1 0 21988 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1189_
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1190_
timestamp 1649977179
transform 1 0 20240 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1191_
timestamp 1649977179
transform -1 0 22172 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1192_
timestamp 1649977179
transform 1 0 17940 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1193_
timestamp 1649977179
transform 1 0 19688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1194_
timestamp 1649977179
transform -1 0 15456 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1195_
timestamp 1649977179
transform -1 0 14996 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a2bb2o_1  _1196_
timestamp 1649977179
transform -1 0 19320 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1197_
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1198_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1199_
timestamp 1649977179
transform 1 0 17664 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1200_
timestamp 1649977179
transform 1 0 17664 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1649977179
transform 1 0 17480 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1202_
timestamp 1649977179
transform 1 0 19320 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1203_
timestamp 1649977179
transform -1 0 22356 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1204_
timestamp 1649977179
transform 1 0 21160 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1205_
timestamp 1649977179
transform 1 0 20976 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1206_
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1207_
timestamp 1649977179
transform -1 0 21068 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1208_
timestamp 1649977179
transform -1 0 20516 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1209_
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1210_
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1211_
timestamp 1649977179
transform -1 0 34684 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1212_
timestamp 1649977179
transform 1 0 18768 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1213_
timestamp 1649977179
transform -1 0 20792 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1214_
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1215_
timestamp 1649977179
transform -1 0 21344 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1216_
timestamp 1649977179
transform 1 0 20332 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1217_
timestamp 1649977179
transform -1 0 20148 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1218_
timestamp 1649977179
transform 1 0 19872 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1219_
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1220_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19504 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1221_
timestamp 1649977179
transform 1 0 27232 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _1222_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 34132 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1223_
timestamp 1649977179
transform -1 0 19504 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1224_
timestamp 1649977179
transform 1 0 35052 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1225_
timestamp 1649977179
transform 1 0 18032 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1226_
timestamp 1649977179
transform -1 0 35420 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1227_
timestamp 1649977179
transform -1 0 37260 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1228_
timestamp 1649977179
transform 1 0 35972 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1229_
timestamp 1649977179
transform -1 0 38548 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1230_
timestamp 1649977179
transform 1 0 35236 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1231_
timestamp 1649977179
transform 1 0 22356 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1232_
timestamp 1649977179
transform 1 0 35880 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1233_
timestamp 1649977179
transform -1 0 36800 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1234_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 41952 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_2  _1235_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30452 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _1236_
timestamp 1649977179
transform 1 0 23184 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1237_
timestamp 1649977179
transform 1 0 35696 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1238_
timestamp 1649977179
transform 1 0 38732 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1239_
timestamp 1649977179
transform 1 0 38548 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1240_
timestamp 1649977179
transform 1 0 37904 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1241_
timestamp 1649977179
transform -1 0 41216 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1242_
timestamp 1649977179
transform 1 0 40204 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1243_
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1244_
timestamp 1649977179
transform 1 0 39836 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1245_
timestamp 1649977179
transform 1 0 39836 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1246_
timestamp 1649977179
transform 1 0 42044 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1247_
timestamp 1649977179
transform -1 0 46184 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_1  _1248_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 41860 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1249_
timestamp 1649977179
transform 1 0 41216 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1250_
timestamp 1649977179
transform 1 0 42504 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1251_
timestamp 1649977179
transform 1 0 39100 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1252_
timestamp 1649977179
transform 1 0 43056 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1253_
timestamp 1649977179
transform -1 0 44804 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1254_
timestamp 1649977179
transform 1 0 42872 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1255_
timestamp 1649977179
transform 1 0 18768 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1256_
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1257_
timestamp 1649977179
transform -1 0 41400 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _1258_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 40480 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1259_
timestamp 1649977179
transform -1 0 29440 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1260_
timestamp 1649977179
transform 1 0 31648 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1261_
timestamp 1649977179
transform 1 0 23092 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1262_
timestamp 1649977179
transform 1 0 37444 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1263_
timestamp 1649977179
transform 1 0 37444 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1264_
timestamp 1649977179
transform -1 0 38272 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1265_
timestamp 1649977179
transform -1 0 40388 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 1649977179
transform -1 0 36892 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1267_
timestamp 1649977179
transform 1 0 39836 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1268_
timestamp 1649977179
transform -1 0 40848 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1269_
timestamp 1649977179
transform 1 0 43884 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1270_
timestamp 1649977179
transform 1 0 45448 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1271_
timestamp 1649977179
transform 1 0 46000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1272_
timestamp 1649977179
transform 1 0 41216 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1273_
timestamp 1649977179
transform 1 0 42412 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1274_
timestamp 1649977179
transform 1 0 42964 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _1275_
timestamp 1649977179
transform 1 0 40848 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1276_
timestamp 1649977179
transform 1 0 39836 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1277_
timestamp 1649977179
transform 1 0 40848 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _1278_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 44988 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1279_
timestamp 1649977179
transform 1 0 39468 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1280_
timestamp 1649977179
transform 1 0 40480 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1281_
timestamp 1649977179
transform 1 0 40112 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1282_
timestamp 1649977179
transform 1 0 40020 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1283_
timestamp 1649977179
transform -1 0 40664 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1284_
timestamp 1649977179
transform -1 0 22264 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1285_
timestamp 1649977179
transform 1 0 23276 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1286_
timestamp 1649977179
transform 1 0 39284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1287_
timestamp 1649977179
transform -1 0 39376 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1288_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 39560 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1289_
timestamp 1649977179
transform 1 0 40664 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1290_
timestamp 1649977179
transform -1 0 39100 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1291_
timestamp 1649977179
transform 1 0 38364 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1292_
timestamp 1649977179
transform 1 0 39836 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1293_
timestamp 1649977179
transform 1 0 39652 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1294_
timestamp 1649977179
transform -1 0 41492 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1295_
timestamp 1649977179
transform 1 0 40480 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1296_
timestamp 1649977179
transform -1 0 41860 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1297_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 38640 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1298_
timestamp 1649977179
transform 1 0 38456 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1299_
timestamp 1649977179
transform 1 0 39468 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1300_
timestamp 1649977179
transform -1 0 40756 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1301_
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1302_
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1303_
timestamp 1649977179
transform 1 0 37260 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1304_
timestamp 1649977179
transform -1 0 38640 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1305_
timestamp 1649977179
transform 1 0 37260 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1306_
timestamp 1649977179
transform -1 0 19780 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1307_
timestamp 1649977179
transform 1 0 37352 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1308_
timestamp 1649977179
transform 1 0 37812 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1309_
timestamp 1649977179
transform 1 0 39836 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1310_
timestamp 1649977179
transform -1 0 42964 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1311_
timestamp 1649977179
transform -1 0 9384 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1312_
timestamp 1649977179
transform 1 0 8004 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1313_
timestamp 1649977179
transform 1 0 8648 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1314_
timestamp 1649977179
transform -1 0 12696 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1315_
timestamp 1649977179
transform 1 0 9752 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1316_
timestamp 1649977179
transform -1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _1317_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10948 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1318_
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1319_
timestamp 1649977179
transform -1 0 13892 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1320_
timestamp 1649977179
transform 1 0 12512 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1321_
timestamp 1649977179
transform -1 0 10856 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1322_
timestamp 1649977179
transform 1 0 7084 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1323_
timestamp 1649977179
transform 1 0 4784 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1324_
timestamp 1649977179
transform 1 0 8096 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1325_
timestamp 1649977179
transform -1 0 11040 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1326_
timestamp 1649977179
transform -1 0 14536 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1327_
timestamp 1649977179
transform 1 0 8924 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1328_
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1329_
timestamp 1649977179
transform 1 0 7912 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1330_
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1331_
timestamp 1649977179
transform -1 0 9016 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1332_
timestamp 1649977179
transform 1 0 25392 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1333_
timestamp 1649977179
transform 1 0 6440 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1334_
timestamp 1649977179
transform 1 0 6716 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1335_
timestamp 1649977179
transform -1 0 8648 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1336_
timestamp 1649977179
transform -1 0 12052 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1337_
timestamp 1649977179
transform 1 0 12788 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1338_
timestamp 1649977179
transform -1 0 11408 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_1  _1339_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10396 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_1  _1340_
timestamp 1649977179
transform -1 0 9752 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1341_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10764 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1342_
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1343_
timestamp 1649977179
transform 1 0 9384 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1344_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1345_
timestamp 1649977179
transform 1 0 6532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1346_
timestamp 1649977179
transform -1 0 8004 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1347_
timestamp 1649977179
transform -1 0 8372 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1348_
timestamp 1649977179
transform 1 0 22632 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1349_
timestamp 1649977179
transform 1 0 10028 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1350_
timestamp 1649977179
transform 1 0 12512 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1351_
timestamp 1649977179
transform -1 0 7728 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1352_
timestamp 1649977179
transform 1 0 6072 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1353_
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1354_
timestamp 1649977179
transform -1 0 7636 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1355_
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1356_
timestamp 1649977179
transform -1 0 9844 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1357_
timestamp 1649977179
transform -1 0 9476 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1358_
timestamp 1649977179
transform 1 0 13064 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1359_
timestamp 1649977179
transform 1 0 12420 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1360_
timestamp 1649977179
transform 1 0 10396 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1361_
timestamp 1649977179
transform -1 0 11592 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1362_
timestamp 1649977179
transform -1 0 12144 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1363_
timestamp 1649977179
transform -1 0 11040 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1364_
timestamp 1649977179
transform 1 0 10396 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1365_
timestamp 1649977179
transform 1 0 7636 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1366_
timestamp 1649977179
transform -1 0 8464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1367_
timestamp 1649977179
transform 1 0 6900 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1368_
timestamp 1649977179
transform 1 0 7268 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1369_
timestamp 1649977179
transform 1 0 7268 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1370_
timestamp 1649977179
transform 1 0 5152 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1371_
timestamp 1649977179
transform 1 0 6808 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1372_
timestamp 1649977179
transform -1 0 8464 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1373_
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1374_
timestamp 1649977179
transform -1 0 9384 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1375_
timestamp 1649977179
transform -1 0 9568 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1376_
timestamp 1649977179
transform -1 0 8556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1377_
timestamp 1649977179
transform -1 0 8464 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1378_
timestamp 1649977179
transform 1 0 7360 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1379_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1380_
timestamp 1649977179
transform -1 0 7176 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1381_
timestamp 1649977179
transform 1 0 6440 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_1  _1382_
timestamp 1649977179
transform -1 0 9568 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1383_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1384_
timestamp 1649977179
transform -1 0 6992 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1385_
timestamp 1649977179
transform 1 0 4784 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1386_
timestamp 1649977179
transform 1 0 5428 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1387_
timestamp 1649977179
transform 1 0 4140 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1388_
timestamp 1649977179
transform -1 0 6624 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1389_
timestamp 1649977179
transform 1 0 5152 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1390_
timestamp 1649977179
transform 1 0 6072 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1391_
timestamp 1649977179
transform -1 0 5152 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1392_
timestamp 1649977179
transform 1 0 4416 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1393_
timestamp 1649977179
transform 1 0 5336 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1394_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1395_
timestamp 1649977179
transform -1 0 36616 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1396_
timestamp 1649977179
transform 1 0 25116 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1397_
timestamp 1649977179
transform 1 0 25300 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1398_
timestamp 1649977179
transform -1 0 26864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1399_
timestamp 1649977179
transform 1 0 24472 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1400_
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1401_
timestamp 1649977179
transform 1 0 32384 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1402_
timestamp 1649977179
transform 1 0 32476 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1403_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 32568 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1404_
timestamp 1649977179
transform 1 0 33304 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1405_
timestamp 1649977179
transform -1 0 47012 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1406_
timestamp 1649977179
transform -1 0 35328 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1407_
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1408_
timestamp 1649977179
transform -1 0 32660 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1409_
timestamp 1649977179
transform 1 0 31096 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1410_
timestamp 1649977179
transform -1 0 32476 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1411_
timestamp 1649977179
transform 1 0 32844 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1412_
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1413_
timestamp 1649977179
transform 1 0 24656 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1414_
timestamp 1649977179
transform -1 0 26128 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1415_
timestamp 1649977179
transform 1 0 22632 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1416_
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1417_
timestamp 1649977179
transform 1 0 23460 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1418_
timestamp 1649977179
transform 1 0 25760 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1419_
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1420_
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1421_
timestamp 1649977179
transform -1 0 29072 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1422_
timestamp 1649977179
transform -1 0 27968 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1423_
timestamp 1649977179
transform 1 0 33120 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1424_
timestamp 1649977179
transform -1 0 44436 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1425_
timestamp 1649977179
transform -1 0 43516 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1426_
timestamp 1649977179
transform 1 0 46092 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1427_
timestamp 1649977179
transform 1 0 25944 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1428_
timestamp 1649977179
transform 1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1429_
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1430_
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1431_
timestamp 1649977179
transform 1 0 27968 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1432_
timestamp 1649977179
transform -1 0 28612 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _1433_
timestamp 1649977179
transform -1 0 28612 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1434_
timestamp 1649977179
transform 1 0 23276 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1435_
timestamp 1649977179
transform -1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1436_
timestamp 1649977179
transform 1 0 25484 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1437_
timestamp 1649977179
transform 1 0 24564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1438_
timestamp 1649977179
transform 1 0 24748 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1439_
timestamp 1649977179
transform 1 0 25668 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1440_
timestamp 1649977179
transform 1 0 23276 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1441_
timestamp 1649977179
transform 1 0 24196 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1442_
timestamp 1649977179
transform -1 0 27232 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1443_
timestamp 1649977179
transform 1 0 28888 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1444_
timestamp 1649977179
transform 1 0 27784 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1445_
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1446_
timestamp 1649977179
transform 1 0 31004 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1447_
timestamp 1649977179
transform 1 0 25760 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1448_
timestamp 1649977179
transform 1 0 25668 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1449_
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1450_
timestamp 1649977179
transform 1 0 26864 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1451_
timestamp 1649977179
transform 1 0 27692 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1452_
timestamp 1649977179
transform 1 0 31924 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1453_
timestamp 1649977179
transform -1 0 35052 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1454_
timestamp 1649977179
transform -1 0 34408 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1455_
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1456_
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1457_
timestamp 1649977179
transform -1 0 30176 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1458_
timestamp 1649977179
transform 1 0 29256 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1459_
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1460_
timestamp 1649977179
transform 1 0 31832 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_2  _1461_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32568 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _1462_
timestamp 1649977179
transform 1 0 25392 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1463_
timestamp 1649977179
transform 1 0 24472 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1464_
timestamp 1649977179
transform 1 0 24472 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1465_
timestamp 1649977179
transform 1 0 25300 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1466_
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1467_
timestamp 1649977179
transform 1 0 27600 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1468_
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1469_
timestamp 1649977179
transform -1 0 29072 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1470_
timestamp 1649977179
transform 1 0 24840 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1471_
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1472_
timestamp 1649977179
transform -1 0 27232 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1473_
timestamp 1649977179
transform 1 0 25760 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1474_
timestamp 1649977179
transform 1 0 27232 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1475_
timestamp 1649977179
transform -1 0 28888 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1476_
timestamp 1649977179
transform 1 0 31096 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1477_
timestamp 1649977179
transform 1 0 32108 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1478_
timestamp 1649977179
transform 1 0 32936 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1479_
timestamp 1649977179
transform -1 0 45724 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1480_
timestamp 1649977179
transform -1 0 16652 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1481_
timestamp 1649977179
transform -1 0 15272 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1482_
timestamp 1649977179
transform 1 0 14536 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1483_
timestamp 1649977179
transform -1 0 13156 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1484_
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1485_
timestamp 1649977179
transform -1 0 10856 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1486_
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1487_
timestamp 1649977179
transform 1 0 8924 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1488_
timestamp 1649977179
transform -1 0 11040 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1489_
timestamp 1649977179
transform -1 0 18308 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1490_
timestamp 1649977179
transform 1 0 10948 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1491_
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1492_
timestamp 1649977179
transform 1 0 14260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1493_
timestamp 1649977179
transform 1 0 14260 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1494_
timestamp 1649977179
transform 1 0 14628 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1495_
timestamp 1649977179
transform -1 0 38732 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _1496_
timestamp 1649977179
transform -1 0 17480 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1497_
timestamp 1649977179
transform -1 0 15456 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1498_
timestamp 1649977179
transform 1 0 15640 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1499_
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1500_
timestamp 1649977179
transform -1 0 17296 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1501_
timestamp 1649977179
transform 1 0 14720 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1502_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1503_
timestamp 1649977179
transform 1 0 16468 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1504_
timestamp 1649977179
transform 1 0 42780 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1505_
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1506_
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1507_
timestamp 1649977179
transform -1 0 16284 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1508_
timestamp 1649977179
transform -1 0 16192 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1509_
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1510_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_2  _1511_
timestamp 1649977179
transform -1 0 16836 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1512_
timestamp 1649977179
transform 1 0 12512 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1513_
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1514_
timestamp 1649977179
transform -1 0 10396 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1515_
timestamp 1649977179
transform 1 0 8280 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1516_
timestamp 1649977179
transform -1 0 9568 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1517_
timestamp 1649977179
transform -1 0 9292 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1518_
timestamp 1649977179
transform -1 0 11776 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1519_
timestamp 1649977179
transform 1 0 11592 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1520_
timestamp 1649977179
transform 1 0 12696 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1521_
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1522_
timestamp 1649977179
transform 1 0 13800 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1523_
timestamp 1649977179
transform 1 0 15180 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1524_
timestamp 1649977179
transform -1 0 14812 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1525_
timestamp 1649977179
transform -1 0 10856 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1526_
timestamp 1649977179
transform -1 0 12144 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1527_
timestamp 1649977179
transform 1 0 9660 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1528_
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1529_
timestamp 1649977179
transform 1 0 17112 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1530_
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1531_
timestamp 1649977179
transform -1 0 15088 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1532_
timestamp 1649977179
transform -1 0 15824 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1533_
timestamp 1649977179
transform -1 0 14352 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1534_
timestamp 1649977179
transform -1 0 15640 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1535_
timestamp 1649977179
transform 1 0 11776 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1536_
timestamp 1649977179
transform -1 0 14812 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1537_
timestamp 1649977179
transform 1 0 12144 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1538_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1539_
timestamp 1649977179
transform 1 0 9200 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1540_
timestamp 1649977179
transform -1 0 12972 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1541_
timestamp 1649977179
transform 1 0 11868 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _1542_
timestamp 1649977179
transform -1 0 12696 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1543_
timestamp 1649977179
transform -1 0 13708 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1544_
timestamp 1649977179
transform 1 0 12788 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1545_
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1546_
timestamp 1649977179
transform 1 0 9476 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1547_
timestamp 1649977179
transform -1 0 12972 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1548_
timestamp 1649977179
transform 1 0 8832 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1549_
timestamp 1649977179
transform -1 0 10948 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1550_
timestamp 1649977179
transform 1 0 8924 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1551_
timestamp 1649977179
transform -1 0 9660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1552_
timestamp 1649977179
transform 1 0 6716 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1553_
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1554_
timestamp 1649977179
transform 1 0 9936 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1555_
timestamp 1649977179
transform -1 0 14628 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1556_
timestamp 1649977179
transform 1 0 12328 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1557_
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1558_
timestamp 1649977179
transform -1 0 43792 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1559_
timestamp 1649977179
transform 1 0 20424 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1560_
timestamp 1649977179
transform 1 0 20516 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1561_
timestamp 1649977179
transform -1 0 22724 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1562_
timestamp 1649977179
transform 1 0 20700 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1563_
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1564_
timestamp 1649977179
transform 1 0 25116 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1565_
timestamp 1649977179
transform 1 0 24104 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1566_
timestamp 1649977179
transform -1 0 26680 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1567_
timestamp 1649977179
transform -1 0 36156 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1568_
timestamp 1649977179
transform 1 0 27508 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1569_
timestamp 1649977179
transform -1 0 28888 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1570_
timestamp 1649977179
transform 1 0 28336 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1571_
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1572_
timestamp 1649977179
transform 1 0 30452 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1573_
timestamp 1649977179
transform 1 0 28428 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1574_
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1575_
timestamp 1649977179
transform 1 0 29716 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1576_
timestamp 1649977179
transform 1 0 30544 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1577_
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1578_
timestamp 1649977179
transform 1 0 25300 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1579_
timestamp 1649977179
transform -1 0 27232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1580_
timestamp 1649977179
transform 1 0 25024 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1581_
timestamp 1649977179
transform -1 0 26864 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1582_
timestamp 1649977179
transform -1 0 26496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1583_
timestamp 1649977179
transform 1 0 27968 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1584_
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1585_
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1586_
timestamp 1649977179
transform -1 0 40388 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1587_
timestamp 1649977179
transform -1 0 40112 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1588_
timestamp 1649977179
transform -1 0 29072 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1589_
timestamp 1649977179
transform 1 0 25300 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1590_
timestamp 1649977179
transform 1 0 25944 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1591_
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1592_
timestamp 1649977179
transform -1 0 25392 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221ai_4  _1593_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 27140 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__nand2_1  _1594_
timestamp 1649977179
transform 1 0 28980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1595_
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1596_
timestamp 1649977179
transform 1 0 28520 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1597_
timestamp 1649977179
transform -1 0 27968 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1598_
timestamp 1649977179
transform 1 0 29072 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1599_
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1600_
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1601_
timestamp 1649977179
transform 1 0 19504 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1602_
timestamp 1649977179
transform -1 0 20056 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1603_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 30176 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1604_
timestamp 1649977179
transform -1 0 30912 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1605_
timestamp 1649977179
transform 1 0 32752 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1606_
timestamp 1649977179
transform -1 0 30176 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1607_
timestamp 1649977179
transform -1 0 30452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1608_
timestamp 1649977179
transform 1 0 31280 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1609_
timestamp 1649977179
transform 1 0 28520 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1610_
timestamp 1649977179
transform 1 0 29072 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1611_
timestamp 1649977179
transform 1 0 30360 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1612_
timestamp 1649977179
transform 1 0 25668 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1613_
timestamp 1649977179
transform -1 0 31188 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1614_
timestamp 1649977179
transform 1 0 25668 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1615_
timestamp 1649977179
transform 1 0 26036 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1616_
timestamp 1649977179
transform 1 0 28152 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1617_
timestamp 1649977179
transform 1 0 28704 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_2  _1618_
timestamp 1649977179
transform 1 0 30452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__xor2_1  _1619_
timestamp 1649977179
transform 1 0 29900 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1620_
timestamp 1649977179
transform 1 0 32476 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1621_
timestamp 1649977179
transform 1 0 32016 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1622_
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1623_
timestamp 1649977179
transform -1 0 32568 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1624_
timestamp 1649977179
transform 1 0 35972 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1625_
timestamp 1649977179
transform -1 0 37904 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1626_
timestamp 1649977179
transform 1 0 30176 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1627_
timestamp 1649977179
transform 1 0 32108 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1628_
timestamp 1649977179
transform 1 0 29348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1629_
timestamp 1649977179
transform 1 0 29808 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1630_
timestamp 1649977179
transform 1 0 31096 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1631_
timestamp 1649977179
transform 1 0 27876 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1632_
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1633_
timestamp 1649977179
transform 1 0 28152 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1634_
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1635_
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1636_
timestamp 1649977179
transform 1 0 33120 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1637_
timestamp 1649977179
transform 1 0 33672 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1638_
timestamp 1649977179
transform 1 0 38640 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1639_
timestamp 1649977179
transform 1 0 48484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1640_
timestamp 1649977179
transform -1 0 42136 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1641_
timestamp 1649977179
transform -1 0 39376 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1642_
timestamp 1649977179
transform -1 0 46368 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1643_
timestamp 1649977179
transform 1 0 44252 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1644_
timestamp 1649977179
transform 1 0 46092 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1645_
timestamp 1649977179
transform -1 0 47196 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1646_
timestamp 1649977179
transform 1 0 38456 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1647_
timestamp 1649977179
transform 1 0 40112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1648_
timestamp 1649977179
transform 1 0 44068 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1649_
timestamp 1649977179
transform -1 0 45264 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1650_
timestamp 1649977179
transform 1 0 35144 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1651_
timestamp 1649977179
transform 1 0 35696 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1652_
timestamp 1649977179
transform 1 0 50140 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1653_
timestamp 1649977179
transform 1 0 52072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1654_
timestamp 1649977179
transform -1 0 48576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1655_
timestamp 1649977179
transform 1 0 42044 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1656_
timestamp 1649977179
transform 1 0 42780 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1657_
timestamp 1649977179
transform 1 0 43516 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1658_
timestamp 1649977179
transform -1 0 39744 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1659_
timestamp 1649977179
transform -1 0 40112 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1660_
timestamp 1649977179
transform 1 0 40940 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1661_
timestamp 1649977179
transform 1 0 44160 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1662_
timestamp 1649977179
transform 1 0 15180 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1663_
timestamp 1649977179
transform 1 0 13984 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1664_
timestamp 1649977179
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1665_
timestamp 1649977179
transform 1 0 12696 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1666_
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1667_
timestamp 1649977179
transform -1 0 18216 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1668_
timestamp 1649977179
transform -1 0 15364 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1669_
timestamp 1649977179
transform 1 0 16468 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1670_
timestamp 1649977179
transform -1 0 16468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1671_
timestamp 1649977179
transform 1 0 18032 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1672_
timestamp 1649977179
transform 1 0 19320 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1673_
timestamp 1649977179
transform -1 0 18676 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1674_
timestamp 1649977179
transform 1 0 14720 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1675_
timestamp 1649977179
transform 1 0 19136 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1676_
timestamp 1649977179
transform -1 0 19320 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1677_
timestamp 1649977179
transform 1 0 16008 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1678_
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1679_
timestamp 1649977179
transform -1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1680_
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1681_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1682_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1683_
timestamp 1649977179
transform 1 0 15364 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1684_
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1685_
timestamp 1649977179
transform -1 0 17112 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1686_
timestamp 1649977179
transform 1 0 13156 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1687_
timestamp 1649977179
transform -1 0 17388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1688_
timestamp 1649977179
transform 1 0 15272 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1689_
timestamp 1649977179
transform -1 0 14352 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1690_
timestamp 1649977179
transform 1 0 15640 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1691_
timestamp 1649977179
transform -1 0 14904 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1692_
timestamp 1649977179
transform 1 0 14628 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1693_
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1694_
timestamp 1649977179
transform 1 0 15272 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1695_
timestamp 1649977179
transform 1 0 15180 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1696_
timestamp 1649977179
transform 1 0 17848 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1697_
timestamp 1649977179
transform 1 0 15272 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1698_
timestamp 1649977179
transform 1 0 14904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1699_
timestamp 1649977179
transform 1 0 16376 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1700_
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1701_
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1702_
timestamp 1649977179
transform 1 0 16928 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1703_
timestamp 1649977179
transform 1 0 16652 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1704_
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1705_
timestamp 1649977179
transform 1 0 31188 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1706_
timestamp 1649977179
transform 1 0 23460 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1707_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1708_
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1709_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1710_
timestamp 1649977179
transform 1 0 36616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1711_
timestamp 1649977179
transform 1 0 43240 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1649977179
transform -1 0 43332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1713_
timestamp 1649977179
transform 1 0 29532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1714_
timestamp 1649977179
transform 1 0 43700 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1715_
timestamp 1649977179
transform -1 0 43516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1716_
timestamp 1649977179
transform 1 0 28244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1717_
timestamp 1649977179
transform 1 0 37260 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1718_
timestamp 1649977179
transform -1 0 37536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1719_
timestamp 1649977179
transform 1 0 27416 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1720_
timestamp 1649977179
transform -1 0 39284 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1721_
timestamp 1649977179
transform 1 0 39836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1722_
timestamp 1649977179
transform 1 0 24840 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1723_
timestamp 1649977179
transform -1 0 38456 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1724_
timestamp 1649977179
transform 1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1725_
timestamp 1649977179
transform -1 0 25300 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1726_
timestamp 1649977179
transform 1 0 36524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1727_
timestamp 1649977179
transform -1 0 35696 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1728_
timestamp 1649977179
transform 1 0 35052 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1729_
timestamp 1649977179
transform 1 0 20148 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1730_
timestamp 1649977179
transform -1 0 41952 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1731_
timestamp 1649977179
transform -1 0 42688 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1732_
timestamp 1649977179
transform 1 0 20976 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1733_
timestamp 1649977179
transform -1 0 41860 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1734_
timestamp 1649977179
transform -1 0 42504 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1735_
timestamp 1649977179
transform 1 0 20056 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1736_
timestamp 1649977179
transform -1 0 41584 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1737_
timestamp 1649977179
transform -1 0 42136 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1738_
timestamp 1649977179
transform 1 0 19596 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1739_
timestamp 1649977179
transform 1 0 36984 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1740_
timestamp 1649977179
transform -1 0 36800 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1741_
timestamp 1649977179
transform 1 0 19596 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1742_
timestamp 1649977179
transform 1 0 34868 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1743_
timestamp 1649977179
transform -1 0 34040 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1744_
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1745_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _1746_
timestamp 1649977179
transform -1 0 24656 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1747_
timestamp 1649977179
transform 1 0 35328 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1748_
timestamp 1649977179
transform 1 0 42136 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1749_
timestamp 1649977179
transform -1 0 41952 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1750_
timestamp 1649977179
transform -1 0 44160 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1751_
timestamp 1649977179
transform 1 0 43976 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1752_
timestamp 1649977179
transform 1 0 37720 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1753_
timestamp 1649977179
transform 1 0 36156 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1754_
timestamp 1649977179
transform -1 0 39284 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1755_
timestamp 1649977179
transform 1 0 38916 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1756_
timestamp 1649977179
transform 1 0 31924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1757_
timestamp 1649977179
transform 1 0 30728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1758_
timestamp 1649977179
transform -1 0 35604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1759_
timestamp 1649977179
transform 1 0 34684 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1760_
timestamp 1649977179
transform -1 0 34776 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1761_
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1762_
timestamp 1649977179
transform 1 0 36248 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1763_
timestamp 1649977179
transform 1 0 35972 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1764_
timestamp 1649977179
transform -1 0 35604 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1765_
timestamp 1649977179
transform 1 0 34132 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1766_
timestamp 1649977179
transform -1 0 33764 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1767_
timestamp 1649977179
transform -1 0 36156 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1768_
timestamp 1649977179
transform 1 0 35696 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1769_
timestamp 1649977179
transform -1 0 35972 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1770_
timestamp 1649977179
transform -1 0 36524 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _1771_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1772_
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1773_
timestamp 1649977179
transform -1 0 9844 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1774_
timestamp 1649977179
transform -1 0 9844 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1775_
timestamp 1649977179
transform 1 0 9292 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1776_
timestamp 1649977179
transform 1 0 6900 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1777_
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1778_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1779_
timestamp 1649977179
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1780_
timestamp 1649977179
transform 1 0 4968 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1781_
timestamp 1649977179
transform -1 0 4968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1782_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1783_
timestamp 1649977179
transform 1 0 5152 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1784_
timestamp 1649977179
transform -1 0 10948 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1785_
timestamp 1649977179
transform 1 0 4968 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1786_
timestamp 1649977179
transform -1 0 3956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1787_
timestamp 1649977179
transform 1 0 11408 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1788_
timestamp 1649977179
transform -1 0 11040 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1789_
timestamp 1649977179
transform 1 0 11960 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1790_
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1791_
timestamp 1649977179
transform 1 0 7268 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1792_
timestamp 1649977179
transform 1 0 7360 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1793_
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1794_
timestamp 1649977179
transform -1 0 11408 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1795_
timestamp 1649977179
transform 1 0 11960 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1796_
timestamp 1649977179
transform 1 0 11592 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1797_
timestamp 1649977179
transform -1 0 16284 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1798_
timestamp 1649977179
transform -1 0 14352 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1799_
timestamp 1649977179
transform 1 0 8096 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1800_
timestamp 1649977179
transform 1 0 9200 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1801_
timestamp 1649977179
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1802_
timestamp 1649977179
transform 1 0 7176 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1803_
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1804_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1805_
timestamp 1649977179
transform 1 0 5244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1806_
timestamp 1649977179
transform 1 0 6716 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1807_
timestamp 1649977179
transform 1 0 5244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1808_
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1809_
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1810_
timestamp 1649977179
transform -1 0 8004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1811_
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1812_
timestamp 1649977179
transform -1 0 4232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1813_
timestamp 1649977179
transform -1 0 5888 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1814_
timestamp 1649977179
transform 1 0 6164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1815_
timestamp 1649977179
transform 1 0 6992 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1816_
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1817_
timestamp 1649977179
transform 1 0 6348 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1818_
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1819_
timestamp 1649977179
transform 1 0 4784 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1820_
timestamp 1649977179
transform -1 0 4692 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1821_
timestamp 1649977179
transform 1 0 10212 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1822_
timestamp 1649977179
transform 1 0 9936 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1823_
timestamp 1649977179
transform 1 0 24932 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1824_
timestamp 1649977179
transform 1 0 32476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1825_
timestamp 1649977179
transform -1 0 34960 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1826_
timestamp 1649977179
transform -1 0 34776 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1827_
timestamp 1649977179
transform -1 0 34224 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1828_
timestamp 1649977179
transform -1 0 34040 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1829_
timestamp 1649977179
transform 1 0 32292 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1830_
timestamp 1649977179
transform -1 0 32568 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1831_
timestamp 1649977179
transform 1 0 29440 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1832_
timestamp 1649977179
transform -1 0 29072 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1833_
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1834_
timestamp 1649977179
transform -1 0 31648 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1835_
timestamp 1649977179
transform -1 0 27692 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1836_
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1837_
timestamp 1649977179
transform 1 0 26036 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1838_
timestamp 1649977179
transform 1 0 27508 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1839_
timestamp 1649977179
transform 1 0 25944 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1840_
timestamp 1649977179
transform 1 0 24748 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1841_
timestamp 1649977179
transform 1 0 24472 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1842_
timestamp 1649977179
transform -1 0 28428 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1843_
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1844_
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1845_
timestamp 1649977179
transform 1 0 24472 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1846_
timestamp 1649977179
transform -1 0 32568 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1847_
timestamp 1649977179
transform -1 0 32384 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _1848_
timestamp 1649977179
transform 1 0 25208 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1849_
timestamp 1649977179
transform 1 0 27048 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1850_
timestamp 1649977179
transform -1 0 31648 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1851_
timestamp 1649977179
transform 1 0 32936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1852_
timestamp 1649977179
transform 1 0 30360 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1853_
timestamp 1649977179
transform -1 0 30636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1854_
timestamp 1649977179
transform -1 0 28152 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1855_
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1856_
timestamp 1649977179
transform -1 0 27784 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1857_
timestamp 1649977179
transform 1 0 27968 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1858_
timestamp 1649977179
transform 1 0 25300 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1859_
timestamp 1649977179
transform 1 0 24656 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1860_
timestamp 1649977179
transform -1 0 24472 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1861_
timestamp 1649977179
transform 1 0 24380 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1862_
timestamp 1649977179
transform -1 0 24840 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1863_
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1864_
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1865_
timestamp 1649977179
transform 1 0 22080 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1866_
timestamp 1649977179
transform 1 0 21896 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1867_
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1868_
timestamp 1649977179
transform 1 0 20976 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1869_
timestamp 1649977179
transform 1 0 23184 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1870_
timestamp 1649977179
transform 1 0 23000 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1871_
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1872_
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _1873_
timestamp 1649977179
transform -1 0 16100 0 1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_2  _1874_
timestamp 1649977179
transform -1 0 14260 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1875_
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1876_
timestamp 1649977179
transform -1 0 12236 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1877_
timestamp 1649977179
transform 1 0 11868 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1878_
timestamp 1649977179
transform -1 0 11040 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1879_
timestamp 1649977179
transform 1 0 10488 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1880_
timestamp 1649977179
transform 1 0 12512 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1881_
timestamp 1649977179
transform -1 0 12144 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1882_
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1883_
timestamp 1649977179
transform 1 0 11960 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1884_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1885_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1886_
timestamp 1649977179
transform -1 0 7912 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1887_
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1888_
timestamp 1649977179
transform 1 0 5244 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1889_
timestamp 1649977179
transform 1 0 5060 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1890_
timestamp 1649977179
transform -1 0 5428 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1891_
timestamp 1649977179
transform -1 0 7452 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1892_
timestamp 1649977179
transform 1 0 6900 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1893_
timestamp 1649977179
transform -1 0 8464 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1894_
timestamp 1649977179
transform 1 0 8188 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1895_
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1896_
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1897_
timestamp 1649977179
transform 1 0 10120 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1898_
timestamp 1649977179
transform 1 0 9660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1899_
timestamp 1649977179
transform 1 0 15640 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1900_
timestamp 1649977179
transform -1 0 14812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1901_
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1902_
timestamp 1649977179
transform -1 0 13616 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1903_
timestamp 1649977179
transform -1 0 15916 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1904_
timestamp 1649977179
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1905_
timestamp 1649977179
transform -1 0 16468 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1906_
timestamp 1649977179
transform -1 0 17112 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1907_
timestamp 1649977179
transform -1 0 15456 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1908_
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1909_
timestamp 1649977179
transform 1 0 13156 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1910_
timestamp 1649977179
transform -1 0 12604 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1911_
timestamp 1649977179
transform -1 0 14628 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1912_
timestamp 1649977179
transform 1 0 10212 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1913_
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1914_
timestamp 1649977179
transform 1 0 15364 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1915_
timestamp 1649977179
transform -1 0 15732 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1916_
timestamp 1649977179
transform 1 0 11776 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1917_
timestamp 1649977179
transform -1 0 11776 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1918_
timestamp 1649977179
transform 1 0 15364 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1919_
timestamp 1649977179
transform 1 0 15272 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1920_
timestamp 1649977179
transform 1 0 13248 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1921_
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1922_
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1923_
timestamp 1649977179
transform 1 0 13340 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _1924_
timestamp 1649977179
transform 1 0 23092 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1925_
timestamp 1649977179
transform -1 0 33948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1926_
timestamp 1649977179
transform -1 0 31372 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1927_
timestamp 1649977179
transform -1 0 31740 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1928_
timestamp 1649977179
transform 1 0 33120 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1929_
timestamp 1649977179
transform -1 0 32844 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1930_
timestamp 1649977179
transform -1 0 33948 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1931_
timestamp 1649977179
transform -1 0 33856 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1932_
timestamp 1649977179
transform 1 0 32936 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1933_
timestamp 1649977179
transform -1 0 33396 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1934_
timestamp 1649977179
transform 1 0 33304 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1935_
timestamp 1649977179
transform 1 0 32568 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1936_
timestamp 1649977179
transform -1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1937_
timestamp 1649977179
transform -1 0 31648 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1938_
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1939_
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1940_
timestamp 1649977179
transform -1 0 31556 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1941_
timestamp 1649977179
transform 1 0 30820 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1942_
timestamp 1649977179
transform 1 0 30636 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1943_
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1944_
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1945_
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1946_
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1947_
timestamp 1649977179
transform -1 0 35972 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1948_
timestamp 1649977179
transform 1 0 36340 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1949_
timestamp 1649977179
transform -1 0 23644 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1950_
timestamp 1649977179
transform 1 0 23184 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1951_
timestamp 1649977179
transform -1 0 25116 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1952_
timestamp 1649977179
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1953_
timestamp 1649977179
transform -1 0 23920 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1954_
timestamp 1649977179
transform -1 0 24012 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1955_
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1956_
timestamp 1649977179
transform -1 0 22724 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1957_
timestamp 1649977179
transform 1 0 21988 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1958_
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1959_
timestamp 1649977179
transform -1 0 25208 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1960_
timestamp 1649977179
transform 1 0 27876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1961_
timestamp 1649977179
transform -1 0 22356 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1962_
timestamp 1649977179
transform -1 0 16836 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1963_
timestamp 1649977179
transform -1 0 16928 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1964_
timestamp 1649977179
transform -1 0 16192 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1965_
timestamp 1649977179
transform 1 0 15640 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1966_
timestamp 1649977179
transform -1 0 15824 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1967_
timestamp 1649977179
transform 1 0 15732 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1968_
timestamp 1649977179
transform 1 0 19872 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1969_
timestamp 1649977179
transform 1 0 18216 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1970_
timestamp 1649977179
transform 1 0 16928 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1971_
timestamp 1649977179
transform -1 0 17388 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1972_
timestamp 1649977179
transform 1 0 22264 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1973_
timestamp 1649977179
transform -1 0 22540 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1974_
timestamp 1649977179
transform -1 0 14536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1975_
timestamp 1649977179
transform 1 0 15640 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _1976_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15456 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1977_
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1978_
timestamp 1649977179
transform -1 0 29716 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1979_
timestamp 1649977179
transform -1 0 29992 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1980_
timestamp 1649977179
transform 1 0 26036 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1981_
timestamp 1649977179
transform -1 0 26036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1982_
timestamp 1649977179
transform -1 0 28060 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1983_
timestamp 1649977179
transform -1 0 27784 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1984_
timestamp 1649977179
transform -1 0 27784 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1985_
timestamp 1649977179
transform 1 0 27968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1986_
timestamp 1649977179
transform -1 0 23736 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1987_
timestamp 1649977179
transform -1 0 23368 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1988_
timestamp 1649977179
transform 1 0 19596 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1989_
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1990_
timestamp 1649977179
transform -1 0 20792 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1991_
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1992_
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1993_
timestamp 1649977179
transform -1 0 21344 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1994_
timestamp 1649977179
transform -1 0 21620 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1995_
timestamp 1649977179
transform -1 0 18768 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1996_
timestamp 1649977179
transform 1 0 18400 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1997_
timestamp 1649977179
transform -1 0 17756 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1998_
timestamp 1649977179
transform -1 0 17572 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1999_
timestamp 1649977179
transform 1 0 17020 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2000_
timestamp 1649977179
transform -1 0 17204 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2001_
timestamp 1649977179
transform -1 0 18124 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2002_
timestamp 1649977179
transform -1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2003_
timestamp 1649977179
transform -1 0 41952 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2004_
timestamp 1649977179
transform 1 0 42412 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2005_
timestamp 1649977179
transform 1 0 42504 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2006_
timestamp 1649977179
transform -1 0 42688 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2007_
timestamp 1649977179
transform 1 0 45816 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2008_
timestamp 1649977179
transform -1 0 45264 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2009_
timestamp 1649977179
transform -1 0 45632 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2010_
timestamp 1649977179
transform 1 0 44252 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2011_
timestamp 1649977179
transform 1 0 41584 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2012_
timestamp 1649977179
transform -1 0 40940 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2013_
timestamp 1649977179
transform -1 0 40480 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2014_
timestamp 1649977179
transform 1 0 44988 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2015_
timestamp 1649977179
transform 1 0 44160 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2016_
timestamp 1649977179
transform -1 0 37352 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2017_
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2018_
timestamp 1649977179
transform 1 0 33764 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2019_
timestamp 1649977179
transform -1 0 37536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2020_
timestamp 1649977179
transform 1 0 45632 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2021_
timestamp 1649977179
transform -1 0 45264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2022_
timestamp 1649977179
transform -1 0 32936 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2023_
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2024_
timestamp 1649977179
transform 1 0 25208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2025_
timestamp 1649977179
transform 1 0 25208 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2026_
timestamp 1649977179
transform -1 0 24656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2027_
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2028_
timestamp 1649977179
transform -1 0 22724 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2029_
timestamp 1649977179
transform -1 0 24656 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2030_
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2031_
timestamp 1649977179
transform -1 0 23000 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2032_
timestamp 1649977179
transform -1 0 19504 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2033_
timestamp 1649977179
transform -1 0 18124 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2034_
timestamp 1649977179
transform 1 0 18400 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _2035_
timestamp 1649977179
transform 1 0 39008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2036_
timestamp 1649977179
transform -1 0 21160 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2037_
timestamp 1649977179
transform 1 0 43424 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2038_
timestamp 1649977179
transform 1 0 31280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2039_
timestamp 1649977179
transform 1 0 29440 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2040_
timestamp 1649977179
transform 1 0 38916 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2041_
timestamp 1649977179
transform -1 0 40296 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2042_
timestamp 1649977179
transform -1 0 38732 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2043_
timestamp 1649977179
transform -1 0 37536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2044_
timestamp 1649977179
transform -1 0 44344 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2045_
timestamp 1649977179
transform 1 0 40388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2046_
timestamp 1649977179
transform 1 0 45632 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2047_
timestamp 1649977179
transform -1 0 45264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2048_
timestamp 1649977179
transform 1 0 46092 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2049_
timestamp 1649977179
transform -1 0 45264 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2050_
timestamp 1649977179
transform 1 0 44252 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2051_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 40572 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2052_
timestamp 1649977179
transform -1 0 40572 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2053_
timestamp 1649977179
transform 1 0 39928 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2054_
timestamp 1649977179
transform -1 0 45356 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _2055_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19044 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2056_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2057_
timestamp 1649977179
transform 1 0 19872 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2058_
timestamp 1649977179
transform 1 0 18584 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2059_
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2060_
timestamp 1649977179
transform 1 0 14720 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2061_
timestamp 1649977179
transform 1 0 14076 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2062_
timestamp 1649977179
transform 1 0 14996 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2063_
timestamp 1649977179
transform 1 0 14444 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2064_
timestamp 1649977179
transform 1 0 15272 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2065_
timestamp 1649977179
transform 1 0 15824 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2066_
timestamp 1649977179
transform 1 0 43608 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2067_
timestamp 1649977179
transform 1 0 43884 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2068_
timestamp 1649977179
transform 1 0 37536 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2069_
timestamp 1649977179
transform 1 0 37904 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2070_
timestamp 1649977179
transform -1 0 39376 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2071_
timestamp 1649977179
transform 1 0 34868 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2072_
timestamp 1649977179
transform -1 0 43884 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2073_
timestamp 1649977179
transform -1 0 43056 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2074_
timestamp 1649977179
transform -1 0 42688 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2075_
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2076_
timestamp 1649977179
transform 1 0 34408 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2077_
timestamp 1649977179
transform 1 0 42412 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2078_
timestamp 1649977179
transform 1 0 43792 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2079_
timestamp 1649977179
transform 1 0 35880 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2080_
timestamp 1649977179
transform 1 0 38456 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2081_
timestamp 1649977179
transform 1 0 30084 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2082_
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2083_
timestamp 1649977179
transform 1 0 36064 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2084_
timestamp 1649977179
transform 1 0 35972 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2085_
timestamp 1649977179
transform 1 0 33856 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2086_
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2087_
timestamp 1649977179
transform -1 0 37628 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2088_
timestamp 1649977179
transform 1 0 9108 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2089_
timestamp 1649977179
transform 1 0 5796 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2090_
timestamp 1649977179
transform 1 0 4784 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2091_
timestamp 1649977179
transform 1 0 4692 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2092_
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2093_
timestamp 1649977179
transform 1 0 4324 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2094_
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2095_
timestamp 1649977179
transform 1 0 10120 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2096_
timestamp 1649977179
transform 1 0 6624 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2097_
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2098_
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2099_
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2100_
timestamp 1649977179
transform 1 0 5336 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2101_
timestamp 1649977179
transform 1 0 5060 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2102_
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2103_
timestamp 1649977179
transform 1 0 5796 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2104_
timestamp 1649977179
transform 1 0 4324 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2105_
timestamp 1649977179
transform -1 0 5796 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2106_
timestamp 1649977179
transform -1 0 6624 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2107_
timestamp 1649977179
transform 1 0 4508 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2108_
timestamp 1649977179
transform 1 0 4416 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2109_
timestamp 1649977179
transform 1 0 9200 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2110_
timestamp 1649977179
transform -1 0 36156 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2111_
timestamp 1649977179
transform -1 0 36156 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2112_
timestamp 1649977179
transform 1 0 32108 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2113_
timestamp 1649977179
transform -1 0 31004 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2114_
timestamp 1649977179
transform 1 0 31464 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2115_
timestamp 1649977179
transform 1 0 25944 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2116_
timestamp 1649977179
transform 1 0 25668 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2117_
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2118_
timestamp 1649977179
transform 1 0 28336 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2119_
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2120_
timestamp 1649977179
transform -1 0 33580 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2121_
timestamp 1649977179
transform -1 0 32660 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2122_
timestamp 1649977179
transform 1 0 30452 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2123_
timestamp 1649977179
transform -1 0 28428 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2124_
timestamp 1649977179
transform -1 0 27600 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2125_
timestamp 1649977179
transform 1 0 24380 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2126_
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2127_
timestamp 1649977179
transform 1 0 20608 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2128_
timestamp 1649977179
transform 1 0 21712 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2129_
timestamp 1649977179
transform 1 0 20608 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2130_
timestamp 1649977179
transform 1 0 22448 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2131_
timestamp 1649977179
transform 1 0 26036 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2132_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2133_
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2134_
timestamp 1649977179
transform 1 0 11868 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2135_
timestamp 1649977179
transform 1 0 11592 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2136_
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2137_
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2138_
timestamp 1649977179
transform 1 0 5244 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2139_
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2140_
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2141_
timestamp 1649977179
transform 1 0 5796 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2142_
timestamp 1649977179
transform 1 0 9200 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2143_
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2144_
timestamp 1649977179
transform -1 0 16100 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2145_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2146_
timestamp 1649977179
transform -1 0 15824 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2147_
timestamp 1649977179
transform -1 0 12880 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2148_
timestamp 1649977179
transform 1 0 5060 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2149_
timestamp 1649977179
transform 1 0 15272 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2150_
timestamp 1649977179
transform -1 0 12236 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2151_
timestamp 1649977179
transform 1 0 14996 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2152_
timestamp 1649977179
transform 1 0 11960 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2153_
timestamp 1649977179
transform 1 0 12144 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2154_
timestamp 1649977179
transform -1 0 33212 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2155_
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2156_
timestamp 1649977179
transform -1 0 36524 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2157_
timestamp 1649977179
transform 1 0 33120 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2158_
timestamp 1649977179
transform 1 0 32200 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2159_
timestamp 1649977179
transform -1 0 31648 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2160_
timestamp 1649977179
transform 1 0 31924 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2161_
timestamp 1649977179
transform 1 0 30452 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2162_
timestamp 1649977179
transform 1 0 31188 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2163_
timestamp 1649977179
transform 1 0 28244 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2164_
timestamp 1649977179
transform 1 0 36064 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2165_
timestamp 1649977179
transform 1 0 24656 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2166_
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2167_
timestamp 1649977179
transform 1 0 22448 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2168_
timestamp 1649977179
transform 1 0 21528 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2169_
timestamp 1649977179
transform -1 0 26496 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2170_
timestamp 1649977179
transform -1 0 18032 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2171_
timestamp 1649977179
transform 1 0 15364 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2172_
timestamp 1649977179
transform 1 0 13892 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2173_
timestamp 1649977179
transform 1 0 18032 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2174_
timestamp 1649977179
transform 1 0 17204 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2175_
timestamp 1649977179
transform 1 0 22172 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2176_
timestamp 1649977179
transform 1 0 30176 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2177_
timestamp 1649977179
transform 1 0 26404 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2178_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 27508 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2179_
timestamp 1649977179
transform -1 0 27600 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2180_
timestamp 1649977179
transform -1 0 26312 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2181_
timestamp 1649977179
transform 1 0 21160 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2182_
timestamp 1649977179
transform -1 0 19780 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _2183_
timestamp 1649977179
transform 1 0 22356 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2184_
timestamp 1649977179
transform 1 0 17296 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _2185_
timestamp 1649977179
transform 1 0 18124 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _2186_
timestamp 1649977179
transform 1 0 17020 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _2187_
timestamp 1649977179
transform 1 0 19228 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _2188_
timestamp 1649977179
transform 1 0 40572 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2189_
timestamp 1649977179
transform 1 0 40480 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _2190_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 40204 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2191_
timestamp 1649977179
transform 1 0 39744 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _2192_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 42688 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__dfrtp_1  _2193_
timestamp 1649977179
transform 1 0 43700 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2194_
timestamp 1649977179
transform 1 0 43608 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _2195_
timestamp 1649977179
transform 1 0 43424 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2196_
timestamp 1649977179
transform 1 0 43424 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _2197_
timestamp 1649977179
transform 1 0 44988 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__dfrtp_1  _2198_
timestamp 1649977179
transform 1 0 43884 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2199_
timestamp 1649977179
transform 1 0 43884 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _2200_
timestamp 1649977179
transform -1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2201_
timestamp 1649977179
transform -1 0 44988 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_4  _2202_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 45724 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxtn_2  _2203_
timestamp 1649977179
transform 1 0 47564 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__dfrtp_1  _2204_
timestamp 1649977179
transform -1 0 41676 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2205_
timestamp 1649977179
transform 1 0 37996 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _2206_
timestamp 1649977179
transform 1 0 37536 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2207_
timestamp 1649977179
transform 1 0 36984 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _2208_
timestamp 1649977179
transform 1 0 38180 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__dfrtp_1  _2209_
timestamp 1649977179
transform 1 0 43608 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2210_
timestamp 1649977179
transform 1 0 43332 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _2211_
timestamp 1649977179
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2212_
timestamp 1649977179
transform 1 0 42780 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2213_
timestamp 1649977179
transform 1 0 45816 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _2214_
timestamp 1649977179
transform -1 0 37260 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2215_
timestamp 1649977179
transform 1 0 33028 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _2216_
timestamp 1649977179
transform 1 0 35052 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2217_
timestamp 1649977179
transform -1 0 34776 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2218_
timestamp 1649977179
transform 1 0 35696 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _2219_
timestamp 1649977179
transform 1 0 35972 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2220_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 43884 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2221_
timestamp 1649977179
transform 1 0 43700 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtp_1  _2222_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 51796 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _2223_
timestamp 1649977179
transform 1 0 31004 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2224_
timestamp 1649977179
transform 1 0 23828 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2225_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22724 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2226_
timestamp 1649977179
transform 1 0 23000 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2227_
timestamp 1649977179
transform 1 0 22632 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2228_
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2229_
timestamp 1649977179
transform 1 0 20792 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2230_
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2231_
timestamp 1649977179
transform 1 0 17848 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2232_
timestamp 1649977179
transform 1 0 15364 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2233_
timestamp 1649977179
transform 1 0 17480 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2234_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2235_
timestamp 1649977179
transform -1 0 45356 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2236_
timestamp 1649977179
transform 1 0 30728 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2237_
timestamp 1649977179
transform 1 0 29072 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2238_
timestamp 1649977179
transform -1 0 40112 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2239_
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2240_
timestamp 1649977179
transform 1 0 35512 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2241_
timestamp 1649977179
transform -1 0 45264 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2242_
timestamp 1649977179
transform 1 0 39836 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2243_
timestamp 1649977179
transform 1 0 42688 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2244_
timestamp 1649977179
transform 1 0 43608 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2245_
timestamp 1649977179
transform 1 0 43884 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2246_
timestamp 1649977179
transform 1 0 43792 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2247_
timestamp 1649977179
transform 1 0 44988 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_1  _2248_
timestamp 1649977179
transform -1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2249_
timestamp 1649977179
transform -1 0 50140 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2250_
timestamp 1649977179
transform -1 0 50048 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2251_
timestamp 1649977179
transform -1 0 48668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _2252_
timestamp 1649977179
transform -1 0 50232 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _2253_
timestamp 1649977179
transform -1 0 49680 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _2254_
timestamp 1649977179
transform -1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  _2470_
timestamp 1649977179
transform -1 0 52992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2471_
timestamp 1649977179
transform -1 0 55568 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2472_
timestamp 1649977179
transform -1 0 60812 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2473_
timestamp 1649977179
transform -1 0 67436 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2474_
timestamp 1649977179
transform -1 0 57960 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2475_
timestamp 1649977179
transform -1 0 67436 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2476_
timestamp 1649977179
transform -1 0 67436 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2477_
timestamp 1649977179
transform -1 0 67436 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _2478_
timestamp 1649977179
transform -1 0 67436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24840 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12328 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1649977179
transform -1 0 12880 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1649977179
transform 1 0 17204 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1649977179
transform 1 0 17296 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1649977179
transform 1 0 12328 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1649977179
transform -1 0 13432 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1649977179
transform 1 0 19412 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1649977179
transform -1 0 19136 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1649977179
transform -1 0 34316 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1649977179
transform 1 0 32108 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1649977179
transform 1 0 38180 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1649977179
transform 1 0 38732 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1649977179
transform 1 0 32660 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1649977179
transform -1 0 34224 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1649977179
transform 1 0 38088 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1649977179
transform 1 0 37904 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1649977179
transform -1 0 56396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1649977179
transform -1 0 46828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 49312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 50140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 47196 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 48484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1649977179
transform -1 0 48300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input9 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12512 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 11684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 12328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 12972 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 10396 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 12788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 11776 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1649977179
transform -1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 12328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 12512 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform 1 0 13800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1649977179
transform -1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform 1 0 14536 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1649977179
transform -1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input32
timestamp 1649977179
transform -1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1649977179
transform -1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1649977179
transform 1 0 15824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 12696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1649977179
transform -1 0 51336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform -1 0 51888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform -1 0 53084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform 1 0 52716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1649977179
transform 1 0 53452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1649977179
transform -1 0 53820 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1649977179
transform -1 0 54556 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1649977179
transform -1 0 54556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1649977179
transform -1 0 55660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 54372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform -1 0 55292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform -1 0 40296 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform -1 0 41032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform -1 0 41768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 43148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform 1 0 43884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform -1 0 43608 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 43976 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform -1 0 46092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform -1 0 46092 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 67804 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 67804 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform 1 0 67804 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 67804 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 67344 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 67344 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 67344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 67344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater71
timestamp 1649977179
transform -1 0 50876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_72 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4600 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_73
timestamp 1649977179
transform 1 0 5612 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_74
timestamp 1649977179
transform -1 0 7820 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_75
timestamp 1649977179
transform -1 0 9568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_76
timestamp 1649977179
transform 1 0 10764 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_77
timestamp 1649977179
transform -1 0 12880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_78
timestamp 1649977179
transform -1 0 14536 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_79
timestamp 1649977179
transform -1 0 16192 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_80
timestamp 1649977179
transform -1 0 17848 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_81
timestamp 1649977179
transform -1 0 19504 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_82
timestamp 1649977179
transform -1 0 21252 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_83
timestamp 1649977179
transform -1 0 22816 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_84
timestamp 1649977179
transform -1 0 24656 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_85
timestamp 1649977179
transform 1 0 25576 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_86
timestamp 1649977179
transform -1 0 27784 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_87
timestamp 1649977179
transform 1 0 28796 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_88
timestamp 1649977179
transform -1 0 31004 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_89
timestamp 1649977179
transform -1 0 32752 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_90
timestamp 1649977179
transform 1 0 33948 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_91
timestamp 1649977179
transform -1 0 36156 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_92
timestamp 1649977179
transform -1 0 37812 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_93
timestamp 1649977179
transform -1 0 40112 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_94
timestamp 1649977179
transform -1 0 41400 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_95
timestamp 1649977179
transform -1 0 42780 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_96
timestamp 1649977179
transform -1 0 44436 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_97
timestamp 1649977179
transform -1 0 46092 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_98
timestamp 1649977179
transform -1 0 47840 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_99
timestamp 1649977179
transform -1 0 49404 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_100
timestamp 1649977179
transform -1 0 51060 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_101
timestamp 1649977179
transform -1 0 52992 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_102
timestamp 1649977179
transform -1 0 54372 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_103
timestamp 1649977179
transform -1 0 56212 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_104
timestamp 1649977179
transform -1 0 58144 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_105
timestamp 1649977179
transform -1 0 59432 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_106
timestamp 1649977179
transform -1 0 61364 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_107
timestamp 1649977179
transform -1 0 63296 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_108
timestamp 1649977179
transform -1 0 64584 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_109
timestamp 1649977179
transform -1 0 65964 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_110
timestamp 1649977179
transform -1 0 5244 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_111
timestamp 1649977179
transform -1 0 6900 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_112
timestamp 1649977179
transform -1 0 8464 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_113
timestamp 1649977179
transform -1 0 10212 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_114
timestamp 1649977179
transform -1 0 11868 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_115
timestamp 1649977179
transform -1 0 13524 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_116
timestamp 1649977179
transform -1 0 15180 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_117
timestamp 1649977179
transform -1 0 16928 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_118
timestamp 1649977179
transform -1 0 18492 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_119
timestamp 1649977179
transform -1 0 20148 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_120
timestamp 1649977179
transform -1 0 22080 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_121
timestamp 1649977179
transform -1 0 23460 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_122
timestamp 1649977179
transform -1 0 25116 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_123
timestamp 1649977179
transform 1 0 26220 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_124
timestamp 1649977179
transform -1 0 28428 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_125
timestamp 1649977179
transform -1 0 30084 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_126
timestamp 1649977179
transform -1 0 31648 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_127
timestamp 1649977179
transform -1 0 33396 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_128
timestamp 1649977179
transform -1 0 35052 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_129
timestamp 1649977179
transform -1 0 36800 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_130
timestamp 1649977179
transform -1 0 38456 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_131
timestamp 1649977179
transform -1 0 40756 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_132
timestamp 1649977179
transform -1 0 41676 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_133
timestamp 1649977179
transform -1 0 43424 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_134
timestamp 1649977179
transform -1 0 45264 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_135
timestamp 1649977179
transform -1 0 46736 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_136
timestamp 1649977179
transform -1 0 48484 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_137
timestamp 1649977179
transform -1 0 50416 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_138
timestamp 1649977179
transform -1 0 51704 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_139
timestamp 1649977179
transform -1 0 53636 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_140
timestamp 1649977179
transform -1 0 55568 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_141
timestamp 1649977179
transform -1 0 56856 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_142
timestamp 1649977179
transform -1 0 58788 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_143
timestamp 1649977179
transform -1 0 60720 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_144
timestamp 1649977179
transform -1 0 62008 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_145
timestamp 1649977179
transform -1 0 63940 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_146
timestamp 1649977179
transform -1 0 64860 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_147
timestamp 1649977179
transform -1 0 66608 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_148
timestamp 1649977179
transform -1 0 59432 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_149
timestamp 1649977179
transform -1 0 58788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_150
timestamp 1649977179
transform -1 0 58788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_151
timestamp 1649977179
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_152
timestamp 1649977179
transform -1 0 22632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_153
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_154
timestamp 1649977179
transform -1 0 23368 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_155
timestamp 1649977179
transform 1 0 22356 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_156
timestamp 1649977179
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_157
timestamp 1649977179
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_158
timestamp 1649977179
transform 1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_159
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_160
timestamp 1649977179
transform 1 0 23000 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_161
timestamp 1649977179
transform 1 0 23644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_162
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_163
timestamp 1649977179
transform 1 0 24288 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_164
timestamp 1649977179
transform 1 0 24932 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_165
timestamp 1649977179
transform -1 0 26496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_166
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_167
timestamp 1649977179
transform 1 0 24932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_168
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_169
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_170
timestamp 1649977179
transform 1 0 26864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_171
timestamp 1649977179
transform -1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_172
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_173
timestamp 1649977179
transform 1 0 27508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_174
timestamp 1649977179
transform 1 0 27140 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_175
timestamp 1649977179
transform 1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_176
timestamp 1649977179
transform 1 0 28796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_177
timestamp 1649977179
transform 1 0 27784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_178
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_179
timestamp 1649977179
transform -1 0 30268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_180
timestamp 1649977179
transform 1 0 27508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_181
timestamp 1649977179
transform 1 0 28428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_182
timestamp 1649977179
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_183
timestamp 1649977179
transform -1 0 31372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_184
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_185
timestamp 1649977179
transform 1 0 30084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_186
timestamp 1649977179
transform -1 0 32200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_187
timestamp 1649977179
transform -1 0 34224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_188
timestamp 1649977179
transform 1 0 30084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_189
timestamp 1649977179
transform 1 0 30728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_190
timestamp 1649977179
transform 1 0 31372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_191
timestamp 1649977179
transform -1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_192
timestamp 1649977179
transform 1 0 32660 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_193
timestamp 1649977179
transform 1 0 33580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_194
timestamp 1649977179
transform 1 0 33304 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_195
timestamp 1649977179
transform -1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_196
timestamp 1649977179
transform 1 0 33948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_197
timestamp 1649977179
transform -1 0 35144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_198
timestamp 1649977179
transform 1 0 34776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_199
timestamp 1649977179
transform -1 0 35788 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_200
timestamp 1649977179
transform 1 0 35420 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_201
timestamp 1649977179
transform -1 0 36340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_202
timestamp 1649977179
transform -1 0 36616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_203
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_204
timestamp 1649977179
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_205
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_206
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_207
timestamp 1649977179
transform -1 0 38180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_208
timestamp 1649977179
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_209
timestamp 1649977179
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_210
timestamp 1649977179
transform -1 0 39468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_211
timestamp 1649977179
transform -1 0 39100 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_212
timestamp 1649977179
transform 1 0 38180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_213
timestamp 1649977179
transform 1 0 39100 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_214
timestamp 1649977179
transform 1 0 35328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_215
timestamp 1649977179
transform -1 0 46736 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_216
timestamp 1649977179
transform -1 0 46460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_217
timestamp 1649977179
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_218
timestamp 1649977179
transform -1 0 48944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_219
timestamp 1649977179
transform -1 0 48484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_220
timestamp 1649977179
transform -1 0 45908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_221
timestamp 1649977179
transform -1 0 48116 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_222
timestamp 1649977179
transform -1 0 46552 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_223
timestamp 1649977179
transform -1 0 46000 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_224
timestamp 1649977179
transform -1 0 46644 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_225
timestamp 1649977179
transform -1 0 47840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_226
timestamp 1649977179
transform -1 0 46828 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_227
timestamp 1649977179
transform -1 0 47840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_228
timestamp 1649977179
transform -1 0 49128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_229
timestamp 1649977179
transform -1 0 48484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_230
timestamp 1649977179
transform -1 0 50416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_231
timestamp 1649977179
transform -1 0 51336 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_232
timestamp 1649977179
transform -1 0 51060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_233
timestamp 1649977179
transform -1 0 52440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_234
timestamp 1649977179
transform -1 0 50784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_235
timestamp 1649977179
transform -1 0 53084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_236
timestamp 1649977179
transform -1 0 52992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_237
timestamp 1649977179
transform -1 0 52072 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_238
timestamp 1649977179
transform -1 0 53636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_239
timestamp 1649977179
transform -1 0 52992 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_240
timestamp 1649977179
transform -1 0 54280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_241
timestamp 1649977179
transform -1 0 53636 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_242
timestamp 1649977179
transform -1 0 55936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_243
timestamp 1649977179
transform -1 0 55568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_244
timestamp 1649977179
transform -1 0 57040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_245
timestamp 1649977179
transform -1 0 56580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_246
timestamp 1649977179
transform -1 0 56212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_247
timestamp 1649977179
transform -1 0 57224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_248
timestamp 1649977179
transform -1 0 56856 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_249
timestamp 1649977179
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_250
timestamp 1649977179
transform -1 0 57500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_251
timestamp 1649977179
transform -1 0 58788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_252
timestamp 1649977179
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_253
timestamp 1649977179
transform -1 0 58144 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_254
timestamp 1649977179
transform 1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_255
timestamp 1649977179
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_256
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_257
timestamp 1649977179
transform 1 0 13064 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_258
timestamp 1649977179
transform 1 0 10764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_259
timestamp 1649977179
transform 1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_260
timestamp 1649977179
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_261
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_262
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_263
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_264
timestamp 1649977179
transform 1 0 14352 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_265
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_266
timestamp 1649977179
transform -1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_267
timestamp 1649977179
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_268
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_269
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_270
timestamp 1649977179
transform 1 0 17204 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_271
timestamp 1649977179
transform 1 0 17112 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_272
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_273
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_274
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_275
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_276
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_277
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_278
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_279
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_280
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_281
timestamp 1649977179
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_282
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_283
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_284
timestamp 1649977179
transform 1 0 20424 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_285
timestamp 1649977179
transform -1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_286
timestamp 1649977179
transform 1 0 21712 0 1 3264
box -38 -48 314 592
<< labels >>
flabel metal2 s 3790 59200 3846 60000 0 FreeSans 224 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 20350 59200 20406 60000 0 FreeSans 224 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 22006 59200 22062 60000 0 FreeSans 224 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 23662 59200 23718 60000 0 FreeSans 224 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 25318 59200 25374 60000 0 FreeSans 224 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 26974 59200 27030 60000 0 FreeSans 224 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 28630 59200 28686 60000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 30286 59200 30342 60000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 31942 59200 31998 60000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 33598 59200 33654 60000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 35254 59200 35310 60000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 5446 59200 5502 60000 0 FreeSans 224 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 36910 59200 36966 60000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 38566 59200 38622 60000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 40222 59200 40278 60000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 41878 59200 41934 60000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 43534 59200 43590 60000 0 FreeSans 224 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 45190 59200 45246 60000 0 FreeSans 224 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 46846 59200 46902 60000 0 FreeSans 224 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 48502 59200 48558 60000 0 FreeSans 224 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 50158 59200 50214 60000 0 FreeSans 224 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 51814 59200 51870 60000 0 FreeSans 224 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 7102 59200 7158 60000 0 FreeSans 224 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 53470 59200 53526 60000 0 FreeSans 224 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 55126 59200 55182 60000 0 FreeSans 224 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 56782 59200 56838 60000 0 FreeSans 224 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 58438 59200 58494 60000 0 FreeSans 224 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 60094 59200 60150 60000 0 FreeSans 224 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 61750 59200 61806 60000 0 FreeSans 224 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 63406 59200 63462 60000 0 FreeSans 224 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 65062 59200 65118 60000 0 FreeSans 224 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 8758 59200 8814 60000 0 FreeSans 224 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 10414 59200 10470 60000 0 FreeSans 224 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 12070 59200 12126 60000 0 FreeSans 224 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 13726 59200 13782 60000 0 FreeSans 224 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 15382 59200 15438 60000 0 FreeSans 224 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 17038 59200 17094 60000 0 FreeSans 224 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 18694 59200 18750 60000 0 FreeSans 224 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 4342 59200 4398 60000 0 FreeSans 224 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 20902 59200 20958 60000 0 FreeSans 224 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 22558 59200 22614 60000 0 FreeSans 224 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 24214 59200 24270 60000 0 FreeSans 224 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 25870 59200 25926 60000 0 FreeSans 224 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 27526 59200 27582 60000 0 FreeSans 224 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 29182 59200 29238 60000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 30838 59200 30894 60000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 32494 59200 32550 60000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 34150 59200 34206 60000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 35806 59200 35862 60000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 5998 59200 6054 60000 0 FreeSans 224 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 37462 59200 37518 60000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 39118 59200 39174 60000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 40774 59200 40830 60000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 42430 59200 42486 60000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 44086 59200 44142 60000 0 FreeSans 224 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 45742 59200 45798 60000 0 FreeSans 224 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 47398 59200 47454 60000 0 FreeSans 224 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 49054 59200 49110 60000 0 FreeSans 224 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 50710 59200 50766 60000 0 FreeSans 224 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 52366 59200 52422 60000 0 FreeSans 224 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 7654 59200 7710 60000 0 FreeSans 224 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 54022 59200 54078 60000 0 FreeSans 224 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 55678 59200 55734 60000 0 FreeSans 224 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 57334 59200 57390 60000 0 FreeSans 224 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 58990 59200 59046 60000 0 FreeSans 224 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 60646 59200 60702 60000 0 FreeSans 224 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 62302 59200 62358 60000 0 FreeSans 224 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 63958 59200 64014 60000 0 FreeSans 224 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 65614 59200 65670 60000 0 FreeSans 224 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 9310 59200 9366 60000 0 FreeSans 224 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 10966 59200 11022 60000 0 FreeSans 224 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 12622 59200 12678 60000 0 FreeSans 224 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 14278 59200 14334 60000 0 FreeSans 224 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 15934 59200 15990 60000 0 FreeSans 224 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 17590 59200 17646 60000 0 FreeSans 224 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 19246 59200 19302 60000 0 FreeSans 224 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 4894 59200 4950 60000 0 FreeSans 224 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 21454 59200 21510 60000 0 FreeSans 224 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 23110 59200 23166 60000 0 FreeSans 224 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 24766 59200 24822 60000 0 FreeSans 224 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 26422 59200 26478 60000 0 FreeSans 224 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 28078 59200 28134 60000 0 FreeSans 224 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 29734 59200 29790 60000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 31390 59200 31446 60000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 33046 59200 33102 60000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 34702 59200 34758 60000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 36358 59200 36414 60000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 6550 59200 6606 60000 0 FreeSans 224 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 38014 59200 38070 60000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 39670 59200 39726 60000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 41326 59200 41382 60000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 42982 59200 43038 60000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 44638 59200 44694 60000 0 FreeSans 224 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 46294 59200 46350 60000 0 FreeSans 224 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 47950 59200 48006 60000 0 FreeSans 224 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 49606 59200 49662 60000 0 FreeSans 224 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 51262 59200 51318 60000 0 FreeSans 224 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 52918 59200 52974 60000 0 FreeSans 224 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 8206 59200 8262 60000 0 FreeSans 224 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 54574 59200 54630 60000 0 FreeSans 224 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 56230 59200 56286 60000 0 FreeSans 224 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 57886 59200 57942 60000 0 FreeSans 224 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 59542 59200 59598 60000 0 FreeSans 224 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 61198 59200 61254 60000 0 FreeSans 224 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 62854 59200 62910 60000 0 FreeSans 224 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 64510 59200 64566 60000 0 FreeSans 224 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 66166 59200 66222 60000 0 FreeSans 224 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 9862 59200 9918 60000 0 FreeSans 224 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 11518 59200 11574 60000 0 FreeSans 224 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 13174 59200 13230 60000 0 FreeSans 224 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 14830 59200 14886 60000 0 FreeSans 224 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 16486 59200 16542 60000 0 FreeSans 224 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 18142 59200 18198 60000 0 FreeSans 224 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 19798 59200 19854 60000 0 FreeSans 224 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 57426 0 57482 800 0 FreeSans 224 90 0 0 irq[0]
port 114 nsew signal tristate
flabel metal2 s 57518 0 57574 800 0 FreeSans 224 90 0 0 irq[1]
port 115 nsew signal tristate
flabel metal2 s 57610 0 57666 800 0 FreeSans 224 90 0 0 irq[2]
port 116 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 117 nsew signal input
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 118 nsew signal input
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 119 nsew signal input
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 120 nsew signal input
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 121 nsew signal input
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 122 nsew signal input
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 123 nsew signal input
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 124 nsew signal input
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 125 nsew signal input
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 126 nsew signal input
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 127 nsew signal input
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 128 nsew signal input
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 129 nsew signal input
flabel metal2 s 52734 0 52790 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 130 nsew signal input
flabel metal2 s 53010 0 53066 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 131 nsew signal input
flabel metal2 s 53286 0 53342 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 132 nsew signal input
flabel metal2 s 53562 0 53618 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 133 nsew signal input
flabel metal2 s 53838 0 53894 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 134 nsew signal input
flabel metal2 s 54114 0 54170 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 135 nsew signal input
flabel metal2 s 54390 0 54446 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 136 nsew signal input
flabel metal2 s 54666 0 54722 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 137 nsew signal input
flabel metal2 s 54942 0 54998 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 138 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 139 nsew signal input
flabel metal2 s 55218 0 55274 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 140 nsew signal input
flabel metal2 s 55494 0 55550 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 141 nsew signal input
flabel metal2 s 55770 0 55826 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 142 nsew signal input
flabel metal2 s 56046 0 56102 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 143 nsew signal input
flabel metal2 s 56322 0 56378 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 144 nsew signal input
flabel metal2 s 56598 0 56654 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 145 nsew signal input
flabel metal2 s 56874 0 56930 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 146 nsew signal input
flabel metal2 s 57150 0 57206 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 147 nsew signal input
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 148 nsew signal input
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 149 nsew signal input
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 150 nsew signal input
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 151 nsew signal input
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 152 nsew signal input
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 153 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 154 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 155 nsew signal input
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 156 nsew signal input
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 157 nsew signal input
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 158 nsew signal input
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 159 nsew signal input
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 160 nsew signal input
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 161 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 162 nsew signal input
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 163 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 164 nsew signal input
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 165 nsew signal input
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 166 nsew signal input
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 167 nsew signal input
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 168 nsew signal input
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 169 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 170 nsew signal input
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 171 nsew signal input
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 172 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 173 nsew signal input
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 174 nsew signal input
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 175 nsew signal input
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 176 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 177 nsew signal input
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 178 nsew signal input
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 179 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 180 nsew signal input
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 181 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 182 nsew signal input
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 183 nsew signal input
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 184 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 185 nsew signal input
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 186 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 187 nsew signal input
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 188 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 189 nsew signal input
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 190 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 191 nsew signal input
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 192 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 193 nsew signal input
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 194 nsew signal input
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 195 nsew signal input
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 196 nsew signal input
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 197 nsew signal input
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 198 nsew signal input
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 199 nsew signal input
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 200 nsew signal input
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 201 nsew signal input
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 202 nsew signal input
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 203 nsew signal input
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 204 nsew signal input
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 205 nsew signal input
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 206 nsew signal input
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 207 nsew signal input
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 208 nsew signal input
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 209 nsew signal input
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 210 nsew signal input
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 211 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 212 nsew signal input
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 213 nsew signal input
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 214 nsew signal input
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 215 nsew signal input
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 216 nsew signal input
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 217 nsew signal input
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 218 nsew signal input
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 219 nsew signal input
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 220 nsew signal input
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 221 nsew signal input
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 222 nsew signal input
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 223 nsew signal input
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 224 nsew signal input
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 225 nsew signal input
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 226 nsew signal input
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 227 nsew signal input
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 228 nsew signal input
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 229 nsew signal input
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 230 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 231 nsew signal input
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 232 nsew signal input
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 233 nsew signal input
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 234 nsew signal input
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 235 nsew signal input
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 236 nsew signal input
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 237 nsew signal input
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 238 nsew signal input
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 239 nsew signal input
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 240 nsew signal input
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 241 nsew signal input
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 242 nsew signal input
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 243 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 244 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 245 nsew signal tristate
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 246 nsew signal tristate
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 247 nsew signal tristate
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 248 nsew signal tristate
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 249 nsew signal tristate
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 250 nsew signal tristate
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 251 nsew signal tristate
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 252 nsew signal tristate
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 253 nsew signal tristate
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 254 nsew signal tristate
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 255 nsew signal tristate
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 256 nsew signal tristate
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 257 nsew signal tristate
flabel metal2 s 52826 0 52882 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 258 nsew signal tristate
flabel metal2 s 53102 0 53158 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 259 nsew signal tristate
flabel metal2 s 53378 0 53434 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 260 nsew signal tristate
flabel metal2 s 53654 0 53710 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 261 nsew signal tristate
flabel metal2 s 53930 0 53986 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 262 nsew signal tristate
flabel metal2 s 54206 0 54262 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 263 nsew signal tristate
flabel metal2 s 54482 0 54538 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 264 nsew signal tristate
flabel metal2 s 54758 0 54814 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 265 nsew signal tristate
flabel metal2 s 55034 0 55090 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 266 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 267 nsew signal tristate
flabel metal2 s 55310 0 55366 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 268 nsew signal tristate
flabel metal2 s 55586 0 55642 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 269 nsew signal tristate
flabel metal2 s 55862 0 55918 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 270 nsew signal tristate
flabel metal2 s 56138 0 56194 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 271 nsew signal tristate
flabel metal2 s 56414 0 56470 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 272 nsew signal tristate
flabel metal2 s 56690 0 56746 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 273 nsew signal tristate
flabel metal2 s 56966 0 57022 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 274 nsew signal tristate
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 275 nsew signal tristate
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 276 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 277 nsew signal tristate
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 278 nsew signal tristate
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 279 nsew signal tristate
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 280 nsew signal tristate
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 281 nsew signal tristate
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 282 nsew signal tristate
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 283 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 284 nsew signal tristate
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 285 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 286 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 287 nsew signal tristate
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 288 nsew signal tristate
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 289 nsew signal tristate
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 290 nsew signal tristate
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 291 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 292 nsew signal tristate
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 293 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 294 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 295 nsew signal tristate
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 296 nsew signal tristate
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 297 nsew signal tristate
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 298 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 299 nsew signal tristate
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 300 nsew signal tristate
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 301 nsew signal tristate
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 302 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 303 nsew signal tristate
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 304 nsew signal tristate
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 305 nsew signal tristate
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 306 nsew signal tristate
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 307 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 308 nsew signal tristate
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 309 nsew signal tristate
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 310 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 311 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 312 nsew signal tristate
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 313 nsew signal tristate
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 314 nsew signal tristate
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 315 nsew signal tristate
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 316 nsew signal tristate
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 317 nsew signal tristate
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 318 nsew signal tristate
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 319 nsew signal tristate
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 320 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 321 nsew signal tristate
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 322 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 323 nsew signal tristate
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 324 nsew signal tristate
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 325 nsew signal tristate
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 326 nsew signal tristate
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 327 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 328 nsew signal tristate
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 329 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 330 nsew signal tristate
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 331 nsew signal tristate
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 332 nsew signal tristate
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 333 nsew signal tristate
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 334 nsew signal tristate
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 335 nsew signal tristate
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 336 nsew signal tristate
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 337 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 338 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 339 nsew signal tristate
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 340 nsew signal tristate
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 341 nsew signal tristate
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 342 nsew signal tristate
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 343 nsew signal tristate
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 344 nsew signal tristate
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 345 nsew signal tristate
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 346 nsew signal tristate
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 347 nsew signal tristate
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 348 nsew signal tristate
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 349 nsew signal tristate
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 350 nsew signal tristate
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 351 nsew signal tristate
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 352 nsew signal tristate
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 353 nsew signal tristate
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 354 nsew signal tristate
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 355 nsew signal tristate
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 356 nsew signal tristate
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 357 nsew signal tristate
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 358 nsew signal tristate
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 359 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 360 nsew signal tristate
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 361 nsew signal tristate
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 362 nsew signal tristate
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 363 nsew signal tristate
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 364 nsew signal tristate
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 365 nsew signal tristate
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 366 nsew signal tristate
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 367 nsew signal tristate
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 368 nsew signal tristate
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 369 nsew signal tristate
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 370 nsew signal tristate
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 371 nsew signal tristate
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 372 nsew signal tristate
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 373 nsew signal input
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 374 nsew signal input
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 375 nsew signal input
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 376 nsew signal input
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 377 nsew signal input
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 378 nsew signal input
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 379 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 380 nsew signal input
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 381 nsew signal input
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 382 nsew signal input
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 383 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 384 nsew signal input
flabel metal2 s 52642 0 52698 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 385 nsew signal input
flabel metal2 s 52918 0 52974 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 386 nsew signal input
flabel metal2 s 53194 0 53250 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 387 nsew signal input
flabel metal2 s 53470 0 53526 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 388 nsew signal input
flabel metal2 s 53746 0 53802 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 389 nsew signal input
flabel metal2 s 54022 0 54078 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 390 nsew signal input
flabel metal2 s 54298 0 54354 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 391 nsew signal input
flabel metal2 s 54574 0 54630 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 392 nsew signal input
flabel metal2 s 54850 0 54906 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 393 nsew signal input
flabel metal2 s 55126 0 55182 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 394 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 395 nsew signal input
flabel metal2 s 55402 0 55458 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 396 nsew signal input
flabel metal2 s 55678 0 55734 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 397 nsew signal input
flabel metal2 s 55954 0 56010 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 398 nsew signal input
flabel metal2 s 56230 0 56286 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 399 nsew signal input
flabel metal2 s 56506 0 56562 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 400 nsew signal input
flabel metal2 s 56782 0 56838 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 401 nsew signal input
flabel metal2 s 57058 0 57114 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 402 nsew signal input
flabel metal2 s 57334 0 57390 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 403 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 404 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 405 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 406 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 407 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 408 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 409 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 410 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 411 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 412 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 413 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 414 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 415 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 416 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 417 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 418 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 419 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 420 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 421 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 422 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 423 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 424 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 425 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 426 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 427 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 428 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 429 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 430 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 431 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 432 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 433 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 434 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 435 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 436 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 437 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 438 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 439 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 440 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 441 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 442 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 443 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 444 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 445 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 446 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 447 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 448 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 449 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 450 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 451 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 452 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 453 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 454 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 455 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 456 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 457 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 458 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 459 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 460 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 461 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 462 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 463 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 464 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 465 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 466 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 467 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 468 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 469 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 470 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 471 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 472 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 473 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 474 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 475 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 476 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 477 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 478 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 479 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 480 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 481 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 482 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 483 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 484 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 485 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 486 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 487 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 488 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 489 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 490 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 491 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 492 nsew signal input
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 493 nsew signal input
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 494 nsew signal input
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 495 nsew signal input
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 496 nsew signal input
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 497 nsew signal input
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 498 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 499 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 500 nsew signal input
flabel metal3 s 69200 18640 70000 18760 0 FreeSans 480 0 0 0 out_1
port 501 nsew signal tristate
flabel metal3 s 69200 26120 70000 26240 0 FreeSans 480 0 0 0 out_2
port 502 nsew signal tristate
flabel metal3 s 69200 33600 70000 33720 0 FreeSans 480 0 0 0 out_3
port 503 nsew signal tristate
flabel metal3 s 69200 41080 70000 41200 0 FreeSans 480 0 0 0 out_4
port 504 nsew signal tristate
flabel metal3 s 69200 48560 70000 48680 0 FreeSans 480 0 0 0 out_5
port 505 nsew signal tristate
flabel metal3 s 69200 56040 70000 56160 0 FreeSans 480 0 0 0 out_7
port 506 nsew signal tristate
flabel metal3 s 69200 11160 70000 11280 0 FreeSans 480 0 0 0 rst
port 507 nsew signal tristate
flabel metal3 s 69200 3680 70000 3800 0 FreeSans 480 0 0 0 serial_data_rlbp_out
port 508 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 509 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 509 nsew power bidirectional
flabel metal4 s 65648 2128 65968 57712 0 FreeSans 1920 90 0 0 vccd1
port 509 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 510 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 510 nsew ground bidirectional
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wb_clk_i
port 511 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wb_rst_i
port 512 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 513 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 514 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 515 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 516 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 517 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 518 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 519 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 520 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 521 nsew signal input
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 522 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 523 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 524 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 525 nsew signal input
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 526 nsew signal input
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 527 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 528 nsew signal input
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 529 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 530 nsew signal input
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 531 nsew signal input
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 532 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 533 nsew signal input
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 534 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 535 nsew signal input
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 536 nsew signal input
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 537 nsew signal input
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 538 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 539 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 540 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 541 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 542 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 543 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 544 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 545 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 546 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 547 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 548 nsew signal input
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 549 nsew signal input
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 550 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 551 nsew signal input
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 552 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 553 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 554 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 555 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 556 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 557 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 558 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 559 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 560 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 561 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 562 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 563 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 564 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 565 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 566 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 567 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 568 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 569 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 570 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 571 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 572 nsew signal input
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 573 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 574 nsew signal input
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 575 nsew signal input
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 576 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 577 nsew signal input
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 578 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 579 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 580 nsew signal tristate
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 581 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 582 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 583 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 584 nsew signal tristate
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 585 nsew signal tristate
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 586 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 587 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 588 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 589 nsew signal tristate
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 590 nsew signal tristate
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 591 nsew signal tristate
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 592 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 593 nsew signal tristate
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 594 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 595 nsew signal tristate
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 596 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 597 nsew signal tristate
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 598 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 599 nsew signal tristate
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 600 nsew signal tristate
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 601 nsew signal tristate
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 602 nsew signal tristate
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 603 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 604 nsew signal tristate
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 605 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 606 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 607 nsew signal tristate
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 608 nsew signal tristate
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 609 nsew signal tristate
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 610 nsew signal tristate
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 611 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 612 nsew signal input
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 613 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 614 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 615 nsew signal input
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_we_i
port 616 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 70000 60000
<< end >>
