magic
tech sky130B
magscale 1 2
timestamp 1662590442
<< viali >>
rect 4353 7361 4387 7395
rect 4997 7361 5031 7395
rect 5825 7361 5859 7395
rect 7113 7361 7147 7395
rect 7573 7361 7607 7395
rect 8401 7361 8435 7395
rect 9137 7361 9171 7395
rect 9873 7361 9907 7395
rect 10517 7361 10551 7395
rect 11897 7361 11931 7395
rect 12633 7361 12667 7395
rect 13277 7361 13311 7395
rect 14657 7361 14691 7395
rect 15485 7361 15519 7395
rect 15945 7361 15979 7395
rect 17233 7361 17267 7395
rect 18061 7361 18095 7395
rect 18705 7361 18739 7395
rect 19533 7361 19567 7395
rect 20177 7361 20211 7395
rect 21281 7361 21315 7395
rect 22293 7361 22327 7395
rect 22937 7361 22971 7395
rect 23673 7361 23707 7395
rect 25145 7361 25179 7395
rect 25605 7361 25639 7395
rect 26433 7361 26467 7395
rect 27721 7361 27755 7395
rect 28365 7361 28399 7395
rect 29009 7361 29043 7395
rect 29837 7361 29871 7395
rect 30573 7361 30607 7395
rect 31217 7361 31251 7395
rect 32137 7361 32171 7395
rect 32781 7361 32815 7395
rect 33517 7361 33551 7395
rect 34713 7361 34747 7395
rect 35357 7361 35391 7395
rect 37289 7361 37323 7395
rect 37933 7361 37967 7395
rect 38577 7361 38611 7395
rect 39865 7361 39899 7395
rect 40509 7361 40543 7395
rect 41153 7361 41187 7395
rect 42441 7361 42475 7395
rect 43729 7361 43763 7395
rect 45017 7361 45051 7395
rect 45661 7361 45695 7395
rect 46305 7361 46339 7395
rect 47593 7361 47627 7395
rect 48237 7361 48271 7395
rect 48881 7361 48915 7395
rect 50169 7361 50203 7395
rect 50813 7361 50847 7395
rect 51457 7361 51491 7395
rect 52745 7361 52779 7395
rect 53389 7361 53423 7395
rect 54033 7361 54067 7395
rect 55321 7361 55355 7395
rect 55965 7361 55999 7395
rect 56609 7361 56643 7395
rect 36001 7293 36035 7327
rect 43085 7225 43119 7259
rect 6377 6817 6411 6851
rect 11437 6817 11471 6851
rect 14197 6817 14231 6851
rect 16957 6817 16991 6851
rect 21097 6817 21131 6851
rect 24409 6817 24443 6851
rect 27077 6817 27111 6851
rect 36277 6817 36311 6851
rect 39865 6817 39899 6851
rect 43637 6817 43671 6851
rect 46397 6817 46431 6851
rect 49157 6817 49191 6851
rect 54217 6817 54251 6851
rect 26525 6681 26559 6715
rect 27813 6681 27847 6715
rect 9965 6613 9999 6647
rect 33517 6613 33551 6647
rect 52193 6613 52227 6647
rect 8217 6205 8251 6239
rect 20729 6205 20763 6239
rect 11897 6137 11931 6171
rect 33885 6137 33919 6171
rect 50537 6137 50571 6171
rect 8769 6069 8803 6103
rect 9321 6069 9355 6103
rect 9781 6069 9815 6103
rect 10517 6069 10551 6103
rect 21189 6069 21223 6103
rect 23305 6069 23339 6103
rect 25697 6069 25731 6103
rect 26341 6069 26375 6103
rect 26985 6069 27019 6103
rect 27997 6069 28031 6103
rect 30481 6069 30515 6103
rect 31033 6069 31067 6103
rect 33241 6069 33275 6103
rect 34621 6069 34655 6103
rect 35081 6069 35115 6103
rect 35725 6069 35759 6103
rect 45569 6069 45603 6103
rect 49893 6069 49927 6103
rect 51181 6069 51215 6103
rect 51917 6069 51951 6103
rect 52745 6069 52779 6103
rect 4813 5865 4847 5899
rect 34713 5865 34747 5899
rect 40509 5865 40543 5899
rect 42625 5865 42659 5899
rect 53665 5865 53699 5899
rect 26433 5797 26467 5831
rect 30941 5797 30975 5831
rect 31033 5797 31067 5831
rect 48145 5797 48179 5831
rect 7205 5729 7239 5763
rect 28181 5729 28215 5763
rect 31677 5729 31711 5763
rect 34897 5729 34931 5763
rect 35265 5729 35299 5763
rect 37565 5729 37599 5763
rect 37657 5729 37691 5763
rect 45937 5729 45971 5763
rect 53021 5729 53055 5763
rect 7757 5661 7791 5695
rect 8401 5661 8435 5695
rect 9413 5661 9447 5695
rect 10149 5661 10183 5695
rect 10977 5661 11011 5695
rect 12081 5661 12115 5695
rect 12909 5661 12943 5695
rect 14841 5661 14875 5695
rect 15853 5661 15887 5695
rect 16497 5661 16531 5695
rect 17049 5661 17083 5695
rect 26893 5661 26927 5695
rect 27721 5661 27755 5695
rect 30941 5661 30975 5695
rect 31769 5661 31803 5695
rect 31953 5661 31987 5695
rect 33425 5661 33459 5695
rect 33517 5661 33551 5695
rect 35725 5661 35759 5695
rect 36277 5661 36311 5695
rect 36461 5661 36495 5695
rect 37289 5661 37323 5695
rect 38209 5661 38243 5695
rect 43085 5661 43119 5695
rect 45293 5661 45327 5695
rect 45477 5661 45511 5695
rect 50353 5661 50387 5695
rect 50997 5661 51031 5695
rect 51733 5661 51767 5695
rect 52377 5661 52411 5695
rect 5917 5593 5951 5627
rect 6469 5593 6503 5627
rect 31217 5593 31251 5627
rect 32137 5593 32171 5627
rect 32689 5593 32723 5627
rect 33701 5593 33735 5627
rect 36369 5593 36403 5627
rect 39957 5593 39991 5627
rect 47593 5593 47627 5627
rect 55873 5593 55907 5627
rect 8217 5525 8251 5559
rect 9597 5525 9631 5559
rect 14381 5525 14415 5559
rect 16313 5525 16347 5559
rect 20085 5525 20119 5559
rect 20729 5525 20763 5559
rect 21557 5525 21591 5559
rect 22385 5525 22419 5559
rect 22937 5525 22971 5559
rect 23489 5525 23523 5559
rect 24685 5525 24719 5559
rect 25145 5525 25179 5559
rect 25789 5525 25823 5559
rect 27537 5525 27571 5559
rect 28825 5525 28859 5559
rect 29745 5525 29779 5559
rect 30389 5525 30423 5559
rect 33425 5525 33459 5559
rect 35081 5525 35115 5559
rect 41705 5525 41739 5559
rect 45385 5525 45419 5559
rect 46489 5525 46523 5559
rect 47041 5525 47075 5559
rect 49617 5525 49651 5559
rect 55321 5525 55355 5559
rect 4353 5321 4387 5355
rect 7573 5321 7607 5355
rect 20729 5321 20763 5355
rect 23857 5321 23891 5355
rect 28365 5321 28399 5355
rect 31309 5321 31343 5355
rect 35173 5321 35207 5355
rect 39313 5321 39347 5355
rect 41705 5321 41739 5355
rect 42625 5321 42659 5355
rect 44649 5321 44683 5355
rect 50905 5321 50939 5355
rect 13461 5253 13495 5287
rect 19073 5253 19107 5287
rect 21189 5253 21223 5287
rect 22753 5253 22787 5287
rect 24501 5253 24535 5287
rect 33149 5253 33183 5287
rect 45293 5253 45327 5287
rect 48329 5253 48363 5287
rect 48545 5253 48579 5287
rect 4261 5185 4295 5219
rect 4353 5185 4387 5219
rect 5181 5185 5215 5219
rect 5273 5185 5307 5219
rect 5365 5185 5399 5219
rect 5549 5185 5583 5219
rect 6469 5185 6503 5219
rect 6929 5185 6963 5219
rect 7757 5185 7791 5219
rect 8401 5185 8435 5219
rect 8861 5185 8895 5219
rect 9505 5185 9539 5219
rect 16129 5185 16163 5219
rect 18245 5185 18279 5219
rect 18797 5185 18831 5219
rect 25145 5185 25179 5219
rect 25789 5185 25823 5219
rect 26985 5185 27019 5219
rect 27241 5185 27275 5219
rect 30481 5185 30515 5219
rect 32137 5185 32171 5219
rect 32321 5185 32355 5219
rect 32965 5185 32999 5219
rect 34161 5185 34195 5219
rect 34989 5185 35023 5219
rect 35265 5185 35299 5219
rect 36001 5185 36035 5219
rect 36737 5185 36771 5219
rect 37657 5185 37691 5219
rect 39305 5185 39339 5219
rect 39497 5185 39531 5219
rect 39957 5185 39991 5219
rect 40178 5185 40212 5219
rect 40509 5185 40543 5219
rect 41061 5185 41095 5219
rect 41245 5185 41279 5219
rect 43453 5185 43487 5219
rect 43637 5185 43671 5219
rect 44557 5185 44591 5219
rect 44741 5185 44775 5219
rect 45201 5185 45235 5219
rect 45477 5185 45511 5219
rect 49157 5185 49191 5219
rect 50721 5185 50755 5219
rect 50905 5185 50939 5219
rect 51365 5185 51399 5219
rect 52009 5185 52043 5219
rect 52745 5185 52779 5219
rect 53573 5185 53607 5219
rect 55137 5185 55171 5219
rect 4077 5117 4111 5151
rect 12633 5117 12667 5151
rect 22293 5117 22327 5151
rect 30757 5117 30791 5151
rect 32229 5117 32263 5151
rect 33977 5117 34011 5151
rect 35817 5117 35851 5151
rect 36185 5117 36219 5151
rect 42441 5117 42475 5151
rect 42809 5117 42843 5151
rect 46581 5117 46615 5151
rect 47041 5117 47075 5151
rect 49801 5117 49835 5151
rect 8217 5049 8251 5083
rect 9045 5049 9079 5083
rect 11897 5049 11931 5083
rect 15485 5049 15519 5083
rect 18061 5049 18095 5083
rect 18889 5049 18923 5083
rect 32781 5049 32815 5083
rect 40233 5049 40267 5083
rect 46857 5049 46891 5083
rect 48697 5049 48731 5083
rect 51549 5049 51583 5083
rect 54033 5049 54067 5083
rect 3249 4981 3283 5015
rect 4905 4981 4939 5015
rect 7113 4981 7147 5015
rect 9689 4981 9723 5015
rect 10333 4981 10367 5015
rect 10977 4981 11011 5015
rect 14197 4981 14231 5015
rect 14841 4981 14875 5015
rect 15945 4981 15979 5015
rect 16773 4981 16807 5015
rect 17233 4981 17267 5015
rect 18981 4981 19015 5015
rect 19993 4981 20027 5015
rect 23397 4981 23431 5015
rect 24961 4981 24995 5015
rect 26433 4981 26467 5015
rect 28825 4981 28859 5015
rect 34345 4981 34379 5015
rect 34805 4981 34839 5015
rect 37565 4981 37599 5015
rect 38209 4981 38243 5015
rect 41245 4981 41279 5015
rect 42809 4981 42843 5015
rect 43453 4981 43487 5015
rect 45661 4981 45695 5015
rect 47593 4981 47627 5015
rect 48513 4981 48547 5015
rect 49341 4981 49375 5015
rect 52101 4981 52135 5015
rect 52837 4981 52871 5015
rect 53389 4981 53423 5015
rect 55321 4981 55355 5015
rect 55781 4981 55815 5015
rect 56333 4981 56367 5015
rect 3249 4777 3283 4811
rect 6561 4777 6595 4811
rect 12725 4777 12759 4811
rect 18153 4777 18187 4811
rect 23857 4777 23891 4811
rect 30113 4777 30147 4811
rect 33149 4777 33183 4811
rect 36921 4777 36955 4811
rect 41061 4777 41095 4811
rect 42551 4777 42585 4811
rect 51181 4777 51215 4811
rect 55689 4777 55723 4811
rect 3157 4709 3191 4743
rect 9321 4709 9355 4743
rect 11805 4709 11839 4743
rect 18613 4709 18647 4743
rect 20637 4709 20671 4743
rect 25053 4709 25087 4743
rect 27629 4709 27663 4743
rect 32597 4709 32631 4743
rect 37841 4709 37875 4743
rect 44281 4709 44315 4743
rect 48605 4709 48639 4743
rect 6469 4641 6503 4675
rect 8401 4641 8435 4675
rect 10425 4641 10459 4675
rect 12633 4641 12667 4675
rect 15301 4641 15335 4675
rect 16957 4641 16991 4675
rect 18337 4641 18371 4675
rect 19257 4641 19291 4675
rect 25881 4641 25915 4675
rect 26157 4641 26191 4675
rect 29561 4641 29595 4675
rect 35173 4641 35207 4675
rect 35449 4641 35483 4675
rect 42809 4641 42843 4675
rect 46029 4641 46063 4675
rect 46305 4641 46339 4675
rect 53113 4641 53147 4675
rect 53757 4641 53791 4675
rect 3249 4573 3283 4607
rect 3801 4573 3835 4607
rect 4445 4573 4479 4607
rect 4712 4573 4746 4607
rect 6561 4573 6595 4607
rect 7573 4573 7607 4607
rect 7757 4573 7791 4607
rect 9965 4573 9999 4607
rect 12449 4573 12483 4607
rect 12725 4573 12759 4607
rect 13553 4573 13587 4607
rect 14473 4573 14507 4607
rect 15761 4573 15795 4607
rect 17601 4573 17635 4607
rect 17693 4573 17727 4607
rect 18429 4573 18463 4607
rect 21373 4573 21407 4607
rect 22385 4573 22419 4607
rect 22477 4573 22511 4607
rect 22569 4573 22603 4607
rect 22753 4573 22787 4607
rect 23213 4573 23247 4607
rect 23397 4573 23431 4607
rect 23489 4573 23523 4607
rect 23581 4573 23615 4607
rect 24409 4573 24443 4607
rect 24593 4573 24627 4607
rect 24685 4573 24719 4607
rect 24777 4573 24811 4607
rect 28273 4573 28307 4607
rect 28825 4573 28859 4607
rect 29929 4573 29963 4607
rect 30757 4573 30791 4607
rect 33885 4573 33919 4607
rect 34161 4573 34195 4607
rect 37657 4573 37691 4607
rect 38393 4573 38427 4607
rect 40049 4573 40083 4607
rect 43453 4573 43487 4607
rect 44281 4573 44315 4607
rect 44465 4573 44499 4607
rect 45201 4573 45235 4607
rect 49341 4573 49375 4607
rect 49617 4573 49651 4607
rect 50169 4573 50203 4607
rect 51273 4573 51307 4607
rect 52837 4573 52871 4607
rect 54033 4573 54067 4607
rect 55505 4573 55539 4607
rect 56149 4573 56183 4607
rect 2973 4505 3007 4539
rect 6285 4505 6319 4539
rect 10692 4505 10726 4539
rect 17417 4505 17451 4539
rect 18153 4505 18187 4539
rect 19524 4505 19558 4539
rect 22109 4505 22143 4539
rect 28181 4505 28215 4539
rect 31002 4505 31036 4539
rect 39957 4505 39991 4539
rect 45109 4505 45143 4539
rect 55321 4505 55355 4539
rect 3985 4437 4019 4471
rect 5825 4437 5859 4471
rect 7113 4437 7147 4471
rect 7665 4437 7699 4471
rect 9781 4437 9815 4471
rect 12265 4437 12299 4471
rect 14657 4437 14691 4471
rect 15945 4437 15979 4471
rect 17693 4437 17727 4471
rect 29745 4437 29779 4471
rect 32137 4437 32171 4471
rect 38945 4437 38979 4471
rect 40601 4437 40635 4471
rect 47777 4437 47811 4471
rect 50353 4437 50387 4471
rect 52101 4437 52135 4471
rect 54769 4437 54803 4471
rect 56701 4437 56735 4471
rect 57253 4437 57287 4471
rect 3709 4233 3743 4267
rect 10609 4233 10643 4267
rect 51089 4233 51123 4267
rect 55045 4233 55079 4267
rect 2697 4165 2731 4199
rect 13369 4165 13403 4199
rect 16037 4165 16071 4199
rect 17877 4165 17911 4199
rect 28549 4165 28583 4199
rect 35909 4165 35943 4199
rect 49065 4165 49099 4199
rect 53021 4165 53055 4199
rect 2881 4097 2915 4131
rect 3433 4097 3467 4131
rect 3525 4097 3559 4131
rect 4169 4097 4203 4131
rect 4425 4097 4459 4131
rect 6561 4097 6595 4131
rect 7389 4097 7423 4131
rect 9606 4097 9640 4131
rect 9873 4097 9907 4131
rect 10793 4097 10827 4131
rect 11805 4097 11839 4131
rect 11897 4097 11931 4131
rect 11989 4097 12023 4131
rect 12173 4097 12207 4131
rect 13093 4097 13127 4131
rect 13185 4097 13219 4131
rect 14657 4097 14691 4131
rect 15117 4097 15151 4131
rect 15761 4097 15795 4131
rect 15853 4097 15887 4131
rect 18153 4097 18187 4131
rect 18797 4097 18831 4131
rect 21833 4097 21867 4131
rect 22017 4097 22051 4131
rect 22109 4097 22143 4131
rect 22201 4097 22235 4131
rect 23581 4097 23615 4131
rect 24133 4097 24167 4131
rect 24389 4097 24423 4131
rect 26249 4097 26283 4131
rect 30757 4097 30791 4131
rect 32597 4097 32631 4131
rect 33425 4097 33459 4131
rect 38209 4097 38243 4131
rect 39129 4097 39163 4131
rect 39221 4097 39255 4131
rect 41705 4097 41739 4131
rect 42901 4097 42935 4131
rect 43821 4097 43855 4131
rect 43913 4097 43947 4131
rect 45753 4097 45787 4131
rect 46581 4097 46615 4131
rect 49341 4097 49375 4131
rect 49801 4097 49835 4131
rect 51273 4097 51307 4131
rect 52745 4097 52779 4131
rect 55873 4097 55907 4131
rect 56701 4097 56735 4131
rect 10977 4029 11011 4063
rect 11529 4029 11563 4063
rect 14013 4029 14047 4063
rect 17969 4029 18003 4063
rect 19073 4029 19107 4063
rect 22477 4029 22511 4063
rect 33701 4029 33735 4063
rect 37289 4029 37323 4063
rect 41429 4029 41463 4063
rect 55597 4029 55631 4063
rect 6745 3961 6779 3995
rect 8033 3961 8067 3995
rect 12909 3961 12943 3995
rect 17417 3961 17451 3995
rect 25513 3961 25547 3995
rect 28089 3961 28123 3995
rect 30941 3961 30975 3995
rect 32781 3961 32815 3995
rect 36553 3961 36587 3995
rect 37565 3961 37599 3995
rect 45109 3961 45143 3995
rect 49893 3961 49927 3995
rect 51733 3961 51767 3995
rect 2145 3893 2179 3927
rect 5549 3893 5583 3927
rect 8493 3893 8527 3927
rect 13093 3893 13127 3927
rect 15301 3893 15335 3927
rect 15945 3893 15979 3927
rect 18153 3893 18187 3927
rect 18337 3893 18371 3927
rect 20545 3893 20579 3927
rect 21281 3893 21315 3927
rect 23397 3893 23431 3927
rect 26433 3893 26467 3927
rect 27169 3893 27203 3927
rect 29837 3893 29871 3927
rect 31401 3893 31435 3927
rect 35173 3893 35207 3927
rect 36001 3893 36035 3927
rect 37749 3893 37783 3927
rect 39957 3893 39991 3927
rect 43085 3893 43119 3927
rect 44465 3893 44499 3927
rect 45937 3893 45971 3927
rect 46673 3893 46707 3927
rect 47593 3893 47627 3927
rect 50445 3893 50479 3927
rect 54493 3893 54527 3927
rect 57253 3893 57287 3927
rect 57897 3893 57931 3927
rect 3801 3689 3835 3723
rect 6377 3689 6411 3723
rect 11805 3689 11839 3723
rect 14473 3689 14507 3723
rect 15945 3689 15979 3723
rect 18245 3689 18279 3723
rect 18705 3689 18739 3723
rect 25329 3689 25363 3723
rect 30941 3689 30975 3723
rect 35449 3689 35483 3723
rect 40049 3689 40083 3723
rect 41153 3689 41187 3723
rect 43913 3689 43947 3723
rect 45753 3689 45787 3723
rect 46949 3689 46983 3723
rect 51641 3689 51675 3723
rect 9137 3621 9171 3655
rect 15485 3621 15519 3655
rect 16405 3621 16439 3655
rect 17785 3621 17819 3655
rect 20361 3621 20395 3655
rect 43453 3621 43487 3655
rect 50169 3621 50203 3655
rect 55321 3621 55355 3655
rect 57805 3621 57839 3655
rect 1501 3553 1535 3587
rect 4261 3553 4295 3587
rect 4445 3553 4479 3587
rect 6285 3553 6319 3587
rect 9873 3553 9907 3587
rect 12357 3553 12391 3587
rect 14263 3553 14297 3587
rect 16037 3553 16071 3587
rect 17141 3553 17175 3587
rect 18337 3553 18371 3587
rect 19717 3553 19751 3587
rect 21189 3553 21223 3587
rect 24777 3553 24811 3587
rect 27261 3553 27295 3587
rect 27537 3553 27571 3587
rect 30389 3553 30423 3587
rect 36001 3553 36035 3587
rect 37749 3553 37783 3587
rect 38669 3553 38703 3587
rect 45201 3553 45235 3587
rect 49065 3553 49099 3587
rect 49341 3553 49375 3587
rect 52285 3553 52319 3587
rect 52561 3553 52595 3587
rect 55873 3553 55907 3587
rect 3065 3485 3099 3519
rect 5273 3485 5307 3519
rect 6377 3485 6411 3519
rect 7757 3485 7791 3519
rect 8401 3485 8435 3519
rect 10609 3485 10643 3519
rect 10701 3485 10735 3519
rect 11345 3485 11379 3519
rect 14105 3485 14139 3519
rect 14473 3485 14507 3519
rect 14657 3485 14691 3519
rect 16221 3485 16255 3519
rect 18521 3485 18555 3519
rect 21005 3485 21039 3519
rect 21649 3485 21683 3519
rect 23121 3485 23155 3519
rect 23857 3485 23891 3519
rect 24961 3485 24995 3519
rect 26065 3485 26099 3519
rect 26801 3485 26835 3519
rect 29561 3485 29595 3519
rect 30573 3485 30607 3519
rect 31401 3485 31435 3519
rect 32321 3485 32355 3519
rect 32781 3485 32815 3519
rect 33425 3485 33459 3519
rect 34713 3485 34747 3519
rect 37105 3485 37139 3519
rect 38945 3485 38979 3519
rect 39865 3485 39899 3519
rect 40509 3485 40543 3519
rect 42533 3485 42567 3519
rect 42809 3485 42843 3519
rect 43269 3485 43303 3519
rect 46581 3485 46615 3519
rect 50905 3485 50939 3519
rect 51181 3485 51215 3519
rect 54585 3485 54619 3519
rect 56517 3485 56551 3519
rect 57345 3485 57379 3519
rect 57989 3485 58023 3519
rect 2605 3417 2639 3451
rect 5917 3417 5951 3451
rect 9689 3417 9723 3451
rect 10425 3417 10459 3451
rect 13185 3417 13219 3451
rect 15945 3417 15979 3451
rect 18245 3417 18279 3451
rect 20821 3417 20855 3451
rect 24869 3417 24903 3451
rect 32229 3417 32263 3451
rect 38853 3417 38887 3451
rect 45293 3417 45327 3451
rect 2053 3349 2087 3383
rect 3157 3349 3191 3383
rect 4169 3349 4203 3383
rect 5457 3349 5491 3383
rect 6561 3349 6595 3383
rect 7113 3349 7147 3383
rect 10701 3349 10735 3383
rect 12173 3349 12207 3383
rect 12265 3349 12299 3383
rect 13093 3349 13127 3383
rect 19901 3349 19935 3383
rect 19993 3349 20027 3383
rect 21833 3349 21867 3383
rect 22937 3349 22971 3383
rect 23673 3349 23707 3383
rect 25881 3349 25915 3383
rect 26617 3349 26651 3383
rect 29009 3349 29043 3383
rect 30481 3349 30515 3383
rect 31585 3349 31619 3383
rect 34069 3349 34103 3383
rect 36185 3349 36219 3383
rect 36277 3349 36311 3383
rect 36645 3349 36679 3383
rect 39313 3349 39347 3383
rect 41797 3349 41831 3383
rect 45385 3349 45419 3383
rect 46949 3349 46983 3383
rect 47133 3349 47167 3383
rect 47593 3349 47627 3383
rect 54033 3349 54067 3383
rect 55689 3349 55723 3383
rect 55781 3349 55815 3383
rect 57161 3349 57195 3383
rect 2973 3145 3007 3179
rect 6837 3145 6871 3179
rect 11621 3145 11655 3179
rect 13461 3145 13495 3179
rect 14749 3145 14783 3179
rect 17693 3145 17727 3179
rect 20821 3145 20855 3179
rect 23857 3145 23891 3179
rect 31217 3145 31251 3179
rect 31585 3145 31619 3179
rect 50282 3145 50316 3179
rect 50445 3145 50479 3179
rect 19686 3077 19720 3111
rect 25145 3077 25179 3111
rect 28641 3077 28675 3111
rect 30389 3077 30423 3111
rect 33885 3077 33919 3111
rect 39957 3077 39991 3111
rect 41797 3077 41831 3111
rect 47041 3077 47075 3111
rect 49525 3077 49559 3111
rect 50077 3077 50111 3111
rect 56057 3077 56091 3111
rect 56149 3077 56183 3111
rect 1869 3009 1903 3043
rect 3433 3009 3467 3043
rect 4353 3009 4387 3043
rect 4629 3009 4663 3043
rect 5273 3009 5307 3043
rect 5641 3009 5675 3043
rect 6469 3009 6503 3043
rect 6653 3009 6687 3043
rect 7021 3009 7055 3043
rect 7849 3009 7883 3043
rect 8769 3009 8803 3043
rect 9689 3009 9723 3043
rect 12265 3009 12299 3043
rect 12817 3009 12851 3043
rect 12909 3009 12943 3043
rect 13277 3009 13311 3043
rect 14381 3009 14415 3043
rect 15577 3009 15611 3043
rect 15945 3009 15979 3043
rect 16037 3009 16071 3043
rect 17509 3009 17543 3043
rect 19441 3009 19475 3043
rect 22201 3009 22235 3043
rect 22937 3009 22971 3043
rect 26065 3009 26099 3043
rect 27261 3009 27295 3043
rect 31125 3009 31159 3043
rect 33609 3009 33643 3043
rect 37289 3009 37323 3043
rect 37933 3009 37967 3043
rect 40049 3009 40083 3043
rect 43729 3009 43763 3043
rect 45661 3009 45695 3043
rect 46305 3009 46339 3043
rect 50905 3009 50939 3043
rect 54953 3009 54987 3043
rect 57897 3009 57931 3043
rect 4537 2941 4571 2975
rect 5181 2941 5215 2975
rect 14473 2941 14507 2975
rect 30941 2941 30975 2975
rect 40509 2941 40543 2975
rect 44373 2941 44407 2975
rect 48881 2941 48915 2975
rect 53389 2941 53423 2975
rect 55229 2941 55263 2975
rect 56241 2941 56275 2975
rect 3617 2873 3651 2907
rect 10977 2873 11011 2907
rect 15393 2873 15427 2907
rect 18337 2873 18371 2907
rect 22017 2873 22051 2907
rect 32781 2873 32815 2907
rect 35817 2873 35851 2907
rect 36461 2873 36495 2907
rect 38577 2873 38611 2907
rect 43085 2873 43119 2907
rect 48237 2873 48271 2907
rect 51549 2873 51583 2907
rect 56885 2873 56919 2907
rect 2421 2805 2455 2839
rect 4169 2805 4203 2839
rect 4353 2805 4387 2839
rect 5641 2805 5675 2839
rect 5825 2805 5859 2839
rect 6561 2805 6595 2839
rect 7665 2805 7699 2839
rect 8585 2805 8619 2839
rect 10333 2805 10367 2839
rect 13277 2805 13311 2839
rect 14381 2805 14415 2839
rect 15577 2805 15611 2839
rect 17049 2805 17083 2839
rect 18981 2805 19015 2839
rect 22753 2805 22787 2839
rect 26249 2805 26283 2839
rect 27077 2805 27111 2839
rect 28181 2805 28215 2839
rect 32137 2805 32171 2839
rect 35357 2805 35391 2839
rect 39221 2805 39255 2839
rect 41153 2805 41187 2839
rect 42441 2805 42475 2839
rect 45017 2805 45051 2839
rect 47593 2805 47627 2839
rect 50261 2805 50295 2839
rect 52745 2805 52779 2839
rect 54217 2805 54251 2839
rect 55689 2805 55723 2839
rect 4077 2601 4111 2635
rect 11529 2601 11563 2635
rect 13185 2601 13219 2635
rect 14197 2601 14231 2635
rect 17417 2601 17451 2635
rect 22201 2601 22235 2635
rect 25789 2601 25823 2635
rect 34069 2601 34103 2635
rect 34713 2601 34747 2635
rect 35357 2601 35391 2635
rect 37933 2601 37967 2635
rect 39221 2601 39255 2635
rect 43729 2601 43763 2635
rect 47593 2601 47627 2635
rect 49525 2601 49559 2635
rect 53389 2601 53423 2635
rect 55597 2601 55631 2635
rect 55781 2601 55815 2635
rect 2605 2533 2639 2567
rect 5825 2533 5859 2567
rect 10977 2533 11011 2567
rect 15485 2533 15519 2567
rect 20637 2533 20671 2567
rect 23765 2533 23799 2567
rect 26157 2533 26191 2567
rect 29009 2533 29043 2567
rect 33425 2533 33459 2567
rect 37289 2533 37323 2567
rect 41153 2533 41187 2567
rect 45017 2533 45051 2567
rect 45661 2533 45695 2567
rect 50169 2533 50203 2567
rect 54677 2533 54711 2567
rect 57897 2533 57931 2567
rect 5181 2465 5215 2499
rect 5549 2465 5583 2499
rect 5666 2465 5700 2499
rect 6653 2465 6687 2499
rect 18061 2465 18095 2499
rect 18705 2465 18739 2499
rect 19993 2465 20027 2499
rect 21281 2465 21315 2499
rect 24501 2465 24535 2499
rect 24685 2465 24719 2499
rect 26985 2465 27019 2499
rect 30297 2465 30331 2499
rect 32137 2465 32171 2499
rect 40509 2465 40543 2499
rect 44465 2465 44499 2499
rect 48237 2465 48271 2499
rect 54033 2465 54067 2499
rect 2421 2397 2455 2431
rect 3065 2397 3099 2431
rect 3893 2397 3927 2431
rect 4721 2397 4755 2431
rect 6561 2397 6595 2431
rect 6745 2397 6779 2431
rect 7481 2397 7515 2431
rect 9229 2397 9263 2431
rect 9689 2397 9723 2431
rect 10793 2397 10827 2431
rect 12265 2397 12299 2431
rect 12725 2397 12759 2431
rect 13093 2397 13127 2431
rect 13369 2397 13403 2431
rect 14841 2397 14875 2431
rect 16129 2397 16163 2431
rect 22385 2397 22419 2431
rect 23121 2397 23155 2431
rect 23581 2397 23615 2431
rect 27241 2397 27275 2431
rect 29837 2397 29871 2431
rect 31033 2397 31067 2431
rect 32781 2397 32815 2431
rect 36001 2397 36035 2431
rect 36737 2397 36771 2431
rect 38577 2397 38611 2431
rect 39865 2397 39899 2431
rect 42441 2397 42475 2431
rect 43085 2397 43119 2431
rect 46305 2397 46339 2431
rect 48881 2397 48915 2431
rect 50813 2397 50847 2431
rect 51457 2397 51491 2431
rect 52745 2397 52779 2431
rect 55321 2397 55355 2431
rect 56241 2397 56275 2431
rect 56885 2397 56919 2431
rect 1961 2329 1995 2363
rect 3249 2261 3283 2295
rect 5457 2261 5491 2295
rect 7711 2261 7745 2295
rect 9045 2261 9079 2295
rect 9873 2261 9907 2295
rect 12909 2261 12943 2295
rect 19349 2261 19383 2295
rect 22937 2261 22971 2295
rect 24777 2261 24811 2295
rect 25145 2261 25179 2295
rect 25605 2261 25639 2295
rect 25789 2261 25823 2295
rect 28365 2261 28399 2295
rect 29653 2261 29687 2295
rect 41797 2261 41831 2295
rect 47041 2261 47075 2295
rect 52101 2261 52135 2295
<< metal1 >>
rect 1104 7642 58880 7664
rect 1104 7590 15398 7642
rect 15450 7590 15462 7642
rect 15514 7590 15526 7642
rect 15578 7590 15590 7642
rect 15642 7590 15654 7642
rect 15706 7590 29846 7642
rect 29898 7590 29910 7642
rect 29962 7590 29974 7642
rect 30026 7590 30038 7642
rect 30090 7590 30102 7642
rect 30154 7590 44294 7642
rect 44346 7590 44358 7642
rect 44410 7590 44422 7642
rect 44474 7590 44486 7642
rect 44538 7590 44550 7642
rect 44602 7590 58880 7642
rect 1104 7568 58880 7590
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4430 7392 4436 7404
rect 4387 7364 4436 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 4430 7352 4436 7364
rect 4488 7352 4494 7404
rect 4982 7392 4988 7404
rect 4943 7364 4988 7392
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 5810 7392 5816 7404
rect 5771 7364 5816 7392
rect 5810 7352 5816 7364
rect 5868 7352 5874 7404
rect 7098 7392 7104 7404
rect 7059 7364 7104 7392
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 7558 7392 7564 7404
rect 7519 7364 7564 7392
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 8386 7392 8392 7404
rect 8347 7364 8392 7392
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 9122 7392 9128 7404
rect 9083 7364 9128 7392
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 9861 7395 9919 7401
rect 9861 7361 9873 7395
rect 9907 7392 9919 7395
rect 9950 7392 9956 7404
rect 9907 7364 9956 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 10410 7352 10416 7404
rect 10468 7392 10474 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 10468 7364 10517 7392
rect 10468 7352 10474 7364
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 11882 7392 11888 7404
rect 11843 7364 11888 7392
rect 10505 7355 10563 7361
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 12618 7392 12624 7404
rect 12579 7364 12624 7392
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 13262 7392 13268 7404
rect 13223 7364 13268 7392
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 14642 7392 14648 7404
rect 14603 7364 14648 7392
rect 14642 7352 14648 7364
rect 14700 7352 14706 7404
rect 15286 7352 15292 7404
rect 15344 7392 15350 7404
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15344 7364 15485 7392
rect 15344 7352 15350 7364
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15930 7392 15936 7404
rect 15891 7364 15936 7392
rect 15473 7355 15531 7361
rect 15930 7352 15936 7364
rect 15988 7352 15994 7404
rect 17218 7392 17224 7404
rect 17179 7364 17224 7392
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 18046 7392 18052 7404
rect 18007 7364 18052 7392
rect 18046 7352 18052 7364
rect 18104 7352 18110 7404
rect 18690 7392 18696 7404
rect 18651 7364 18696 7392
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 19518 7392 19524 7404
rect 19479 7364 19524 7392
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 20162 7392 20168 7404
rect 20123 7364 20168 7392
rect 20162 7352 20168 7364
rect 20220 7352 20226 7404
rect 21266 7392 21272 7404
rect 21227 7364 21272 7392
rect 21266 7352 21272 7364
rect 21324 7352 21330 7404
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 22370 7392 22376 7404
rect 22327 7364 22376 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 22370 7352 22376 7364
rect 22428 7352 22434 7404
rect 22922 7392 22928 7404
rect 22883 7364 22928 7392
rect 22922 7352 22928 7364
rect 22980 7352 22986 7404
rect 23658 7392 23664 7404
rect 23619 7364 23664 7392
rect 23658 7352 23664 7364
rect 23716 7352 23722 7404
rect 25130 7392 25136 7404
rect 25091 7364 25136 7392
rect 25130 7352 25136 7364
rect 25188 7352 25194 7404
rect 25590 7392 25596 7404
rect 25551 7364 25596 7392
rect 25590 7352 25596 7364
rect 25648 7352 25654 7404
rect 26418 7392 26424 7404
rect 26379 7364 26424 7392
rect 26418 7352 26424 7364
rect 26476 7352 26482 7404
rect 27706 7392 27712 7404
rect 27667 7364 27712 7392
rect 27706 7352 27712 7364
rect 27764 7352 27770 7404
rect 28350 7392 28356 7404
rect 28311 7364 28356 7392
rect 28350 7352 28356 7364
rect 28408 7352 28414 7404
rect 28994 7392 29000 7404
rect 28955 7364 29000 7392
rect 28994 7352 29000 7364
rect 29052 7352 29058 7404
rect 29730 7352 29736 7404
rect 29788 7392 29794 7404
rect 29825 7395 29883 7401
rect 29825 7392 29837 7395
rect 29788 7364 29837 7392
rect 29788 7352 29794 7364
rect 29825 7361 29837 7364
rect 29871 7361 29883 7395
rect 30558 7392 30564 7404
rect 30519 7364 30564 7392
rect 29825 7355 29883 7361
rect 30558 7352 30564 7364
rect 30616 7352 30622 7404
rect 31202 7392 31208 7404
rect 31163 7364 31208 7392
rect 31202 7352 31208 7364
rect 31260 7352 31266 7404
rect 32122 7392 32128 7404
rect 32083 7364 32128 7392
rect 32122 7352 32128 7364
rect 32180 7352 32186 7404
rect 32766 7392 32772 7404
rect 32727 7364 32772 7392
rect 32766 7352 32772 7364
rect 32824 7352 32830 7404
rect 33410 7352 33416 7404
rect 33468 7392 33474 7404
rect 33505 7395 33563 7401
rect 33505 7392 33517 7395
rect 33468 7364 33517 7392
rect 33468 7352 33474 7364
rect 33505 7361 33517 7364
rect 33551 7361 33563 7395
rect 33505 7355 33563 7361
rect 33870 7352 33876 7404
rect 33928 7392 33934 7404
rect 34701 7395 34759 7401
rect 34701 7392 34713 7395
rect 33928 7364 34713 7392
rect 33928 7352 33934 7364
rect 34701 7361 34713 7364
rect 34747 7361 34759 7395
rect 34701 7355 34759 7361
rect 34790 7352 34796 7404
rect 34848 7392 34854 7404
rect 35345 7395 35403 7401
rect 35345 7392 35357 7395
rect 34848 7364 35357 7392
rect 34848 7352 34854 7364
rect 35345 7361 35357 7364
rect 35391 7361 35403 7395
rect 35345 7355 35403 7361
rect 36630 7352 36636 7404
rect 36688 7392 36694 7404
rect 37277 7395 37335 7401
rect 37277 7392 37289 7395
rect 36688 7364 37289 7392
rect 36688 7352 36694 7364
rect 37277 7361 37289 7364
rect 37323 7361 37335 7395
rect 37277 7355 37335 7361
rect 37550 7352 37556 7404
rect 37608 7392 37614 7404
rect 37921 7395 37979 7401
rect 37921 7392 37933 7395
rect 37608 7364 37933 7392
rect 37608 7352 37614 7364
rect 37921 7361 37933 7364
rect 37967 7361 37979 7395
rect 37921 7355 37979 7361
rect 38010 7352 38016 7404
rect 38068 7392 38074 7404
rect 38565 7395 38623 7401
rect 38565 7392 38577 7395
rect 38068 7364 38577 7392
rect 38068 7352 38074 7364
rect 38565 7361 38577 7364
rect 38611 7361 38623 7395
rect 38565 7355 38623 7361
rect 38930 7352 38936 7404
rect 38988 7392 38994 7404
rect 39853 7395 39911 7401
rect 39853 7392 39865 7395
rect 38988 7364 39865 7392
rect 38988 7352 38994 7364
rect 39853 7361 39865 7364
rect 39899 7361 39911 7395
rect 40494 7392 40500 7404
rect 40455 7364 40500 7392
rect 39853 7355 39911 7361
rect 40494 7352 40500 7364
rect 40552 7352 40558 7404
rect 41138 7392 41144 7404
rect 41099 7364 41144 7392
rect 41138 7352 41144 7364
rect 41196 7352 41202 7404
rect 41690 7352 41696 7404
rect 41748 7392 41754 7404
rect 42429 7395 42487 7401
rect 42429 7392 42441 7395
rect 41748 7364 42441 7392
rect 41748 7352 41754 7364
rect 42429 7361 42441 7364
rect 42475 7361 42487 7395
rect 42429 7355 42487 7361
rect 43070 7352 43076 7404
rect 43128 7392 43134 7404
rect 43717 7395 43775 7401
rect 43717 7392 43729 7395
rect 43128 7364 43729 7392
rect 43128 7352 43134 7364
rect 43717 7361 43729 7364
rect 43763 7361 43775 7395
rect 43717 7355 43775 7361
rect 44634 7352 44640 7404
rect 44692 7392 44698 7404
rect 45005 7395 45063 7401
rect 45005 7392 45017 7395
rect 44692 7364 45017 7392
rect 44692 7352 44698 7364
rect 45005 7361 45017 7364
rect 45051 7361 45063 7395
rect 45005 7355 45063 7361
rect 45186 7352 45192 7404
rect 45244 7392 45250 7404
rect 45649 7395 45707 7401
rect 45649 7392 45661 7395
rect 45244 7364 45661 7392
rect 45244 7352 45250 7364
rect 45649 7361 45661 7364
rect 45695 7361 45707 7395
rect 45649 7355 45707 7361
rect 45830 7352 45836 7404
rect 45888 7392 45894 7404
rect 46293 7395 46351 7401
rect 46293 7392 46305 7395
rect 45888 7364 46305 7392
rect 45888 7352 45894 7364
rect 46293 7361 46305 7364
rect 46339 7361 46351 7395
rect 47578 7392 47584 7404
rect 47539 7364 47584 7392
rect 46293 7355 46351 7361
rect 47578 7352 47584 7364
rect 47636 7352 47642 7404
rect 47670 7352 47676 7404
rect 47728 7392 47734 7404
rect 48225 7395 48283 7401
rect 48225 7392 48237 7395
rect 47728 7364 48237 7392
rect 47728 7352 47734 7364
rect 48225 7361 48237 7364
rect 48271 7361 48283 7395
rect 48866 7392 48872 7404
rect 48827 7364 48872 7392
rect 48225 7355 48283 7361
rect 48866 7352 48872 7364
rect 48924 7352 48930 7404
rect 50154 7392 50160 7404
rect 50115 7364 50160 7392
rect 50154 7352 50160 7364
rect 50212 7352 50218 7404
rect 50430 7352 50436 7404
rect 50488 7392 50494 7404
rect 50801 7395 50859 7401
rect 50801 7392 50813 7395
rect 50488 7364 50813 7392
rect 50488 7352 50494 7364
rect 50801 7361 50813 7364
rect 50847 7361 50859 7395
rect 51442 7392 51448 7404
rect 51403 7364 51448 7392
rect 50801 7355 50859 7361
rect 51442 7352 51448 7364
rect 51500 7352 51506 7404
rect 52178 7352 52184 7404
rect 52236 7392 52242 7404
rect 52733 7395 52791 7401
rect 52733 7392 52745 7395
rect 52236 7364 52745 7392
rect 52236 7352 52242 7364
rect 52733 7361 52745 7364
rect 52779 7361 52791 7395
rect 52733 7355 52791 7361
rect 53098 7352 53104 7404
rect 53156 7392 53162 7404
rect 53377 7395 53435 7401
rect 53377 7392 53389 7395
rect 53156 7364 53389 7392
rect 53156 7352 53162 7364
rect 53377 7361 53389 7364
rect 53423 7361 53435 7395
rect 53377 7355 53435 7361
rect 53466 7352 53472 7404
rect 53524 7392 53530 7404
rect 54021 7395 54079 7401
rect 54021 7392 54033 7395
rect 53524 7364 54033 7392
rect 53524 7352 53530 7364
rect 54021 7361 54033 7364
rect 54067 7361 54079 7395
rect 54021 7355 54079 7361
rect 55214 7352 55220 7404
rect 55272 7392 55278 7404
rect 55309 7395 55367 7401
rect 55309 7392 55321 7395
rect 55272 7364 55321 7392
rect 55272 7352 55278 7364
rect 55309 7361 55321 7364
rect 55355 7361 55367 7395
rect 55309 7355 55367 7361
rect 55490 7352 55496 7404
rect 55548 7392 55554 7404
rect 55953 7395 56011 7401
rect 55953 7392 55965 7395
rect 55548 7364 55965 7392
rect 55548 7352 55554 7364
rect 55953 7361 55965 7364
rect 55999 7361 56011 7395
rect 55953 7355 56011 7361
rect 56226 7352 56232 7404
rect 56284 7392 56290 7404
rect 56597 7395 56655 7401
rect 56597 7392 56609 7395
rect 56284 7364 56609 7392
rect 56284 7352 56290 7364
rect 56597 7361 56609 7364
rect 56643 7361 56655 7395
rect 56597 7355 56655 7361
rect 35250 7284 35256 7336
rect 35308 7324 35314 7336
rect 35989 7327 36047 7333
rect 35989 7324 36001 7327
rect 35308 7296 36001 7324
rect 35308 7284 35314 7296
rect 35989 7293 36001 7296
rect 36035 7293 36047 7327
rect 35989 7287 36047 7293
rect 42426 7216 42432 7268
rect 42484 7256 42490 7268
rect 43073 7259 43131 7265
rect 43073 7256 43085 7259
rect 42484 7228 43085 7256
rect 42484 7216 42490 7228
rect 43073 7225 43085 7228
rect 43119 7225 43131 7259
rect 43073 7219 43131 7225
rect 1104 7098 58880 7120
rect 1104 7046 8174 7098
rect 8226 7046 8238 7098
rect 8290 7046 8302 7098
rect 8354 7046 8366 7098
rect 8418 7046 8430 7098
rect 8482 7046 22622 7098
rect 22674 7046 22686 7098
rect 22738 7046 22750 7098
rect 22802 7046 22814 7098
rect 22866 7046 22878 7098
rect 22930 7046 37070 7098
rect 37122 7046 37134 7098
rect 37186 7046 37198 7098
rect 37250 7046 37262 7098
rect 37314 7046 37326 7098
rect 37378 7046 51518 7098
rect 51570 7046 51582 7098
rect 51634 7046 51646 7098
rect 51698 7046 51710 7098
rect 51762 7046 51774 7098
rect 51826 7046 58880 7098
rect 1104 7024 58880 7046
rect 6362 6848 6368 6860
rect 6323 6820 6368 6848
rect 6362 6808 6368 6820
rect 6420 6808 6426 6860
rect 11422 6848 11428 6860
rect 11383 6820 11428 6848
rect 11422 6808 11428 6820
rect 11480 6808 11486 6860
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 14148 6820 14197 6848
rect 14148 6808 14154 6820
rect 14185 6817 14197 6820
rect 14231 6817 14243 6851
rect 16942 6848 16948 6860
rect 16903 6820 16948 6848
rect 14185 6811 14243 6817
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 20990 6808 20996 6860
rect 21048 6848 21054 6860
rect 21085 6851 21143 6857
rect 21085 6848 21097 6851
rect 21048 6820 21097 6848
rect 21048 6808 21054 6820
rect 21085 6817 21097 6820
rect 21131 6817 21143 6851
rect 24394 6848 24400 6860
rect 24355 6820 24400 6848
rect 21085 6811 21143 6817
rect 24394 6808 24400 6820
rect 24452 6808 24458 6860
rect 26970 6808 26976 6860
rect 27028 6848 27034 6860
rect 27065 6851 27123 6857
rect 27065 6848 27077 6851
rect 27028 6820 27077 6848
rect 27028 6808 27034 6820
rect 27065 6817 27077 6820
rect 27111 6817 27123 6851
rect 36262 6848 36268 6860
rect 36223 6820 36268 6848
rect 27065 6811 27123 6817
rect 36262 6808 36268 6820
rect 36320 6808 36326 6860
rect 39390 6808 39396 6860
rect 39448 6848 39454 6860
rect 39853 6851 39911 6857
rect 39853 6848 39865 6851
rect 39448 6820 39865 6848
rect 39448 6808 39454 6820
rect 39853 6817 39865 6820
rect 39899 6817 39911 6851
rect 43622 6848 43628 6860
rect 43583 6820 43628 6848
rect 39853 6811 39911 6817
rect 43622 6808 43628 6820
rect 43680 6808 43686 6860
rect 46290 6808 46296 6860
rect 46348 6848 46354 6860
rect 46385 6851 46443 6857
rect 46385 6848 46397 6851
rect 46348 6820 46397 6848
rect 46348 6808 46354 6820
rect 46385 6817 46397 6820
rect 46431 6817 46443 6851
rect 46385 6811 46443 6817
rect 49050 6808 49056 6860
rect 49108 6848 49114 6860
rect 49145 6851 49203 6857
rect 49145 6848 49157 6851
rect 49108 6820 49157 6848
rect 49108 6808 49114 6820
rect 49145 6817 49157 6820
rect 49191 6817 49203 6851
rect 54202 6848 54208 6860
rect 54163 6820 54208 6848
rect 49145 6811 49203 6817
rect 54202 6808 54208 6820
rect 54260 6808 54266 6860
rect 26513 6715 26571 6721
rect 26513 6681 26525 6715
rect 26559 6712 26571 6715
rect 27338 6712 27344 6724
rect 26559 6684 27344 6712
rect 26559 6681 26571 6684
rect 26513 6675 26571 6681
rect 27338 6672 27344 6684
rect 27396 6712 27402 6724
rect 27801 6715 27859 6721
rect 27801 6712 27813 6715
rect 27396 6684 27813 6712
rect 27396 6672 27402 6684
rect 27801 6681 27813 6684
rect 27847 6712 27859 6715
rect 47026 6712 47032 6724
rect 27847 6684 47032 6712
rect 27847 6681 27859 6684
rect 27801 6675 27859 6681
rect 47026 6672 47032 6684
rect 47084 6712 47090 6724
rect 48130 6712 48136 6724
rect 47084 6684 48136 6712
rect 47084 6672 47090 6684
rect 48130 6672 48136 6684
rect 48188 6672 48194 6724
rect 9858 6604 9864 6656
rect 9916 6644 9922 6656
rect 9953 6647 10011 6653
rect 9953 6644 9965 6647
rect 9916 6616 9965 6644
rect 9916 6604 9922 6616
rect 9953 6613 9965 6616
rect 9999 6613 10011 6647
rect 33502 6644 33508 6656
rect 33463 6616 33508 6644
rect 9953 6607 10011 6613
rect 33502 6604 33508 6616
rect 33560 6604 33566 6656
rect 52178 6644 52184 6656
rect 52139 6616 52184 6644
rect 52178 6604 52184 6616
rect 52236 6604 52242 6656
rect 1104 6554 58880 6576
rect 1104 6502 15398 6554
rect 15450 6502 15462 6554
rect 15514 6502 15526 6554
rect 15578 6502 15590 6554
rect 15642 6502 15654 6554
rect 15706 6502 29846 6554
rect 29898 6502 29910 6554
rect 29962 6502 29974 6554
rect 30026 6502 30038 6554
rect 30090 6502 30102 6554
rect 30154 6502 44294 6554
rect 44346 6502 44358 6554
rect 44410 6502 44422 6554
rect 44474 6502 44486 6554
rect 44538 6502 44550 6554
rect 44602 6502 58880 6554
rect 1104 6480 58880 6502
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6236 8263 6239
rect 8662 6236 8668 6248
rect 8251 6208 8668 6236
rect 8251 6205 8263 6208
rect 8205 6199 8263 6205
rect 8662 6196 8668 6208
rect 8720 6196 8726 6248
rect 20717 6239 20775 6245
rect 20717 6205 20729 6239
rect 20763 6236 20775 6239
rect 20806 6236 20812 6248
rect 20763 6208 20812 6236
rect 20763 6205 20775 6208
rect 20717 6199 20775 6205
rect 20806 6196 20812 6208
rect 20864 6196 20870 6248
rect 30282 6196 30288 6248
rect 30340 6236 30346 6248
rect 30340 6208 33456 6236
rect 30340 6196 30346 6208
rect 9858 6128 9864 6180
rect 9916 6168 9922 6180
rect 11885 6171 11943 6177
rect 11885 6168 11897 6171
rect 9916 6140 11897 6168
rect 9916 6128 9922 6140
rect 11885 6137 11897 6140
rect 11931 6137 11943 6171
rect 11885 6131 11943 6137
rect 8754 6100 8760 6112
rect 8715 6072 8760 6100
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 9306 6100 9312 6112
rect 9267 6072 9312 6100
rect 9306 6060 9312 6072
rect 9364 6060 9370 6112
rect 9490 6060 9496 6112
rect 9548 6100 9554 6112
rect 9769 6103 9827 6109
rect 9769 6100 9781 6103
rect 9548 6072 9781 6100
rect 9548 6060 9554 6072
rect 9769 6069 9781 6072
rect 9815 6069 9827 6103
rect 10502 6100 10508 6112
rect 10463 6072 10508 6100
rect 9769 6063 9827 6069
rect 10502 6060 10508 6072
rect 10560 6060 10566 6112
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 21177 6103 21235 6109
rect 21177 6100 21189 6103
rect 20772 6072 21189 6100
rect 20772 6060 20778 6072
rect 21177 6069 21189 6072
rect 21223 6069 21235 6103
rect 23290 6100 23296 6112
rect 23251 6072 23296 6100
rect 21177 6063 21235 6069
rect 23290 6060 23296 6072
rect 23348 6060 23354 6112
rect 25130 6060 25136 6112
rect 25188 6100 25194 6112
rect 25685 6103 25743 6109
rect 25685 6100 25697 6103
rect 25188 6072 25697 6100
rect 25188 6060 25194 6072
rect 25685 6069 25697 6072
rect 25731 6100 25743 6103
rect 26329 6103 26387 6109
rect 26329 6100 26341 6103
rect 25731 6072 26341 6100
rect 25731 6069 25743 6072
rect 25685 6063 25743 6069
rect 26329 6069 26341 6072
rect 26375 6100 26387 6103
rect 26970 6100 26976 6112
rect 26375 6072 26976 6100
rect 26375 6069 26387 6072
rect 26329 6063 26387 6069
rect 26970 6060 26976 6072
rect 27028 6060 27034 6112
rect 27985 6103 28043 6109
rect 27985 6069 27997 6103
rect 28031 6100 28043 6103
rect 28258 6100 28264 6112
rect 28031 6072 28264 6100
rect 28031 6069 28043 6072
rect 27985 6063 28043 6069
rect 28258 6060 28264 6072
rect 28316 6060 28322 6112
rect 30466 6100 30472 6112
rect 30427 6072 30472 6100
rect 30466 6060 30472 6072
rect 30524 6060 30530 6112
rect 31021 6103 31079 6109
rect 31021 6069 31033 6103
rect 31067 6100 31079 6103
rect 31754 6100 31760 6112
rect 31067 6072 31760 6100
rect 31067 6069 31079 6072
rect 31021 6063 31079 6069
rect 31754 6060 31760 6072
rect 31812 6060 31818 6112
rect 33226 6100 33232 6112
rect 33187 6072 33232 6100
rect 33226 6060 33232 6072
rect 33284 6060 33290 6112
rect 33428 6100 33456 6208
rect 38378 6196 38384 6248
rect 38436 6236 38442 6248
rect 42978 6236 42984 6248
rect 38436 6208 42984 6236
rect 38436 6196 38442 6208
rect 42978 6196 42984 6208
rect 43036 6196 43042 6248
rect 33502 6128 33508 6180
rect 33560 6168 33566 6180
rect 33873 6171 33931 6177
rect 33873 6168 33885 6171
rect 33560 6140 33885 6168
rect 33560 6128 33566 6140
rect 33873 6137 33885 6140
rect 33919 6168 33931 6171
rect 33919 6140 35756 6168
rect 33919 6137 33931 6140
rect 33873 6131 33931 6137
rect 35728 6112 35756 6140
rect 40034 6128 40040 6180
rect 40092 6168 40098 6180
rect 50525 6171 50583 6177
rect 50525 6168 50537 6171
rect 40092 6140 50537 6168
rect 40092 6128 40098 6140
rect 50525 6137 50537 6140
rect 50571 6168 50583 6171
rect 50890 6168 50896 6180
rect 50571 6140 50896 6168
rect 50571 6137 50583 6140
rect 50525 6131 50583 6137
rect 50890 6128 50896 6140
rect 50948 6128 50954 6180
rect 34606 6100 34612 6112
rect 33428 6072 34612 6100
rect 34606 6060 34612 6072
rect 34664 6060 34670 6112
rect 35066 6100 35072 6112
rect 35027 6072 35072 6100
rect 35066 6060 35072 6072
rect 35124 6060 35130 6112
rect 35710 6100 35716 6112
rect 35671 6072 35716 6100
rect 35710 6060 35716 6072
rect 35768 6060 35774 6112
rect 35802 6060 35808 6112
rect 35860 6100 35866 6112
rect 36262 6100 36268 6112
rect 35860 6072 36268 6100
rect 35860 6060 35866 6072
rect 36262 6060 36268 6072
rect 36320 6100 36326 6112
rect 39758 6100 39764 6112
rect 36320 6072 39764 6100
rect 36320 6060 36326 6072
rect 39758 6060 39764 6072
rect 39816 6060 39822 6112
rect 45554 6100 45560 6112
rect 45515 6072 45560 6100
rect 45554 6060 45560 6072
rect 45612 6060 45618 6112
rect 46934 6060 46940 6112
rect 46992 6100 46998 6112
rect 49881 6103 49939 6109
rect 49881 6100 49893 6103
rect 46992 6072 49893 6100
rect 46992 6060 46998 6072
rect 49881 6069 49893 6072
rect 49927 6069 49939 6103
rect 49881 6063 49939 6069
rect 51169 6103 51227 6109
rect 51169 6069 51181 6103
rect 51215 6100 51227 6103
rect 51350 6100 51356 6112
rect 51215 6072 51356 6100
rect 51215 6069 51227 6072
rect 51169 6063 51227 6069
rect 51350 6060 51356 6072
rect 51408 6060 51414 6112
rect 51905 6103 51963 6109
rect 51905 6069 51917 6103
rect 51951 6100 51963 6103
rect 51994 6100 52000 6112
rect 51951 6072 52000 6100
rect 51951 6069 51963 6072
rect 51905 6063 51963 6069
rect 51994 6060 52000 6072
rect 52052 6100 52058 6112
rect 52733 6103 52791 6109
rect 52733 6100 52745 6103
rect 52052 6072 52745 6100
rect 52052 6060 52058 6072
rect 52733 6069 52745 6072
rect 52779 6069 52791 6103
rect 52733 6063 52791 6069
rect 1104 6010 58880 6032
rect 1104 5958 8174 6010
rect 8226 5958 8238 6010
rect 8290 5958 8302 6010
rect 8354 5958 8366 6010
rect 8418 5958 8430 6010
rect 8482 5958 22622 6010
rect 22674 5958 22686 6010
rect 22738 5958 22750 6010
rect 22802 5958 22814 6010
rect 22866 5958 22878 6010
rect 22930 5958 37070 6010
rect 37122 5958 37134 6010
rect 37186 5958 37198 6010
rect 37250 5958 37262 6010
rect 37314 5958 37326 6010
rect 37378 5958 51518 6010
rect 51570 5958 51582 6010
rect 51634 5958 51646 6010
rect 51698 5958 51710 6010
rect 51762 5958 51774 6010
rect 51826 5958 58880 6010
rect 1104 5936 58880 5958
rect 4801 5899 4859 5905
rect 4801 5865 4813 5899
rect 4847 5896 4859 5899
rect 5442 5896 5448 5908
rect 4847 5868 5448 5896
rect 4847 5865 4859 5868
rect 4801 5859 4859 5865
rect 5442 5856 5448 5868
rect 5500 5896 5506 5908
rect 10502 5896 10508 5908
rect 5500 5868 10508 5896
rect 5500 5856 5506 5868
rect 10502 5856 10508 5868
rect 10560 5896 10566 5908
rect 20806 5896 20812 5908
rect 10560 5868 20812 5896
rect 10560 5856 10566 5868
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 31846 5856 31852 5908
rect 31904 5896 31910 5908
rect 33042 5896 33048 5908
rect 31904 5868 33048 5896
rect 31904 5856 31910 5868
rect 33042 5856 33048 5868
rect 33100 5856 33106 5908
rect 34698 5896 34704 5908
rect 34659 5868 34704 5896
rect 34698 5856 34704 5868
rect 34756 5896 34762 5908
rect 35526 5896 35532 5908
rect 34756 5868 35532 5896
rect 34756 5856 34762 5868
rect 35526 5856 35532 5868
rect 35584 5856 35590 5908
rect 35710 5856 35716 5908
rect 35768 5896 35774 5908
rect 40497 5899 40555 5905
rect 40497 5896 40509 5899
rect 35768 5868 40509 5896
rect 35768 5856 35774 5868
rect 40497 5865 40509 5868
rect 40543 5896 40555 5899
rect 41690 5896 41696 5908
rect 40543 5868 41696 5896
rect 40543 5865 40555 5868
rect 40497 5859 40555 5865
rect 41690 5856 41696 5868
rect 41748 5856 41754 5908
rect 42613 5899 42671 5905
rect 42613 5865 42625 5899
rect 42659 5896 42671 5899
rect 42978 5896 42984 5908
rect 42659 5868 42984 5896
rect 42659 5865 42671 5868
rect 42613 5859 42671 5865
rect 42978 5856 42984 5868
rect 43036 5896 43042 5908
rect 49786 5896 49792 5908
rect 43036 5868 49792 5896
rect 43036 5856 43042 5868
rect 49786 5856 49792 5868
rect 49844 5856 49850 5908
rect 52178 5856 52184 5908
rect 52236 5896 52242 5908
rect 53653 5899 53711 5905
rect 53653 5896 53665 5899
rect 52236 5868 53665 5896
rect 52236 5856 52242 5868
rect 53653 5865 53665 5868
rect 53699 5865 53711 5899
rect 53653 5859 53711 5865
rect 4338 5788 4344 5840
rect 4396 5828 4402 5840
rect 26421 5831 26479 5837
rect 4396 5800 12434 5828
rect 4396 5788 4402 5800
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 7834 5760 7840 5772
rect 7239 5732 7840 5760
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5692 7803 5695
rect 8018 5692 8024 5704
rect 7791 5664 8024 5692
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 8018 5652 8024 5664
rect 8076 5692 8082 5704
rect 8389 5695 8447 5701
rect 8389 5692 8401 5695
rect 8076 5664 8401 5692
rect 8076 5652 8082 5664
rect 8389 5661 8401 5664
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 9401 5695 9459 5701
rect 9401 5692 9413 5695
rect 9364 5664 9413 5692
rect 9364 5652 9370 5664
rect 9401 5661 9413 5664
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 10042 5652 10048 5704
rect 10100 5692 10106 5704
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 10100 5664 10149 5692
rect 10100 5652 10106 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10870 5652 10876 5704
rect 10928 5692 10934 5704
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 10928 5664 10977 5692
rect 10928 5652 10934 5664
rect 10965 5661 10977 5664
rect 11011 5661 11023 5695
rect 12066 5692 12072 5704
rect 12027 5664 12072 5692
rect 10965 5655 11023 5661
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 4154 5584 4160 5636
rect 4212 5624 4218 5636
rect 5905 5627 5963 5633
rect 5905 5624 5917 5627
rect 4212 5596 5917 5624
rect 4212 5584 4218 5596
rect 5905 5593 5917 5596
rect 5951 5624 5963 5627
rect 6457 5627 6515 5633
rect 6457 5624 6469 5627
rect 5951 5596 6469 5624
rect 5951 5593 5963 5596
rect 5905 5587 5963 5593
rect 6457 5593 6469 5596
rect 6503 5624 6515 5627
rect 9858 5624 9864 5636
rect 6503 5596 9864 5624
rect 6503 5593 6515 5596
rect 6457 5587 6515 5593
rect 9858 5584 9864 5596
rect 9916 5584 9922 5636
rect 12406 5624 12434 5800
rect 26421 5797 26433 5831
rect 26467 5828 26479 5831
rect 27706 5828 27712 5840
rect 26467 5800 27712 5828
rect 26467 5797 26479 5800
rect 26421 5791 26479 5797
rect 27706 5788 27712 5800
rect 27764 5788 27770 5840
rect 30929 5831 30987 5837
rect 30929 5797 30941 5831
rect 30975 5797 30987 5831
rect 30929 5791 30987 5797
rect 27614 5720 27620 5772
rect 27672 5760 27678 5772
rect 28169 5763 28227 5769
rect 28169 5760 28181 5763
rect 27672 5732 28181 5760
rect 27672 5720 27678 5732
rect 28169 5729 28181 5732
rect 28215 5729 28227 5763
rect 30944 5760 30972 5791
rect 31018 5788 31024 5840
rect 31076 5828 31082 5840
rect 31076 5800 31121 5828
rect 31076 5788 31082 5800
rect 34606 5788 34612 5840
rect 34664 5828 34670 5840
rect 48130 5828 48136 5840
rect 34664 5800 45324 5828
rect 48091 5800 48136 5828
rect 34664 5788 34670 5800
rect 31662 5760 31668 5772
rect 30944 5732 31064 5760
rect 31623 5732 31668 5760
rect 28169 5723 28227 5729
rect 12802 5652 12808 5704
rect 12860 5692 12866 5704
rect 12897 5695 12955 5701
rect 12897 5692 12909 5695
rect 12860 5664 12909 5692
rect 12860 5652 12866 5664
rect 12897 5661 12909 5664
rect 12943 5661 12955 5695
rect 12897 5655 12955 5661
rect 14734 5652 14740 5704
rect 14792 5692 14798 5704
rect 14829 5695 14887 5701
rect 14829 5692 14841 5695
rect 14792 5664 14841 5692
rect 14792 5652 14798 5664
rect 14829 5661 14841 5664
rect 14875 5661 14887 5695
rect 14829 5655 14887 5661
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5692 15899 5695
rect 16206 5692 16212 5704
rect 15887 5664 16212 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 16206 5652 16212 5664
rect 16264 5692 16270 5704
rect 16485 5695 16543 5701
rect 16485 5692 16497 5695
rect 16264 5664 16497 5692
rect 16264 5652 16270 5664
rect 16485 5661 16497 5664
rect 16531 5661 16543 5695
rect 16485 5655 16543 5661
rect 16942 5652 16948 5704
rect 17000 5692 17006 5704
rect 17037 5695 17095 5701
rect 17037 5692 17049 5695
rect 17000 5664 17049 5692
rect 17000 5652 17006 5664
rect 17037 5661 17049 5664
rect 17083 5661 17095 5695
rect 17037 5655 17095 5661
rect 26786 5652 26792 5704
rect 26844 5692 26850 5704
rect 26881 5695 26939 5701
rect 26881 5692 26893 5695
rect 26844 5664 26893 5692
rect 26844 5652 26850 5664
rect 26881 5661 26893 5664
rect 26927 5661 26939 5695
rect 26881 5655 26939 5661
rect 27709 5695 27767 5701
rect 27709 5661 27721 5695
rect 27755 5692 27767 5695
rect 29730 5692 29736 5704
rect 27755 5664 29736 5692
rect 27755 5661 27767 5664
rect 27709 5655 27767 5661
rect 29730 5652 29736 5664
rect 29788 5652 29794 5704
rect 30929 5695 30987 5701
rect 30929 5692 30941 5695
rect 30392 5664 30941 5692
rect 22738 5624 22744 5636
rect 12406 5596 22744 5624
rect 22738 5584 22744 5596
rect 22796 5584 22802 5636
rect 30392 5568 30420 5664
rect 30929 5661 30941 5664
rect 30975 5661 30987 5695
rect 31036 5692 31064 5732
rect 31662 5720 31668 5732
rect 31720 5720 31726 5772
rect 32048 5732 32628 5760
rect 31757 5695 31815 5701
rect 31757 5692 31769 5695
rect 31036 5664 31769 5692
rect 30929 5655 30987 5661
rect 31757 5661 31769 5664
rect 31803 5661 31815 5695
rect 31757 5655 31815 5661
rect 31941 5695 31999 5701
rect 31941 5661 31953 5695
rect 31987 5686 31999 5695
rect 32048 5686 32076 5732
rect 31987 5661 32076 5686
rect 31941 5658 32076 5661
rect 31941 5655 31999 5658
rect 7742 5516 7748 5568
rect 7800 5556 7806 5568
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 7800 5528 8217 5556
rect 7800 5516 7806 5528
rect 8205 5525 8217 5528
rect 8251 5525 8263 5559
rect 8205 5519 8263 5525
rect 9585 5559 9643 5565
rect 9585 5525 9597 5559
rect 9631 5556 9643 5559
rect 12894 5556 12900 5568
rect 9631 5528 12900 5556
rect 9631 5525 9643 5528
rect 9585 5519 9643 5525
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 14366 5556 14372 5568
rect 14327 5528 14372 5556
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 16298 5556 16304 5568
rect 16259 5528 16304 5556
rect 16298 5516 16304 5528
rect 16356 5516 16362 5568
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 20073 5559 20131 5565
rect 20073 5556 20085 5559
rect 20036 5528 20085 5556
rect 20036 5516 20042 5528
rect 20073 5525 20085 5528
rect 20119 5525 20131 5559
rect 20714 5556 20720 5568
rect 20675 5528 20720 5556
rect 20073 5519 20131 5525
rect 20714 5516 20720 5528
rect 20772 5516 20778 5568
rect 21545 5559 21603 5565
rect 21545 5525 21557 5559
rect 21591 5556 21603 5559
rect 21634 5556 21640 5568
rect 21591 5528 21640 5556
rect 21591 5525 21603 5528
rect 21545 5519 21603 5525
rect 21634 5516 21640 5528
rect 21692 5516 21698 5568
rect 22373 5559 22431 5565
rect 22373 5525 22385 5559
rect 22419 5556 22431 5559
rect 22462 5556 22468 5568
rect 22419 5528 22468 5556
rect 22419 5525 22431 5528
rect 22373 5519 22431 5525
rect 22462 5516 22468 5528
rect 22520 5516 22526 5568
rect 22925 5559 22983 5565
rect 22925 5525 22937 5559
rect 22971 5556 22983 5559
rect 23014 5556 23020 5568
rect 22971 5528 23020 5556
rect 22971 5525 22983 5528
rect 22925 5519 22983 5525
rect 23014 5516 23020 5528
rect 23072 5516 23078 5568
rect 23474 5556 23480 5568
rect 23435 5528 23480 5556
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 24673 5559 24731 5565
rect 24673 5525 24685 5559
rect 24719 5556 24731 5559
rect 24762 5556 24768 5568
rect 24719 5528 24768 5556
rect 24719 5525 24731 5528
rect 24673 5519 24731 5525
rect 24762 5516 24768 5528
rect 24820 5516 24826 5568
rect 25130 5556 25136 5568
rect 25091 5528 25136 5556
rect 25130 5516 25136 5528
rect 25188 5516 25194 5568
rect 25222 5516 25228 5568
rect 25280 5556 25286 5568
rect 25777 5559 25835 5565
rect 25777 5556 25789 5559
rect 25280 5528 25789 5556
rect 25280 5516 25286 5528
rect 25777 5525 25789 5528
rect 25823 5556 25835 5559
rect 26694 5556 26700 5568
rect 25823 5528 26700 5556
rect 25823 5525 25835 5528
rect 25777 5519 25835 5525
rect 26694 5516 26700 5528
rect 26752 5516 26758 5568
rect 26878 5516 26884 5568
rect 26936 5556 26942 5568
rect 27525 5559 27583 5565
rect 27525 5556 27537 5559
rect 26936 5528 27537 5556
rect 26936 5516 26942 5528
rect 27525 5525 27537 5528
rect 27571 5525 27583 5559
rect 28810 5556 28816 5568
rect 28771 5528 28816 5556
rect 27525 5519 27583 5525
rect 28810 5516 28816 5528
rect 28868 5516 28874 5568
rect 29454 5516 29460 5568
rect 29512 5556 29518 5568
rect 29733 5559 29791 5565
rect 29733 5556 29745 5559
rect 29512 5528 29745 5556
rect 29512 5516 29518 5528
rect 29733 5525 29745 5528
rect 29779 5525 29791 5559
rect 30374 5556 30380 5568
rect 30335 5528 30380 5556
rect 29733 5519 29791 5525
rect 30374 5516 30380 5528
rect 30432 5516 30438 5568
rect 30944 5556 30972 5655
rect 31205 5627 31263 5633
rect 31205 5593 31217 5627
rect 31251 5624 31263 5627
rect 31846 5624 31852 5636
rect 31251 5596 31852 5624
rect 31251 5593 31263 5596
rect 31205 5587 31263 5593
rect 31846 5584 31852 5596
rect 31904 5584 31910 5636
rect 32122 5624 32128 5636
rect 32083 5596 32128 5624
rect 32122 5584 32128 5596
rect 32180 5584 32186 5636
rect 32600 5624 32628 5732
rect 33042 5720 33048 5772
rect 33100 5760 33106 5772
rect 34882 5760 34888 5772
rect 33100 5732 34888 5760
rect 33100 5720 33106 5732
rect 34882 5720 34888 5732
rect 34940 5720 34946 5772
rect 35176 5760 35204 5800
rect 35253 5763 35311 5769
rect 35253 5760 35265 5763
rect 35176 5732 35265 5760
rect 35253 5729 35265 5732
rect 35299 5729 35311 5763
rect 35802 5760 35808 5772
rect 35253 5723 35311 5729
rect 35452 5732 35808 5760
rect 32858 5652 32864 5704
rect 32916 5692 32922 5704
rect 33413 5695 33471 5701
rect 33413 5692 33425 5695
rect 32916 5664 33425 5692
rect 32916 5652 32922 5664
rect 33413 5661 33425 5664
rect 33459 5661 33471 5695
rect 33413 5655 33471 5661
rect 33505 5695 33563 5701
rect 33505 5661 33517 5695
rect 33551 5692 33563 5695
rect 34146 5692 34152 5704
rect 33551 5664 34152 5692
rect 33551 5661 33563 5664
rect 33505 5655 33563 5661
rect 34146 5652 34152 5664
rect 34204 5652 34210 5704
rect 35452 5692 35480 5732
rect 35802 5720 35808 5732
rect 35860 5720 35866 5772
rect 37553 5763 37611 5769
rect 37553 5760 37565 5763
rect 36096 5732 37565 5760
rect 35268 5664 35480 5692
rect 32677 5627 32735 5633
rect 32677 5624 32689 5627
rect 32600 5596 32689 5624
rect 32677 5593 32689 5596
rect 32723 5624 32735 5627
rect 33689 5627 33747 5633
rect 32723 5596 33640 5624
rect 32723 5593 32735 5596
rect 32677 5587 32735 5593
rect 32030 5556 32036 5568
rect 30944 5528 32036 5556
rect 32030 5516 32036 5528
rect 32088 5516 32094 5568
rect 33410 5556 33416 5568
rect 33371 5528 33416 5556
rect 33410 5516 33416 5528
rect 33468 5516 33474 5568
rect 33612 5556 33640 5596
rect 33689 5593 33701 5627
rect 33735 5624 33747 5627
rect 35268 5624 35296 5664
rect 35526 5652 35532 5704
rect 35584 5692 35590 5704
rect 35713 5695 35771 5701
rect 35713 5692 35725 5695
rect 35584 5664 35725 5692
rect 35584 5652 35590 5664
rect 35713 5661 35725 5664
rect 35759 5692 35771 5695
rect 35759 5686 35848 5692
rect 36096 5686 36124 5732
rect 37553 5729 37565 5732
rect 37599 5729 37611 5763
rect 37553 5723 37611 5729
rect 37645 5763 37703 5769
rect 37645 5729 37657 5763
rect 37691 5760 37703 5763
rect 40126 5760 40132 5772
rect 37691 5732 40132 5760
rect 37691 5729 37703 5732
rect 37645 5723 37703 5729
rect 36262 5692 36268 5704
rect 35759 5664 36124 5686
rect 36223 5664 36268 5692
rect 35759 5661 35771 5664
rect 35713 5655 35771 5661
rect 35820 5658 36124 5664
rect 36262 5652 36268 5664
rect 36320 5652 36326 5704
rect 36446 5692 36452 5704
rect 36407 5664 36452 5692
rect 36446 5652 36452 5664
rect 36504 5692 36510 5704
rect 37277 5695 37335 5701
rect 37277 5692 37289 5695
rect 36504 5664 37289 5692
rect 36504 5652 36510 5664
rect 37277 5661 37289 5664
rect 37323 5661 37335 5695
rect 37568 5692 37596 5723
rect 40126 5720 40132 5732
rect 40184 5720 40190 5772
rect 45296 5760 45324 5800
rect 48130 5788 48136 5800
rect 48188 5788 48194 5840
rect 45925 5763 45983 5769
rect 45925 5760 45937 5763
rect 45296 5732 45937 5760
rect 38197 5695 38255 5701
rect 38197 5692 38209 5695
rect 37568 5664 38209 5692
rect 37277 5655 37335 5661
rect 38197 5661 38209 5664
rect 38243 5692 38255 5695
rect 42794 5692 42800 5704
rect 38243 5664 42800 5692
rect 38243 5661 38255 5664
rect 38197 5655 38255 5661
rect 33735 5596 35296 5624
rect 33735 5593 33747 5596
rect 33689 5587 33747 5593
rect 35342 5584 35348 5636
rect 35400 5624 35406 5636
rect 36357 5627 36415 5633
rect 36357 5624 36369 5627
rect 35400 5596 36369 5624
rect 35400 5584 35406 5596
rect 36357 5593 36369 5596
rect 36403 5593 36415 5627
rect 37292 5624 37320 5655
rect 42794 5652 42800 5664
rect 42852 5692 42858 5704
rect 45296 5701 45324 5732
rect 45925 5729 45937 5732
rect 45971 5729 45983 5763
rect 45925 5723 45983 5729
rect 52270 5720 52276 5772
rect 52328 5760 52334 5772
rect 53009 5763 53067 5769
rect 53009 5760 53021 5763
rect 52328 5732 53021 5760
rect 52328 5720 52334 5732
rect 53009 5729 53021 5732
rect 53055 5729 53067 5763
rect 53009 5723 53067 5729
rect 43073 5695 43131 5701
rect 43073 5692 43085 5695
rect 42852 5664 43085 5692
rect 42852 5652 42858 5664
rect 43073 5661 43085 5664
rect 43119 5661 43131 5695
rect 43073 5655 43131 5661
rect 45281 5695 45339 5701
rect 45281 5661 45293 5695
rect 45327 5661 45339 5695
rect 45281 5655 45339 5661
rect 45465 5695 45523 5701
rect 45465 5661 45477 5695
rect 45511 5692 45523 5695
rect 45554 5692 45560 5704
rect 45511 5664 45560 5692
rect 45511 5661 45523 5664
rect 45465 5655 45523 5661
rect 39850 5624 39856 5636
rect 37292 5596 39856 5624
rect 36357 5587 36415 5593
rect 39850 5584 39856 5596
rect 39908 5584 39914 5636
rect 39945 5627 40003 5633
rect 39945 5593 39957 5627
rect 39991 5624 40003 5627
rect 40034 5624 40040 5636
rect 39991 5596 40040 5624
rect 39991 5593 40003 5596
rect 39945 5587 40003 5593
rect 35069 5559 35127 5565
rect 35069 5556 35081 5559
rect 33612 5528 35081 5556
rect 35069 5525 35081 5528
rect 35115 5556 35127 5559
rect 39960 5556 39988 5587
rect 40034 5584 40040 5596
rect 40092 5624 40098 5636
rect 40494 5624 40500 5636
rect 40092 5596 40500 5624
rect 40092 5584 40098 5596
rect 40494 5584 40500 5596
rect 40552 5584 40558 5636
rect 43088 5624 43116 5655
rect 45480 5624 45508 5655
rect 45554 5652 45560 5664
rect 45612 5652 45618 5704
rect 50246 5652 50252 5704
rect 50304 5692 50310 5704
rect 50341 5695 50399 5701
rect 50341 5692 50353 5695
rect 50304 5664 50353 5692
rect 50304 5652 50310 5664
rect 50341 5661 50353 5664
rect 50387 5661 50399 5695
rect 50341 5655 50399 5661
rect 50522 5652 50528 5704
rect 50580 5692 50586 5704
rect 50985 5695 51043 5701
rect 50985 5692 50997 5695
rect 50580 5664 50997 5692
rect 50580 5652 50586 5664
rect 50985 5661 50997 5664
rect 51031 5661 51043 5695
rect 50985 5655 51043 5661
rect 51442 5652 51448 5704
rect 51500 5692 51506 5704
rect 51721 5695 51779 5701
rect 51721 5692 51733 5695
rect 51500 5664 51733 5692
rect 51500 5652 51506 5664
rect 51721 5661 51733 5664
rect 51767 5661 51779 5695
rect 51721 5655 51779 5661
rect 51902 5652 51908 5704
rect 51960 5692 51966 5704
rect 52365 5695 52423 5701
rect 52365 5692 52377 5695
rect 51960 5664 52377 5692
rect 51960 5652 51966 5664
rect 52365 5661 52377 5664
rect 52411 5661 52423 5695
rect 52365 5655 52423 5661
rect 47581 5627 47639 5633
rect 47581 5624 47593 5627
rect 43088 5596 45508 5624
rect 46492 5596 47593 5624
rect 35115 5528 39988 5556
rect 41693 5559 41751 5565
rect 35115 5525 35127 5528
rect 35069 5519 35127 5525
rect 41693 5525 41705 5559
rect 41739 5556 41751 5559
rect 43070 5556 43076 5568
rect 41739 5528 43076 5556
rect 41739 5525 41751 5528
rect 41693 5519 41751 5525
rect 43070 5516 43076 5528
rect 43128 5516 43134 5568
rect 45186 5516 45192 5568
rect 45244 5556 45250 5568
rect 45373 5559 45431 5565
rect 45373 5556 45385 5559
rect 45244 5528 45385 5556
rect 45244 5516 45250 5528
rect 45373 5525 45385 5528
rect 45419 5525 45431 5559
rect 45373 5519 45431 5525
rect 46014 5516 46020 5568
rect 46072 5556 46078 5568
rect 46492 5565 46520 5596
rect 47581 5593 47593 5596
rect 47627 5624 47639 5627
rect 49694 5624 49700 5636
rect 47627 5596 49700 5624
rect 47627 5593 47639 5596
rect 47581 5587 47639 5593
rect 49694 5584 49700 5596
rect 49752 5584 49758 5636
rect 54754 5584 54760 5636
rect 54812 5624 54818 5636
rect 55861 5627 55919 5633
rect 55861 5624 55873 5627
rect 54812 5596 55873 5624
rect 54812 5584 54818 5596
rect 55861 5593 55873 5596
rect 55907 5593 55919 5627
rect 55861 5587 55919 5593
rect 46477 5559 46535 5565
rect 46477 5556 46489 5559
rect 46072 5528 46489 5556
rect 46072 5516 46078 5528
rect 46477 5525 46489 5528
rect 46523 5525 46535 5559
rect 46477 5519 46535 5525
rect 46934 5516 46940 5568
rect 46992 5556 46998 5568
rect 47029 5559 47087 5565
rect 47029 5556 47041 5559
rect 46992 5528 47041 5556
rect 46992 5516 46998 5528
rect 47029 5525 47041 5528
rect 47075 5525 47087 5559
rect 47029 5519 47087 5525
rect 49605 5559 49663 5565
rect 49605 5525 49617 5559
rect 49651 5556 49663 5559
rect 49786 5556 49792 5568
rect 49651 5528 49792 5556
rect 49651 5525 49663 5528
rect 49605 5519 49663 5525
rect 49786 5516 49792 5528
rect 49844 5516 49850 5568
rect 55214 5516 55220 5568
rect 55272 5556 55278 5568
rect 55309 5559 55367 5565
rect 55309 5556 55321 5559
rect 55272 5528 55321 5556
rect 55272 5516 55278 5528
rect 55309 5525 55321 5528
rect 55355 5525 55367 5559
rect 55309 5519 55367 5525
rect 1104 5466 58880 5488
rect 1104 5414 15398 5466
rect 15450 5414 15462 5466
rect 15514 5414 15526 5466
rect 15578 5414 15590 5466
rect 15642 5414 15654 5466
rect 15706 5414 29846 5466
rect 29898 5414 29910 5466
rect 29962 5414 29974 5466
rect 30026 5414 30038 5466
rect 30090 5414 30102 5466
rect 30154 5414 44294 5466
rect 44346 5414 44358 5466
rect 44410 5414 44422 5466
rect 44474 5414 44486 5466
rect 44538 5414 44550 5466
rect 44602 5414 58880 5466
rect 1104 5392 58880 5414
rect 4338 5352 4344 5364
rect 4299 5324 4344 5352
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 5442 5312 5448 5364
rect 5500 5352 5506 5364
rect 7561 5355 7619 5361
rect 7561 5352 7573 5355
rect 5500 5324 7573 5352
rect 5500 5312 5506 5324
rect 7561 5321 7573 5324
rect 7607 5321 7619 5355
rect 7561 5315 7619 5321
rect 9858 5312 9864 5364
rect 9916 5352 9922 5364
rect 19242 5352 19248 5364
rect 9916 5324 19248 5352
rect 9916 5312 9922 5324
rect 19242 5312 19248 5324
rect 19300 5352 19306 5364
rect 20714 5352 20720 5364
rect 19300 5324 20720 5352
rect 19300 5312 19306 5324
rect 20714 5312 20720 5324
rect 20772 5352 20778 5364
rect 23845 5355 23903 5361
rect 23845 5352 23857 5355
rect 20772 5324 23857 5352
rect 20772 5312 20778 5324
rect 23845 5321 23857 5324
rect 23891 5352 23903 5355
rect 24118 5352 24124 5364
rect 23891 5324 24124 5352
rect 23891 5321 23903 5324
rect 23845 5315 23903 5321
rect 24118 5312 24124 5324
rect 24176 5352 24182 5364
rect 25130 5352 25136 5364
rect 24176 5324 25136 5352
rect 24176 5312 24182 5324
rect 25130 5312 25136 5324
rect 25188 5312 25194 5364
rect 25774 5312 25780 5364
rect 25832 5352 25838 5364
rect 28353 5355 28411 5361
rect 28353 5352 28365 5355
rect 25832 5324 28365 5352
rect 25832 5312 25838 5324
rect 28353 5321 28365 5324
rect 28399 5352 28411 5355
rect 29546 5352 29552 5364
rect 28399 5324 29552 5352
rect 28399 5321 28411 5324
rect 28353 5315 28411 5321
rect 29546 5312 29552 5324
rect 29604 5312 29610 5364
rect 31018 5312 31024 5364
rect 31076 5352 31082 5364
rect 31297 5355 31355 5361
rect 31297 5352 31309 5355
rect 31076 5324 31309 5352
rect 31076 5312 31082 5324
rect 31297 5321 31309 5324
rect 31343 5321 31355 5355
rect 35161 5355 35219 5361
rect 31297 5315 31355 5321
rect 32324 5324 35112 5352
rect 6270 5284 6276 5296
rect 4264 5256 6276 5284
rect 4264 5225 4292 5256
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 6546 5244 6552 5296
rect 6604 5284 6610 5296
rect 12710 5284 12716 5296
rect 6604 5256 12716 5284
rect 6604 5244 6610 5256
rect 12710 5244 12716 5256
rect 12768 5244 12774 5296
rect 13446 5284 13452 5296
rect 13407 5256 13452 5284
rect 13446 5244 13452 5256
rect 13504 5244 13510 5296
rect 18322 5244 18328 5296
rect 18380 5284 18386 5296
rect 19061 5287 19119 5293
rect 19061 5284 19073 5287
rect 18380 5256 19073 5284
rect 18380 5244 18386 5256
rect 19061 5253 19073 5256
rect 19107 5253 19119 5287
rect 19061 5247 19119 5253
rect 20806 5244 20812 5296
rect 20864 5284 20870 5296
rect 21174 5284 21180 5296
rect 20864 5256 21180 5284
rect 20864 5244 20870 5256
rect 21174 5244 21180 5256
rect 21232 5244 21238 5296
rect 22738 5284 22744 5296
rect 22699 5256 22744 5284
rect 22738 5244 22744 5256
rect 22796 5284 22802 5296
rect 23382 5284 23388 5296
rect 22796 5256 23388 5284
rect 22796 5244 22802 5256
rect 23382 5244 23388 5256
rect 23440 5244 23446 5296
rect 24489 5287 24547 5293
rect 24489 5253 24501 5287
rect 24535 5284 24547 5287
rect 25222 5284 25228 5296
rect 24535 5256 25228 5284
rect 24535 5253 24547 5256
rect 24489 5247 24547 5253
rect 25222 5244 25228 5256
rect 25280 5244 25286 5296
rect 28166 5284 28172 5296
rect 25792 5256 28172 5284
rect 4249 5219 4307 5225
rect 4249 5185 4261 5219
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4614 5216 4620 5228
rect 4387 5188 4620 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 5166 5216 5172 5228
rect 5127 5188 5172 5216
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 4062 5148 4068 5160
rect 4023 5120 4068 5148
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4430 5108 4436 5160
rect 4488 5148 4494 5160
rect 5276 5148 5304 5179
rect 5350 5176 5356 5228
rect 5408 5216 5414 5228
rect 5408 5188 5453 5216
rect 5408 5176 5414 5188
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 6457 5219 6515 5225
rect 5592 5188 5637 5216
rect 5592 5176 5598 5188
rect 6457 5185 6469 5219
rect 6503 5216 6515 5219
rect 6917 5219 6975 5225
rect 6917 5216 6929 5219
rect 6503 5188 6929 5216
rect 6503 5185 6515 5188
rect 6457 5179 6515 5185
rect 6917 5185 6929 5188
rect 6963 5216 6975 5219
rect 7006 5216 7012 5228
rect 6963 5188 7012 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5216 7803 5219
rect 7834 5216 7840 5228
rect 7791 5188 7840 5216
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 7834 5176 7840 5188
rect 7892 5176 7898 5228
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 8662 5216 8668 5228
rect 8435 5188 8668 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 8754 5176 8760 5228
rect 8812 5216 8818 5228
rect 8849 5219 8907 5225
rect 8849 5216 8861 5219
rect 8812 5188 8861 5216
rect 8812 5176 8818 5188
rect 8849 5185 8861 5188
rect 8895 5216 8907 5219
rect 9214 5216 9220 5228
rect 8895 5188 9220 5216
rect 8895 5185 8907 5188
rect 8849 5179 8907 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 9490 5216 9496 5228
rect 9451 5188 9496 5216
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 11790 5176 11796 5228
rect 11848 5216 11854 5228
rect 16117 5219 16175 5225
rect 11848 5188 12558 5216
rect 11848 5176 11854 5188
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16758 5216 16764 5228
rect 16163 5188 16764 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 17954 5176 17960 5228
rect 18012 5216 18018 5228
rect 18233 5219 18291 5225
rect 18233 5216 18245 5219
rect 18012 5188 18245 5216
rect 18012 5176 18018 5188
rect 18233 5185 18245 5188
rect 18279 5185 18291 5219
rect 18233 5179 18291 5185
rect 18785 5219 18843 5225
rect 18785 5185 18797 5219
rect 18831 5185 18843 5219
rect 18785 5179 18843 5185
rect 25133 5219 25191 5225
rect 25133 5185 25145 5219
rect 25179 5216 25191 5219
rect 25314 5216 25320 5228
rect 25179 5188 25320 5216
rect 25179 5185 25191 5188
rect 25133 5179 25191 5185
rect 4488 5120 5304 5148
rect 4488 5108 4494 5120
rect 5552 5080 5580 5176
rect 12342 5148 12348 5160
rect 9048 5120 12348 5148
rect 4448 5052 5580 5080
rect 3237 5015 3295 5021
rect 3237 4981 3249 5015
rect 3283 5012 3295 5015
rect 3418 5012 3424 5024
rect 3283 4984 3424 5012
rect 3283 4981 3295 4984
rect 3237 4975 3295 4981
rect 3418 4972 3424 4984
rect 3476 5012 3482 5024
rect 4448 5012 4476 5052
rect 7190 5040 7196 5092
rect 7248 5080 7254 5092
rect 9048 5089 9076 5120
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 12618 5148 12624 5160
rect 12579 5120 12624 5148
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 16482 5108 16488 5160
rect 16540 5148 16546 5160
rect 18800 5148 18828 5179
rect 25314 5176 25320 5188
rect 25372 5176 25378 5228
rect 25792 5225 25820 5256
rect 28166 5244 28172 5256
rect 28224 5244 28230 5296
rect 25777 5219 25835 5225
rect 25777 5185 25789 5219
rect 25823 5185 25835 5219
rect 26970 5216 26976 5228
rect 26931 5188 26976 5216
rect 25777 5179 25835 5185
rect 26970 5176 26976 5188
rect 27028 5176 27034 5228
rect 27229 5219 27287 5225
rect 27229 5216 27241 5219
rect 27080 5188 27241 5216
rect 16540 5120 18828 5148
rect 16540 5108 16546 5120
rect 22186 5108 22192 5160
rect 22244 5148 22250 5160
rect 22281 5151 22339 5157
rect 22281 5148 22293 5151
rect 22244 5120 22293 5148
rect 22244 5108 22250 5120
rect 22281 5117 22293 5120
rect 22327 5148 22339 5151
rect 24762 5148 24768 5160
rect 22327 5120 24768 5148
rect 22327 5117 22339 5120
rect 22281 5111 22339 5117
rect 24762 5108 24768 5120
rect 24820 5108 24826 5160
rect 25038 5108 25044 5160
rect 25096 5148 25102 5160
rect 27080 5148 27108 5188
rect 27229 5185 27241 5188
rect 27275 5185 27287 5219
rect 27229 5179 27287 5185
rect 30469 5219 30527 5225
rect 30469 5185 30481 5219
rect 30515 5216 30527 5219
rect 31662 5216 31668 5228
rect 30515 5188 31668 5216
rect 30515 5185 30527 5188
rect 30469 5179 30527 5185
rect 31662 5176 31668 5188
rect 31720 5176 31726 5228
rect 32122 5216 32128 5228
rect 32083 5188 32128 5216
rect 32122 5176 32128 5188
rect 32180 5176 32186 5228
rect 32324 5225 32352 5324
rect 33137 5287 33195 5293
rect 33137 5253 33149 5287
rect 33183 5284 33195 5287
rect 33410 5284 33416 5296
rect 33183 5256 33416 5284
rect 33183 5253 33195 5256
rect 33137 5247 33195 5253
rect 33410 5244 33416 5256
rect 33468 5284 33474 5296
rect 35084 5284 35112 5324
rect 35161 5321 35173 5355
rect 35207 5352 35219 5355
rect 39301 5355 39359 5361
rect 39301 5352 39313 5355
rect 35207 5324 39313 5352
rect 35207 5321 35219 5324
rect 35161 5315 35219 5321
rect 39301 5321 39313 5324
rect 39347 5352 39359 5355
rect 41690 5352 41696 5364
rect 39347 5324 39988 5352
rect 41651 5324 41696 5352
rect 39347 5321 39359 5324
rect 39301 5315 39359 5321
rect 33468 5256 35020 5284
rect 35084 5256 39528 5284
rect 33468 5244 33474 5256
rect 32309 5219 32367 5225
rect 32309 5185 32321 5219
rect 32355 5185 32367 5219
rect 32309 5179 32367 5185
rect 32953 5219 33011 5225
rect 32953 5185 32965 5219
rect 32999 5216 33011 5219
rect 33226 5216 33232 5228
rect 32999 5188 33232 5216
rect 32999 5185 33011 5188
rect 32953 5179 33011 5185
rect 33226 5176 33232 5188
rect 33284 5216 33290 5228
rect 33870 5216 33876 5228
rect 33284 5188 33876 5216
rect 33284 5176 33290 5188
rect 33870 5176 33876 5188
rect 33928 5176 33934 5228
rect 34146 5176 34152 5228
rect 34204 5216 34210 5228
rect 34992 5225 35020 5256
rect 34977 5219 35035 5225
rect 34204 5188 34297 5216
rect 34204 5176 34210 5188
rect 34977 5185 34989 5219
rect 35023 5185 35035 5219
rect 34977 5179 35035 5185
rect 35253 5219 35311 5225
rect 35253 5185 35265 5219
rect 35299 5216 35311 5219
rect 35342 5216 35348 5228
rect 35299 5188 35348 5216
rect 35299 5185 35311 5188
rect 35253 5179 35311 5185
rect 35342 5176 35348 5188
rect 35400 5176 35406 5228
rect 36004 5225 36032 5256
rect 39500 5228 39528 5256
rect 35989 5219 36047 5225
rect 35989 5185 36001 5219
rect 36035 5185 36047 5219
rect 36722 5216 36728 5228
rect 36683 5188 36728 5216
rect 35989 5179 36047 5185
rect 36722 5176 36728 5188
rect 36780 5176 36786 5228
rect 37645 5219 37703 5225
rect 37645 5185 37657 5219
rect 37691 5216 37703 5219
rect 38654 5216 38660 5228
rect 37691 5188 38660 5216
rect 37691 5185 37703 5188
rect 37645 5179 37703 5185
rect 38654 5176 38660 5188
rect 38712 5176 38718 5228
rect 38746 5176 38752 5228
rect 38804 5216 38810 5228
rect 39293 5219 39351 5225
rect 39293 5216 39305 5219
rect 38804 5188 39305 5216
rect 38804 5176 38810 5188
rect 39293 5185 39305 5188
rect 39339 5185 39351 5219
rect 39293 5179 39351 5185
rect 39482 5176 39488 5228
rect 39540 5216 39546 5228
rect 39960 5225 39988 5324
rect 41690 5312 41696 5324
rect 41748 5312 41754 5364
rect 42610 5352 42616 5364
rect 42571 5324 42616 5352
rect 42610 5312 42616 5324
rect 42668 5312 42674 5364
rect 44637 5355 44695 5361
rect 44637 5321 44649 5355
rect 44683 5352 44695 5355
rect 50893 5355 50951 5361
rect 44683 5324 45508 5352
rect 44683 5321 44695 5324
rect 44637 5315 44695 5321
rect 42426 5284 42432 5296
rect 40052 5256 42432 5284
rect 39945 5219 40003 5225
rect 39540 5188 39585 5216
rect 39540 5176 39546 5188
rect 39945 5185 39957 5219
rect 39991 5185 40003 5219
rect 39945 5179 40003 5185
rect 25096 5120 27108 5148
rect 25096 5108 25102 5120
rect 29454 5108 29460 5160
rect 29512 5148 29518 5160
rect 30282 5148 30288 5160
rect 29512 5120 30288 5148
rect 29512 5108 29518 5120
rect 30282 5108 30288 5120
rect 30340 5148 30346 5160
rect 30745 5151 30803 5157
rect 30745 5148 30757 5151
rect 30340 5120 30757 5148
rect 30340 5108 30346 5120
rect 30745 5117 30757 5120
rect 30791 5117 30803 5151
rect 30745 5111 30803 5117
rect 32217 5151 32275 5157
rect 32217 5117 32229 5151
rect 32263 5148 32275 5151
rect 32858 5148 32864 5160
rect 32263 5120 32864 5148
rect 32263 5117 32275 5120
rect 32217 5111 32275 5117
rect 32858 5108 32864 5120
rect 32916 5108 32922 5160
rect 33962 5148 33968 5160
rect 33875 5120 33968 5148
rect 33962 5108 33968 5120
rect 34020 5108 34026 5160
rect 8205 5083 8263 5089
rect 8205 5080 8217 5083
rect 7248 5052 8217 5080
rect 7248 5040 7254 5052
rect 8205 5049 8217 5052
rect 8251 5049 8263 5083
rect 8205 5043 8263 5049
rect 9033 5083 9091 5089
rect 9033 5049 9045 5083
rect 9079 5049 9091 5083
rect 9033 5043 9091 5049
rect 11885 5083 11943 5089
rect 11885 5049 11897 5083
rect 11931 5080 11943 5083
rect 12434 5080 12440 5092
rect 11931 5052 12440 5080
rect 11931 5049 11943 5052
rect 11885 5043 11943 5049
rect 12434 5040 12440 5052
rect 12492 5040 12498 5092
rect 15473 5083 15531 5089
rect 15473 5049 15485 5083
rect 15519 5080 15531 5083
rect 16022 5080 16028 5092
rect 15519 5052 16028 5080
rect 15519 5049 15531 5052
rect 15473 5043 15531 5049
rect 16022 5040 16028 5052
rect 16080 5040 16086 5092
rect 17586 5040 17592 5092
rect 17644 5080 17650 5092
rect 18049 5083 18107 5089
rect 18049 5080 18061 5083
rect 17644 5052 18061 5080
rect 17644 5040 17650 5052
rect 18049 5049 18061 5052
rect 18095 5080 18107 5083
rect 18877 5083 18935 5089
rect 18877 5080 18889 5083
rect 18095 5052 18889 5080
rect 18095 5049 18107 5052
rect 18049 5043 18107 5049
rect 18877 5049 18889 5052
rect 18923 5049 18935 5083
rect 18877 5043 18935 5049
rect 19150 5040 19156 5092
rect 19208 5080 19214 5092
rect 24578 5080 24584 5092
rect 19208 5052 24584 5080
rect 19208 5040 19214 5052
rect 24578 5040 24584 5052
rect 24636 5040 24642 5092
rect 29730 5040 29736 5092
rect 29788 5080 29794 5092
rect 32769 5083 32827 5089
rect 32769 5080 32781 5083
rect 29788 5052 32781 5080
rect 29788 5040 29794 5052
rect 32769 5049 32781 5052
rect 32815 5049 32827 5083
rect 32769 5043 32827 5049
rect 3476 4984 4476 5012
rect 3476 4972 3482 4984
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 4893 5015 4951 5021
rect 4893 5012 4905 5015
rect 4764 4984 4905 5012
rect 4764 4972 4770 4984
rect 4893 4981 4905 4984
rect 4939 4981 4951 5015
rect 7098 5012 7104 5024
rect 7059 4984 7104 5012
rect 4893 4975 4951 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 9677 5015 9735 5021
rect 9677 4981 9689 5015
rect 9723 5012 9735 5015
rect 10226 5012 10232 5024
rect 9723 4984 10232 5012
rect 9723 4981 9735 4984
rect 9677 4975 9735 4981
rect 10226 4972 10232 4984
rect 10284 4972 10290 5024
rect 10321 5015 10379 5021
rect 10321 4981 10333 5015
rect 10367 5012 10379 5015
rect 10594 5012 10600 5024
rect 10367 4984 10600 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 10594 4972 10600 4984
rect 10652 4972 10658 5024
rect 10962 5012 10968 5024
rect 10923 4984 10968 5012
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 14185 5015 14243 5021
rect 14185 4981 14197 5015
rect 14231 5012 14243 5015
rect 14458 5012 14464 5024
rect 14231 4984 14464 5012
rect 14231 4981 14243 4984
rect 14185 4975 14243 4981
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 14829 5015 14887 5021
rect 14829 4981 14841 5015
rect 14875 5012 14887 5015
rect 15010 5012 15016 5024
rect 14875 4984 15016 5012
rect 14875 4981 14887 4984
rect 14829 4975 14887 4981
rect 15010 4972 15016 4984
rect 15068 4972 15074 5024
rect 15746 4972 15752 5024
rect 15804 5012 15810 5024
rect 15933 5015 15991 5021
rect 15933 5012 15945 5015
rect 15804 4984 15945 5012
rect 15804 4972 15810 4984
rect 15933 4981 15945 4984
rect 15979 4981 15991 5015
rect 16758 5012 16764 5024
rect 16719 4984 16764 5012
rect 15933 4975 15991 4981
rect 16758 4972 16764 4984
rect 16816 4972 16822 5024
rect 17126 4972 17132 5024
rect 17184 5012 17190 5024
rect 17221 5015 17279 5021
rect 17221 5012 17233 5015
rect 17184 4984 17233 5012
rect 17184 4972 17190 4984
rect 17221 4981 17233 4984
rect 17267 4981 17279 5015
rect 18966 5012 18972 5024
rect 18927 4984 18972 5012
rect 17221 4975 17279 4981
rect 18966 4972 18972 4984
rect 19024 4972 19030 5024
rect 19886 4972 19892 5024
rect 19944 5012 19950 5024
rect 19981 5015 20039 5021
rect 19981 5012 19993 5015
rect 19944 4984 19993 5012
rect 19944 4972 19950 4984
rect 19981 4981 19993 4984
rect 20027 4981 20039 5015
rect 19981 4975 20039 4981
rect 22094 4972 22100 5024
rect 22152 5012 22158 5024
rect 23014 5012 23020 5024
rect 22152 4984 23020 5012
rect 22152 4972 22158 4984
rect 23014 4972 23020 4984
rect 23072 4972 23078 5024
rect 23385 5015 23443 5021
rect 23385 4981 23397 5015
rect 23431 5012 23443 5015
rect 23842 5012 23848 5024
rect 23431 4984 23848 5012
rect 23431 4981 23443 4984
rect 23385 4975 23443 4981
rect 23842 4972 23848 4984
rect 23900 4972 23906 5024
rect 24946 5012 24952 5024
rect 24907 4984 24952 5012
rect 24946 4972 24952 4984
rect 25004 4972 25010 5024
rect 26421 5015 26479 5021
rect 26421 4981 26433 5015
rect 26467 5012 26479 5015
rect 27154 5012 27160 5024
rect 26467 4984 27160 5012
rect 26467 4981 26479 4984
rect 26421 4975 26479 4981
rect 27154 4972 27160 4984
rect 27212 4972 27218 5024
rect 28442 4972 28448 5024
rect 28500 5012 28506 5024
rect 28813 5015 28871 5021
rect 28813 5012 28825 5015
rect 28500 4984 28825 5012
rect 28500 4972 28506 4984
rect 28813 4981 28825 4984
rect 28859 4981 28871 5015
rect 28813 4975 28871 4981
rect 31662 4972 31668 5024
rect 31720 5012 31726 5024
rect 33980 5012 34008 5108
rect 34164 5080 34192 5176
rect 34882 5108 34888 5160
rect 34940 5148 34946 5160
rect 35802 5148 35808 5160
rect 34940 5120 35808 5148
rect 34940 5108 34946 5120
rect 35802 5108 35808 5120
rect 35860 5108 35866 5160
rect 36173 5151 36231 5157
rect 36173 5117 36185 5151
rect 36219 5148 36231 5151
rect 40052 5148 40080 5256
rect 42426 5244 42432 5256
rect 42484 5244 42490 5296
rect 45281 5287 45339 5293
rect 45281 5284 45293 5287
rect 42536 5256 43668 5284
rect 40126 5176 40132 5228
rect 40184 5225 40190 5228
rect 40184 5219 40224 5225
rect 40212 5185 40224 5219
rect 40494 5216 40500 5228
rect 40455 5188 40500 5216
rect 40184 5179 40224 5185
rect 40184 5176 40190 5179
rect 40494 5176 40500 5188
rect 40552 5176 40558 5228
rect 41046 5216 41052 5228
rect 41007 5188 41052 5216
rect 41046 5176 41052 5188
rect 41104 5176 41110 5228
rect 41230 5176 41236 5228
rect 41288 5216 41294 5228
rect 42536 5216 42564 5256
rect 43438 5216 43444 5228
rect 41288 5188 42564 5216
rect 43399 5188 43444 5216
rect 41288 5176 41294 5188
rect 43438 5176 43444 5188
rect 43496 5176 43502 5228
rect 43640 5225 43668 5256
rect 44560 5256 45293 5284
rect 44560 5228 44588 5256
rect 45281 5253 45293 5256
rect 45327 5253 45339 5287
rect 45281 5247 45339 5253
rect 43625 5219 43683 5225
rect 43625 5185 43637 5219
rect 43671 5185 43683 5219
rect 44542 5216 44548 5228
rect 44503 5188 44548 5216
rect 43625 5179 43683 5185
rect 44542 5176 44548 5188
rect 44600 5176 44606 5228
rect 44726 5216 44732 5228
rect 44687 5188 44732 5216
rect 44726 5176 44732 5188
rect 44784 5176 44790 5228
rect 45186 5216 45192 5228
rect 45147 5188 45192 5216
rect 45186 5176 45192 5188
rect 45244 5176 45250 5228
rect 45480 5225 45508 5324
rect 50893 5321 50905 5355
rect 50939 5352 50951 5355
rect 54018 5352 54024 5364
rect 50939 5324 54024 5352
rect 50939 5321 50951 5324
rect 50893 5315 50951 5321
rect 54018 5312 54024 5324
rect 54076 5312 54082 5364
rect 48314 5284 48320 5296
rect 48275 5256 48320 5284
rect 48314 5244 48320 5256
rect 48372 5244 48378 5296
rect 48533 5287 48591 5293
rect 48533 5253 48545 5287
rect 48579 5284 48591 5287
rect 51166 5284 51172 5296
rect 48579 5256 51172 5284
rect 48579 5253 48591 5256
rect 48533 5247 48591 5253
rect 51166 5244 51172 5256
rect 51224 5244 51230 5296
rect 55398 5284 55404 5296
rect 51368 5256 55404 5284
rect 45465 5219 45523 5225
rect 45465 5185 45477 5219
rect 45511 5216 45523 5219
rect 46382 5216 46388 5228
rect 45511 5188 46388 5216
rect 45511 5185 45523 5188
rect 45465 5179 45523 5185
rect 46382 5176 46388 5188
rect 46440 5176 46446 5228
rect 49145 5220 49203 5225
rect 49068 5219 49203 5220
rect 49068 5216 49157 5219
rect 47044 5192 49157 5216
rect 47044 5188 49096 5192
rect 36219 5120 40080 5148
rect 36219 5117 36231 5120
rect 36173 5111 36231 5117
rect 40678 5108 40684 5160
rect 40736 5148 40742 5160
rect 42429 5151 42487 5157
rect 42429 5148 42441 5151
rect 40736 5120 42441 5148
rect 40736 5108 40742 5120
rect 42429 5117 42441 5120
rect 42475 5117 42487 5151
rect 42429 5111 42487 5117
rect 42794 5108 42800 5160
rect 42852 5148 42858 5160
rect 47044 5157 47072 5188
rect 49145 5185 49157 5192
rect 49191 5185 49203 5219
rect 50709 5219 50767 5225
rect 50709 5216 50721 5219
rect 49145 5179 49203 5185
rect 49252 5188 50721 5216
rect 46569 5151 46627 5157
rect 46569 5148 46581 5151
rect 42852 5120 42897 5148
rect 45296 5120 46581 5148
rect 42852 5108 42858 5120
rect 34164 5052 38332 5080
rect 34330 5012 34336 5024
rect 31720 4984 34008 5012
rect 34291 4984 34336 5012
rect 31720 4972 31726 4984
rect 34330 4972 34336 4984
rect 34388 4972 34394 5024
rect 34793 5015 34851 5021
rect 34793 4981 34805 5015
rect 34839 5012 34851 5015
rect 35434 5012 35440 5024
rect 34839 4984 35440 5012
rect 34839 4981 34851 4984
rect 34793 4975 34851 4981
rect 35434 4972 35440 4984
rect 35492 4972 35498 5024
rect 37550 5012 37556 5024
rect 37511 4984 37556 5012
rect 37550 4972 37556 4984
rect 37608 4972 37614 5024
rect 38194 5012 38200 5024
rect 38155 4984 38200 5012
rect 38194 4972 38200 4984
rect 38252 4972 38258 5024
rect 38304 5012 38332 5052
rect 40218 5040 40224 5092
rect 40276 5080 40282 5092
rect 44542 5080 44548 5092
rect 40276 5052 40321 5080
rect 42812 5052 44548 5080
rect 40276 5040 40282 5052
rect 39206 5012 39212 5024
rect 38304 4984 39212 5012
rect 39206 4972 39212 4984
rect 39264 4972 39270 5024
rect 39758 4972 39764 5024
rect 39816 5012 39822 5024
rect 41233 5015 41291 5021
rect 41233 5012 41245 5015
rect 39816 4984 41245 5012
rect 39816 4972 39822 4984
rect 41233 4981 41245 4984
rect 41279 4981 41291 5015
rect 41233 4975 41291 4981
rect 42426 4972 42432 5024
rect 42484 5012 42490 5024
rect 42812 5021 42840 5052
rect 44542 5040 44548 5052
rect 44600 5040 44606 5092
rect 42797 5015 42855 5021
rect 42797 5012 42809 5015
rect 42484 4984 42809 5012
rect 42484 4972 42490 4984
rect 42797 4981 42809 4984
rect 42843 4981 42855 5015
rect 43438 5012 43444 5024
rect 43399 4984 43444 5012
rect 42797 4975 42855 4981
rect 43438 4972 43444 4984
rect 43496 4972 43502 5024
rect 44634 4972 44640 5024
rect 44692 5012 44698 5024
rect 45296 5012 45324 5120
rect 46569 5117 46581 5120
rect 46615 5117 46627 5151
rect 46569 5111 46627 5117
rect 47029 5151 47087 5157
rect 47029 5117 47041 5151
rect 47075 5117 47087 5151
rect 49252 5148 49280 5188
rect 50709 5185 50721 5188
rect 50755 5185 50767 5219
rect 50890 5216 50896 5228
rect 50851 5188 50896 5216
rect 50709 5179 50767 5185
rect 50890 5176 50896 5188
rect 50948 5176 50954 5228
rect 51368 5225 51396 5256
rect 55398 5244 55404 5256
rect 55456 5244 55462 5296
rect 51353 5219 51411 5225
rect 51353 5185 51365 5219
rect 51399 5185 51411 5219
rect 51994 5216 52000 5228
rect 51907 5188 52000 5216
rect 51353 5179 51411 5185
rect 51994 5176 52000 5188
rect 52052 5216 52058 5228
rect 52733 5219 52791 5225
rect 52733 5216 52745 5219
rect 52052 5188 52745 5216
rect 52052 5176 52058 5188
rect 52733 5185 52745 5188
rect 52779 5185 52791 5219
rect 52733 5179 52791 5185
rect 53561 5219 53619 5225
rect 53561 5185 53573 5219
rect 53607 5185 53619 5219
rect 53561 5179 53619 5185
rect 55125 5219 55183 5225
rect 55125 5185 55137 5219
rect 55171 5216 55183 5219
rect 55674 5216 55680 5228
rect 55171 5188 55680 5216
rect 55171 5185 55183 5188
rect 55125 5179 55183 5185
rect 47029 5111 47087 5117
rect 48516 5120 49280 5148
rect 45370 5040 45376 5092
rect 45428 5080 45434 5092
rect 46845 5083 46903 5089
rect 46845 5080 46857 5083
rect 45428 5052 46857 5080
rect 45428 5040 45434 5052
rect 46845 5049 46857 5052
rect 46891 5049 46903 5083
rect 46845 5043 46903 5049
rect 47118 5040 47124 5092
rect 47176 5080 47182 5092
rect 48516 5080 48544 5120
rect 49326 5108 49332 5160
rect 49384 5148 49390 5160
rect 49789 5151 49847 5157
rect 49789 5148 49801 5151
rect 49384 5120 49801 5148
rect 49384 5108 49390 5120
rect 49789 5117 49801 5120
rect 49835 5117 49847 5151
rect 49789 5111 49847 5117
rect 51258 5108 51264 5160
rect 51316 5148 51322 5160
rect 52012 5148 52040 5176
rect 51316 5120 52040 5148
rect 53576 5148 53604 5179
rect 55674 5176 55680 5188
rect 55732 5176 55738 5228
rect 55582 5148 55588 5160
rect 53576 5120 55588 5148
rect 51316 5108 51322 5120
rect 55582 5108 55588 5120
rect 55640 5108 55646 5160
rect 47176 5052 48544 5080
rect 47176 5040 47182 5052
rect 44692 4984 45324 5012
rect 45649 5015 45707 5021
rect 44692 4972 44698 4984
rect 45649 4981 45661 5015
rect 45695 5012 45707 5015
rect 46290 5012 46296 5024
rect 45695 4984 46296 5012
rect 45695 4981 45707 4984
rect 45649 4975 45707 4981
rect 46290 4972 46296 4984
rect 46348 4972 46354 5024
rect 46750 4972 46756 5024
rect 46808 5012 46814 5024
rect 48516 5021 48544 5052
rect 48685 5083 48743 5089
rect 48685 5049 48697 5083
rect 48731 5080 48743 5083
rect 50154 5080 50160 5092
rect 48731 5052 50160 5080
rect 48731 5049 48743 5052
rect 48685 5043 48743 5049
rect 50154 5040 50160 5052
rect 50212 5040 50218 5092
rect 51537 5083 51595 5089
rect 51537 5049 51549 5083
rect 51583 5080 51595 5083
rect 52546 5080 52552 5092
rect 51583 5052 52552 5080
rect 51583 5049 51595 5052
rect 51537 5043 51595 5049
rect 52546 5040 52552 5052
rect 52604 5040 52610 5092
rect 52730 5040 52736 5092
rect 52788 5080 52794 5092
rect 54021 5083 54079 5089
rect 54021 5080 54033 5083
rect 52788 5052 54033 5080
rect 52788 5040 52794 5052
rect 54021 5049 54033 5052
rect 54067 5049 54079 5083
rect 54021 5043 54079 5049
rect 47581 5015 47639 5021
rect 47581 5012 47593 5015
rect 46808 4984 47593 5012
rect 46808 4972 46814 4984
rect 47581 4981 47593 4984
rect 47627 4981 47639 5015
rect 47581 4975 47639 4981
rect 48501 5015 48559 5021
rect 48501 4981 48513 5015
rect 48547 4981 48559 5015
rect 48501 4975 48559 4981
rect 49329 5015 49387 5021
rect 49329 4981 49341 5015
rect 49375 5012 49387 5015
rect 49602 5012 49608 5024
rect 49375 4984 49608 5012
rect 49375 4981 49387 4984
rect 49329 4975 49387 4981
rect 49602 4972 49608 4984
rect 49660 4972 49666 5024
rect 52089 5015 52147 5021
rect 52089 4981 52101 5015
rect 52135 5012 52147 5015
rect 52638 5012 52644 5024
rect 52135 4984 52644 5012
rect 52135 4981 52147 4984
rect 52089 4975 52147 4981
rect 52638 4972 52644 4984
rect 52696 4972 52702 5024
rect 52822 5012 52828 5024
rect 52783 4984 52828 5012
rect 52822 4972 52828 4984
rect 52880 4972 52886 5024
rect 53006 4972 53012 5024
rect 53064 5012 53070 5024
rect 53377 5015 53435 5021
rect 53377 5012 53389 5015
rect 53064 4984 53389 5012
rect 53064 4972 53070 4984
rect 53377 4981 53389 4984
rect 53423 4981 53435 5015
rect 55306 5012 55312 5024
rect 55267 4984 55312 5012
rect 53377 4975 53435 4981
rect 55306 4972 55312 4984
rect 55364 4972 55370 5024
rect 55766 5012 55772 5024
rect 55727 4984 55772 5012
rect 55766 4972 55772 4984
rect 55824 5012 55830 5024
rect 56321 5015 56379 5021
rect 56321 5012 56333 5015
rect 55824 4984 56333 5012
rect 55824 4972 55830 4984
rect 56321 4981 56333 4984
rect 56367 4981 56379 5015
rect 56321 4975 56379 4981
rect 1104 4922 58880 4944
rect 1104 4870 8174 4922
rect 8226 4870 8238 4922
rect 8290 4870 8302 4922
rect 8354 4870 8366 4922
rect 8418 4870 8430 4922
rect 8482 4870 22622 4922
rect 22674 4870 22686 4922
rect 22738 4870 22750 4922
rect 22802 4870 22814 4922
rect 22866 4870 22878 4922
rect 22930 4870 37070 4922
rect 37122 4870 37134 4922
rect 37186 4870 37198 4922
rect 37250 4870 37262 4922
rect 37314 4870 37326 4922
rect 37378 4870 51518 4922
rect 51570 4870 51582 4922
rect 51634 4870 51646 4922
rect 51698 4870 51710 4922
rect 51762 4870 51774 4922
rect 51826 4870 58880 4922
rect 1104 4848 58880 4870
rect 3237 4811 3295 4817
rect 3237 4777 3249 4811
rect 3283 4808 3295 4811
rect 4246 4808 4252 4820
rect 3283 4780 4252 4808
rect 3283 4777 3295 4780
rect 3237 4771 3295 4777
rect 4246 4768 4252 4780
rect 4304 4768 4310 4820
rect 4614 4808 4620 4820
rect 4448 4780 4620 4808
rect 3145 4743 3203 4749
rect 3145 4709 3157 4743
rect 3191 4740 3203 4743
rect 4448 4740 4476 4780
rect 4614 4768 4620 4780
rect 4672 4808 4678 4820
rect 6549 4811 6607 4817
rect 4672 4780 6500 4808
rect 4672 4768 4678 4780
rect 3191 4712 4476 4740
rect 3191 4709 3203 4712
rect 3145 4703 3203 4709
rect 6472 4681 6500 4780
rect 6549 4777 6561 4811
rect 6595 4808 6607 4811
rect 11698 4808 11704 4820
rect 6595 4780 11704 4808
rect 6595 4777 6607 4780
rect 6549 4771 6607 4777
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 12713 4811 12771 4817
rect 12713 4777 12725 4811
rect 12759 4808 12771 4811
rect 13078 4808 13084 4820
rect 12759 4780 13084 4808
rect 12759 4777 12771 4780
rect 12713 4771 12771 4777
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 18138 4808 18144 4820
rect 18099 4780 18144 4808
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 18966 4768 18972 4820
rect 19024 4808 19030 4820
rect 23845 4811 23903 4817
rect 19024 4780 22508 4808
rect 19024 4768 19030 4780
rect 9309 4743 9367 4749
rect 9309 4709 9321 4743
rect 9355 4740 9367 4743
rect 10318 4740 10324 4752
rect 9355 4712 10324 4740
rect 9355 4709 9367 4712
rect 9309 4703 9367 4709
rect 10318 4700 10324 4712
rect 10376 4700 10382 4752
rect 11790 4740 11796 4752
rect 11751 4712 11796 4740
rect 11790 4700 11796 4712
rect 11848 4700 11854 4752
rect 12986 4700 12992 4752
rect 13044 4740 13050 4752
rect 16114 4740 16120 4752
rect 13044 4712 16120 4740
rect 13044 4700 13050 4712
rect 16114 4700 16120 4712
rect 16172 4700 16178 4752
rect 18046 4740 18052 4752
rect 17696 4712 18052 4740
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4672 6515 4675
rect 8294 4672 8300 4684
rect 6503 4644 8300 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 9398 4672 9404 4684
rect 8435 4644 9404 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 9398 4632 9404 4644
rect 9456 4632 9462 4684
rect 9858 4632 9864 4684
rect 9916 4672 9922 4684
rect 10413 4675 10471 4681
rect 10413 4672 10425 4675
rect 9916 4644 10425 4672
rect 9916 4632 9922 4644
rect 10413 4641 10425 4644
rect 10459 4641 10471 4675
rect 10413 4635 10471 4641
rect 12621 4675 12679 4681
rect 12621 4641 12633 4675
rect 12667 4672 12679 4675
rect 13170 4672 13176 4684
rect 12667 4644 13176 4672
rect 12667 4641 12679 4644
rect 12621 4635 12679 4641
rect 13170 4632 13176 4644
rect 13228 4632 13234 4684
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 16666 4672 16672 4684
rect 15335 4644 16672 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 16945 4675 17003 4681
rect 16945 4641 16957 4675
rect 16991 4672 17003 4675
rect 17402 4672 17408 4684
rect 16991 4644 17408 4672
rect 16991 4641 17003 4644
rect 16945 4635 17003 4641
rect 17402 4632 17408 4644
rect 17460 4632 17466 4684
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 3786 4604 3792 4616
rect 3292 4576 3337 4604
rect 3747 4576 3792 4604
rect 3292 4564 3298 4576
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 4154 4564 4160 4616
rect 4212 4604 4218 4616
rect 4706 4613 4712 4616
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4212 4576 4445 4604
rect 4212 4564 4218 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4700 4604 4712 4613
rect 4667 4576 4712 4604
rect 4433 4567 4491 4573
rect 4700 4567 4712 4576
rect 4706 4564 4712 4567
rect 4764 4564 4770 4616
rect 5810 4564 5816 4616
rect 5868 4604 5874 4616
rect 6546 4604 6552 4616
rect 5868 4576 6552 4604
rect 5868 4564 5874 4576
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7561 4607 7619 4613
rect 7561 4604 7573 4607
rect 7156 4576 7573 4604
rect 7156 4564 7162 4576
rect 7561 4573 7573 4576
rect 7607 4573 7619 4607
rect 7742 4604 7748 4616
rect 7703 4576 7748 4604
rect 7561 4567 7619 4573
rect 7742 4564 7748 4576
rect 7800 4564 7806 4616
rect 9950 4604 9956 4616
rect 9911 4576 9956 4604
rect 9950 4564 9956 4576
rect 10008 4564 10014 4616
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 12437 4607 12495 4613
rect 10284 4576 12388 4604
rect 10284 4564 10290 4576
rect 2961 4539 3019 4545
rect 2961 4505 2973 4539
rect 3007 4536 3019 4539
rect 4062 4536 4068 4548
rect 3007 4508 4068 4536
rect 3007 4505 3019 4508
rect 2961 4499 3019 4505
rect 4062 4496 4068 4508
rect 4120 4496 4126 4548
rect 6270 4536 6276 4548
rect 6231 4508 6276 4536
rect 6270 4496 6276 4508
rect 6328 4496 6334 4548
rect 9674 4536 9680 4548
rect 6932 4508 9680 4536
rect 3973 4471 4031 4477
rect 3973 4437 3985 4471
rect 4019 4468 4031 4471
rect 4246 4468 4252 4480
rect 4019 4440 4252 4468
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 5813 4471 5871 4477
rect 5813 4468 5825 4471
rect 5224 4440 5825 4468
rect 5224 4428 5230 4440
rect 5813 4437 5825 4440
rect 5859 4468 5871 4471
rect 6932 4468 6960 4508
rect 9674 4496 9680 4508
rect 9732 4496 9738 4548
rect 10680 4539 10738 4545
rect 10680 4505 10692 4539
rect 10726 4536 10738 4539
rect 11514 4536 11520 4548
rect 10726 4508 11520 4536
rect 10726 4505 10738 4508
rect 10680 4499 10738 4505
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 5859 4440 6960 4468
rect 7101 4471 7159 4477
rect 5859 4437 5871 4440
rect 5813 4431 5871 4437
rect 7101 4437 7113 4471
rect 7147 4468 7159 4471
rect 7282 4468 7288 4480
rect 7147 4440 7288 4468
rect 7147 4437 7159 4440
rect 7101 4431 7159 4437
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 7650 4468 7656 4480
rect 7611 4440 7656 4468
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 9582 4428 9588 4480
rect 9640 4468 9646 4480
rect 9769 4471 9827 4477
rect 9769 4468 9781 4471
rect 9640 4440 9781 4468
rect 9640 4428 9646 4440
rect 9769 4437 9781 4440
rect 9815 4437 9827 4471
rect 9769 4431 9827 4437
rect 11974 4428 11980 4480
rect 12032 4468 12038 4480
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 12032 4440 12265 4468
rect 12032 4428 12038 4440
rect 12253 4437 12265 4440
rect 12299 4437 12311 4471
rect 12360 4468 12388 4576
rect 12437 4573 12449 4607
rect 12483 4573 12495 4607
rect 12710 4604 12716 4616
rect 12671 4576 12716 4604
rect 12437 4567 12495 4573
rect 12452 4536 12480 4567
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4604 13599 4607
rect 14182 4604 14188 4616
rect 13587 4576 14188 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14366 4564 14372 4616
rect 14424 4604 14430 4616
rect 14461 4607 14519 4613
rect 14461 4604 14473 4607
rect 14424 4576 14473 4604
rect 14424 4564 14430 4576
rect 14461 4573 14473 4576
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 12618 4536 12624 4548
rect 12452 4508 12624 4536
rect 12618 4496 12624 4508
rect 12676 4496 12682 4548
rect 14476 4536 14504 4567
rect 15378 4564 15384 4616
rect 15436 4604 15442 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15436 4576 15761 4604
rect 15436 4564 15442 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 17586 4604 17592 4616
rect 17547 4576 17592 4604
rect 15749 4567 15807 4573
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 17696 4613 17724 4712
rect 18046 4700 18052 4712
rect 18104 4700 18110 4752
rect 18601 4743 18659 4749
rect 18601 4709 18613 4743
rect 18647 4740 18659 4743
rect 20625 4743 20683 4749
rect 18647 4712 19104 4740
rect 18647 4709 18659 4712
rect 18601 4703 18659 4709
rect 18322 4672 18328 4684
rect 17788 4644 18328 4672
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4573 17739 4607
rect 17681 4567 17739 4573
rect 15838 4536 15844 4548
rect 14476 4508 15844 4536
rect 15838 4496 15844 4508
rect 15896 4496 15902 4548
rect 16114 4496 16120 4548
rect 16172 4536 16178 4548
rect 17405 4539 17463 4545
rect 17405 4536 17417 4539
rect 16172 4508 17417 4536
rect 16172 4496 16178 4508
rect 17405 4505 17417 4508
rect 17451 4536 17463 4539
rect 17788 4536 17816 4644
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 18414 4604 18420 4616
rect 18375 4576 18420 4604
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 19076 4604 19104 4712
rect 20625 4709 20637 4743
rect 20671 4740 20683 4743
rect 22094 4740 22100 4752
rect 20671 4712 22100 4740
rect 20671 4709 20683 4712
rect 20625 4703 20683 4709
rect 22094 4700 22100 4712
rect 22152 4740 22158 4752
rect 22152 4712 22416 4740
rect 22152 4700 22158 4712
rect 19242 4672 19248 4684
rect 19203 4644 19248 4672
rect 19242 4632 19248 4644
rect 19300 4632 19306 4684
rect 21192 4644 22324 4672
rect 21192 4604 21220 4644
rect 19076 4576 21220 4604
rect 21266 4564 21272 4616
rect 21324 4604 21330 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 21324 4576 21373 4604
rect 21324 4564 21330 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 17451 4508 17816 4536
rect 17451 4505 17463 4508
rect 17405 4499 17463 4505
rect 17954 4496 17960 4548
rect 18012 4536 18018 4548
rect 18141 4539 18199 4545
rect 18141 4536 18153 4539
rect 18012 4508 18153 4536
rect 18012 4496 18018 4508
rect 18141 4505 18153 4508
rect 18187 4505 18199 4539
rect 18141 4499 18199 4505
rect 19512 4539 19570 4545
rect 19512 4505 19524 4539
rect 19558 4536 19570 4539
rect 22097 4539 22155 4545
rect 22097 4536 22109 4539
rect 19558 4508 22109 4536
rect 19558 4505 19570 4508
rect 19512 4499 19570 4505
rect 22097 4505 22109 4508
rect 22143 4505 22155 4539
rect 22296 4536 22324 4644
rect 22388 4613 22416 4712
rect 22480 4613 22508 4780
rect 23216 4780 23704 4808
rect 22373 4607 22431 4613
rect 22373 4573 22385 4607
rect 22419 4573 22431 4607
rect 22373 4567 22431 4573
rect 22465 4607 22523 4613
rect 22465 4573 22477 4607
rect 22511 4573 22523 4607
rect 22465 4567 22523 4573
rect 22554 4564 22560 4616
rect 22612 4604 22618 4616
rect 22612 4576 22657 4604
rect 22612 4564 22618 4576
rect 22738 4564 22744 4616
rect 22796 4604 22802 4616
rect 23216 4613 23244 4780
rect 23382 4700 23388 4752
rect 23440 4700 23446 4752
rect 23400 4672 23428 4700
rect 23676 4672 23704 4780
rect 23845 4777 23857 4811
rect 23891 4808 23903 4811
rect 30101 4811 30159 4817
rect 23891 4780 27568 4808
rect 23891 4777 23903 4780
rect 23845 4771 23903 4777
rect 25038 4740 25044 4752
rect 24999 4712 25044 4740
rect 25038 4700 25044 4712
rect 25096 4700 25102 4752
rect 23400 4644 23520 4672
rect 23676 4644 24440 4672
rect 23492 4613 23520 4644
rect 23201 4607 23259 4613
rect 23201 4604 23213 4607
rect 22796 4576 23213 4604
rect 22796 4564 22802 4576
rect 23201 4573 23213 4576
rect 23247 4573 23259 4607
rect 23201 4567 23259 4573
rect 23385 4607 23443 4613
rect 23385 4573 23397 4607
rect 23431 4573 23443 4607
rect 23385 4567 23443 4573
rect 23477 4607 23535 4613
rect 23477 4573 23489 4607
rect 23523 4573 23535 4607
rect 23477 4567 23535 4573
rect 23569 4607 23627 4613
rect 23569 4573 23581 4607
rect 23615 4604 23627 4607
rect 24210 4604 24216 4616
rect 23615 4576 24216 4604
rect 23615 4573 23627 4576
rect 23569 4567 23627 4573
rect 23400 4536 23428 4567
rect 24210 4564 24216 4576
rect 24268 4564 24274 4616
rect 24412 4613 24440 4644
rect 25130 4632 25136 4684
rect 25188 4672 25194 4684
rect 25869 4675 25927 4681
rect 25869 4672 25881 4675
rect 25188 4644 25881 4672
rect 25188 4632 25194 4644
rect 25869 4641 25881 4644
rect 25915 4641 25927 4675
rect 25869 4635 25927 4641
rect 26145 4675 26203 4681
rect 26145 4641 26157 4675
rect 26191 4672 26203 4675
rect 26878 4672 26884 4684
rect 26191 4644 26884 4672
rect 26191 4641 26203 4644
rect 26145 4635 26203 4641
rect 26878 4632 26884 4644
rect 26936 4632 26942 4684
rect 27540 4672 27568 4780
rect 30101 4777 30113 4811
rect 30147 4808 30159 4811
rect 30282 4808 30288 4820
rect 30147 4780 30288 4808
rect 30147 4777 30159 4780
rect 30101 4771 30159 4777
rect 30282 4768 30288 4780
rect 30340 4768 30346 4820
rect 33137 4811 33195 4817
rect 33137 4808 33149 4811
rect 30668 4780 33149 4808
rect 27617 4743 27675 4749
rect 27617 4709 27629 4743
rect 27663 4740 27675 4743
rect 29454 4740 29460 4752
rect 27663 4712 29460 4740
rect 27663 4709 27675 4712
rect 27617 4703 27675 4709
rect 29454 4700 29460 4712
rect 29512 4700 29518 4752
rect 30668 4740 30696 4780
rect 33137 4777 33149 4780
rect 33183 4777 33195 4811
rect 35618 4808 35624 4820
rect 33137 4771 33195 4777
rect 35176 4780 35624 4808
rect 29564 4712 30696 4740
rect 29564 4684 29592 4712
rect 32122 4700 32128 4752
rect 32180 4740 32186 4752
rect 32585 4743 32643 4749
rect 32585 4740 32597 4743
rect 32180 4712 32597 4740
rect 32180 4700 32186 4712
rect 32585 4709 32597 4712
rect 32631 4709 32643 4743
rect 32585 4703 32643 4709
rect 29546 4672 29552 4684
rect 27540 4644 28396 4672
rect 29507 4644 29552 4672
rect 24397 4607 24455 4613
rect 24397 4573 24409 4607
rect 24443 4573 24455 4607
rect 24578 4604 24584 4616
rect 24539 4576 24584 4604
rect 24397 4567 24455 4573
rect 24578 4564 24584 4576
rect 24636 4564 24642 4616
rect 24673 4607 24731 4613
rect 24673 4573 24685 4607
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4604 24823 4607
rect 25774 4604 25780 4616
rect 24811 4576 25780 4604
rect 24811 4573 24823 4576
rect 24765 4567 24823 4573
rect 22296 4508 23428 4536
rect 22097 4499 22155 4505
rect 12710 4468 12716 4480
rect 12360 4440 12716 4468
rect 12253 4431 12311 4437
rect 12710 4428 12716 4440
rect 12768 4428 12774 4480
rect 14645 4471 14703 4477
rect 14645 4437 14657 4471
rect 14691 4468 14703 4471
rect 15194 4468 15200 4480
rect 14691 4440 15200 4468
rect 14691 4437 14703 4440
rect 14645 4431 14703 4437
rect 15194 4428 15200 4440
rect 15252 4428 15258 4480
rect 15930 4468 15936 4480
rect 15891 4440 15936 4468
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 17681 4471 17739 4477
rect 17681 4437 17693 4471
rect 17727 4468 17739 4471
rect 24688 4468 24716 4567
rect 25774 4564 25780 4576
rect 25832 4564 25838 4616
rect 28258 4604 28264 4616
rect 28219 4576 28264 4604
rect 28258 4564 28264 4576
rect 28316 4564 28322 4616
rect 28169 4539 28227 4545
rect 28169 4536 28181 4539
rect 27370 4508 28181 4536
rect 28169 4505 28181 4508
rect 28215 4505 28227 4539
rect 28368 4536 28396 4644
rect 29546 4632 29552 4644
rect 29604 4632 29610 4684
rect 35176 4681 35204 4780
rect 35618 4768 35624 4780
rect 35676 4768 35682 4820
rect 35802 4768 35808 4820
rect 35860 4808 35866 4820
rect 36909 4811 36967 4817
rect 36909 4808 36921 4811
rect 35860 4780 36921 4808
rect 35860 4768 35866 4780
rect 36909 4777 36921 4780
rect 36955 4808 36967 4811
rect 38746 4808 38752 4820
rect 36955 4780 38752 4808
rect 36955 4777 36967 4780
rect 36909 4771 36967 4777
rect 38746 4768 38752 4780
rect 38804 4768 38810 4820
rect 39482 4768 39488 4820
rect 39540 4808 39546 4820
rect 41049 4811 41107 4817
rect 41049 4808 41061 4811
rect 39540 4780 41061 4808
rect 39540 4768 39546 4780
rect 41049 4777 41061 4780
rect 41095 4808 41107 4811
rect 41230 4808 41236 4820
rect 41095 4780 41236 4808
rect 41095 4777 41107 4780
rect 41049 4771 41107 4777
rect 41230 4768 41236 4780
rect 41288 4768 41294 4820
rect 42426 4808 42432 4820
rect 41386 4780 42432 4808
rect 37829 4743 37887 4749
rect 37829 4709 37841 4743
rect 37875 4740 37887 4743
rect 38654 4740 38660 4752
rect 37875 4712 38660 4740
rect 37875 4709 37887 4712
rect 37829 4703 37887 4709
rect 38654 4700 38660 4712
rect 38712 4740 38718 4752
rect 39114 4740 39120 4752
rect 38712 4712 39120 4740
rect 38712 4700 38718 4712
rect 39114 4700 39120 4712
rect 39172 4700 39178 4752
rect 39206 4700 39212 4752
rect 39264 4740 39270 4752
rect 41386 4740 41414 4780
rect 42426 4768 42432 4780
rect 42484 4768 42490 4820
rect 42539 4811 42597 4817
rect 42539 4777 42551 4811
rect 42585 4808 42597 4811
rect 43438 4808 43444 4820
rect 42585 4780 43444 4808
rect 42585 4777 42597 4780
rect 42539 4771 42597 4777
rect 43438 4768 43444 4780
rect 43496 4768 43502 4820
rect 44358 4768 44364 4820
rect 44416 4808 44422 4820
rect 48314 4808 48320 4820
rect 44416 4780 48320 4808
rect 44416 4768 44422 4780
rect 48314 4768 48320 4780
rect 48372 4768 48378 4820
rect 51166 4808 51172 4820
rect 51127 4780 51172 4808
rect 51166 4768 51172 4780
rect 51224 4768 51230 4820
rect 52454 4768 52460 4820
rect 52512 4808 52518 4820
rect 55674 4808 55680 4820
rect 52512 4780 53144 4808
rect 55635 4780 55680 4808
rect 52512 4768 52518 4780
rect 39264 4712 41414 4740
rect 39264 4700 39270 4712
rect 42886 4700 42892 4752
rect 42944 4740 42950 4752
rect 44269 4743 44327 4749
rect 44269 4740 44281 4743
rect 42944 4712 44281 4740
rect 42944 4700 42950 4712
rect 44269 4709 44281 4712
rect 44315 4709 44327 4743
rect 48590 4740 48596 4752
rect 48551 4712 48596 4740
rect 44269 4703 44327 4709
rect 48590 4700 48596 4712
rect 48648 4700 48654 4752
rect 49602 4700 49608 4752
rect 49660 4740 49666 4752
rect 49660 4712 51074 4740
rect 49660 4700 49666 4712
rect 35161 4675 35219 4681
rect 35161 4641 35173 4675
rect 35207 4641 35219 4675
rect 35434 4672 35440 4684
rect 35395 4644 35440 4672
rect 35161 4635 35219 4641
rect 35434 4632 35440 4644
rect 35492 4632 35498 4684
rect 38746 4632 38752 4684
rect 38804 4672 38810 4684
rect 41046 4672 41052 4684
rect 38804 4644 41052 4672
rect 38804 4632 38810 4644
rect 41046 4632 41052 4644
rect 41104 4632 41110 4684
rect 41782 4632 41788 4684
rect 41840 4672 41846 4684
rect 42797 4675 42855 4681
rect 42797 4672 42809 4675
rect 41840 4644 42809 4672
rect 41840 4632 41846 4644
rect 42797 4641 42809 4644
rect 42843 4672 42855 4675
rect 46014 4672 46020 4684
rect 42843 4644 46020 4672
rect 42843 4641 42855 4644
rect 42797 4635 42855 4641
rect 46014 4632 46020 4644
rect 46072 4632 46078 4684
rect 46290 4672 46296 4684
rect 46251 4644 46296 4672
rect 46290 4632 46296 4644
rect 46348 4632 46354 4684
rect 46382 4632 46388 4684
rect 46440 4672 46446 4684
rect 46440 4644 48314 4672
rect 46440 4632 46446 4644
rect 28718 4564 28724 4616
rect 28776 4604 28782 4616
rect 28813 4607 28871 4613
rect 28813 4604 28825 4607
rect 28776 4576 28825 4604
rect 28776 4564 28782 4576
rect 28813 4573 28825 4576
rect 28859 4573 28871 4607
rect 28813 4567 28871 4573
rect 29917 4607 29975 4613
rect 29917 4573 29929 4607
rect 29963 4604 29975 4607
rect 30650 4604 30656 4616
rect 29963 4576 30656 4604
rect 29963 4573 29975 4576
rect 29917 4567 29975 4573
rect 30650 4564 30656 4576
rect 30708 4564 30714 4616
rect 30745 4607 30803 4613
rect 30745 4573 30757 4607
rect 30791 4604 30803 4607
rect 31386 4604 31392 4616
rect 30791 4576 31392 4604
rect 30791 4573 30803 4576
rect 30745 4567 30803 4573
rect 31386 4564 31392 4576
rect 31444 4564 31450 4616
rect 33870 4604 33876 4616
rect 33831 4576 33876 4604
rect 33870 4564 33876 4576
rect 33928 4564 33934 4616
rect 34149 4607 34207 4613
rect 34149 4573 34161 4607
rect 34195 4604 34207 4607
rect 35066 4604 35072 4616
rect 34195 4576 35072 4604
rect 34195 4573 34207 4576
rect 34149 4567 34207 4573
rect 35066 4564 35072 4576
rect 35124 4604 35130 4616
rect 37550 4604 37556 4616
rect 35124 4576 35204 4604
rect 36570 4576 37556 4604
rect 35124 4564 35130 4576
rect 30990 4539 31048 4545
rect 30990 4536 31002 4539
rect 28368 4508 31002 4536
rect 28169 4499 28227 4505
rect 30990 4505 31002 4508
rect 31036 4505 31048 4539
rect 34422 4536 34428 4548
rect 30990 4499 31048 4505
rect 31726 4508 34428 4536
rect 17727 4440 24716 4468
rect 17727 4437 17739 4440
rect 17681 4431 17739 4437
rect 26142 4428 26148 4480
rect 26200 4468 26206 4480
rect 29733 4471 29791 4477
rect 29733 4468 29745 4471
rect 26200 4440 29745 4468
rect 26200 4428 26206 4440
rect 29733 4437 29745 4440
rect 29779 4468 29791 4471
rect 31726 4468 31754 4508
rect 34422 4496 34428 4508
rect 34480 4496 34486 4548
rect 35176 4536 35204 4576
rect 37550 4564 37556 4576
rect 37608 4564 37614 4616
rect 37642 4564 37648 4616
rect 37700 4604 37706 4616
rect 38378 4604 38384 4616
rect 37700 4576 38384 4604
rect 37700 4564 37706 4576
rect 38378 4564 38384 4576
rect 38436 4564 38442 4616
rect 40037 4607 40095 4613
rect 40037 4573 40049 4607
rect 40083 4604 40095 4607
rect 40083 4576 40632 4604
rect 40083 4573 40095 4576
rect 40037 4567 40095 4573
rect 35710 4536 35716 4548
rect 35176 4508 35716 4536
rect 35710 4496 35716 4508
rect 35768 4496 35774 4548
rect 39945 4539 40003 4545
rect 39945 4536 39957 4539
rect 36832 4508 39957 4536
rect 29779 4440 31754 4468
rect 32125 4471 32183 4477
rect 29779 4437 29791 4440
rect 29733 4431 29791 4437
rect 32125 4437 32137 4471
rect 32171 4468 32183 4471
rect 32582 4468 32588 4480
rect 32171 4440 32588 4468
rect 32171 4437 32183 4440
rect 32125 4431 32183 4437
rect 32582 4428 32588 4440
rect 32640 4428 32646 4480
rect 35802 4428 35808 4480
rect 35860 4468 35866 4480
rect 36832 4468 36860 4508
rect 39945 4505 39957 4508
rect 39991 4505 40003 4539
rect 39945 4499 40003 4505
rect 40604 4480 40632 4576
rect 43346 4564 43352 4616
rect 43404 4604 43410 4616
rect 43441 4607 43499 4613
rect 43441 4604 43453 4607
rect 43404 4576 43453 4604
rect 43404 4564 43410 4576
rect 43441 4573 43453 4576
rect 43487 4573 43499 4607
rect 43441 4567 43499 4573
rect 44269 4607 44327 4613
rect 44269 4573 44281 4607
rect 44315 4604 44327 4607
rect 44358 4604 44364 4616
rect 44315 4576 44364 4604
rect 44315 4573 44327 4576
rect 44269 4567 44327 4573
rect 44358 4564 44364 4576
rect 44416 4564 44422 4616
rect 44453 4607 44511 4613
rect 44453 4573 44465 4607
rect 44499 4604 44511 4607
rect 44634 4604 44640 4616
rect 44499 4576 44640 4604
rect 44499 4573 44511 4576
rect 44453 4567 44511 4573
rect 44634 4564 44640 4576
rect 44692 4564 44698 4616
rect 45186 4604 45192 4616
rect 45147 4576 45192 4604
rect 45186 4564 45192 4576
rect 45244 4564 45250 4616
rect 48286 4604 48314 4644
rect 49329 4607 49387 4613
rect 49329 4604 49341 4607
rect 48286 4576 49341 4604
rect 49329 4573 49341 4576
rect 49375 4573 49387 4607
rect 49602 4604 49608 4616
rect 49563 4576 49608 4604
rect 49329 4567 49387 4573
rect 49602 4564 49608 4576
rect 49660 4564 49666 4616
rect 50154 4604 50160 4616
rect 50115 4576 50160 4604
rect 50154 4564 50160 4576
rect 50212 4564 50218 4616
rect 51046 4604 51074 4712
rect 53116 4681 53144 4780
rect 55674 4768 55680 4780
rect 55732 4768 55738 4820
rect 53101 4675 53159 4681
rect 53101 4641 53113 4675
rect 53147 4672 53159 4675
rect 53742 4672 53748 4684
rect 53147 4644 53748 4672
rect 53147 4641 53159 4644
rect 53101 4635 53159 4641
rect 53742 4632 53748 4644
rect 53800 4632 53806 4684
rect 51261 4607 51319 4613
rect 51261 4604 51273 4607
rect 51046 4576 51273 4604
rect 51261 4573 51273 4576
rect 51307 4604 51319 4607
rect 52825 4607 52883 4613
rect 52825 4604 52837 4607
rect 51307 4576 52837 4604
rect 51307 4573 51319 4576
rect 51261 4567 51319 4573
rect 52825 4573 52837 4576
rect 52871 4573 52883 4607
rect 54018 4604 54024 4616
rect 53979 4576 54024 4604
rect 52825 4567 52883 4573
rect 45097 4539 45155 4545
rect 45097 4536 45109 4539
rect 42090 4508 42472 4536
rect 38930 4468 38936 4480
rect 35860 4440 36860 4468
rect 38891 4440 38936 4468
rect 35860 4428 35866 4440
rect 38930 4428 38936 4440
rect 38988 4428 38994 4480
rect 40586 4468 40592 4480
rect 40547 4440 40592 4468
rect 40586 4428 40592 4440
rect 40644 4428 40650 4480
rect 42444 4468 42472 4508
rect 43548 4508 45109 4536
rect 43548 4468 43576 4508
rect 45097 4505 45109 4508
rect 45143 4505 45155 4539
rect 49878 4536 49884 4548
rect 47518 4508 49884 4536
rect 45097 4499 45155 4505
rect 49878 4496 49884 4508
rect 49936 4496 49942 4548
rect 42444 4440 43576 4468
rect 45554 4428 45560 4480
rect 45612 4468 45618 4480
rect 47765 4471 47823 4477
rect 47765 4468 47777 4471
rect 45612 4440 47777 4468
rect 45612 4428 45618 4440
rect 47765 4437 47777 4440
rect 47811 4437 47823 4471
rect 47765 4431 47823 4437
rect 50341 4471 50399 4477
rect 50341 4437 50353 4471
rect 50387 4468 50399 4471
rect 50890 4468 50896 4480
rect 50387 4440 50896 4468
rect 50387 4437 50399 4440
rect 50341 4431 50399 4437
rect 50890 4428 50896 4440
rect 50948 4428 50954 4480
rect 52086 4468 52092 4480
rect 52047 4440 52092 4468
rect 52086 4428 52092 4440
rect 52144 4428 52150 4480
rect 52840 4468 52868 4567
rect 54018 4564 54024 4576
rect 54076 4564 54082 4616
rect 55490 4604 55496 4616
rect 55451 4576 55496 4604
rect 55490 4564 55496 4576
rect 55548 4604 55554 4616
rect 56137 4607 56195 4613
rect 56137 4604 56149 4607
rect 55548 4576 56149 4604
rect 55548 4564 55554 4576
rect 56137 4573 56149 4576
rect 56183 4573 56195 4607
rect 56137 4567 56195 4573
rect 55309 4539 55367 4545
rect 55309 4536 55321 4539
rect 54128 4508 55321 4536
rect 54128 4468 54156 4508
rect 55309 4505 55321 4508
rect 55355 4505 55367 4539
rect 55309 4499 55367 4505
rect 54754 4468 54760 4480
rect 52840 4440 54156 4468
rect 54715 4440 54760 4468
rect 54754 4428 54760 4440
rect 54812 4428 54818 4480
rect 56594 4428 56600 4480
rect 56652 4468 56658 4480
rect 56689 4471 56747 4477
rect 56689 4468 56701 4471
rect 56652 4440 56701 4468
rect 56652 4428 56658 4440
rect 56689 4437 56701 4440
rect 56735 4437 56747 4471
rect 57238 4468 57244 4480
rect 57199 4440 57244 4468
rect 56689 4431 56747 4437
rect 57238 4428 57244 4440
rect 57296 4428 57302 4480
rect 1104 4378 58880 4400
rect 1104 4326 15398 4378
rect 15450 4326 15462 4378
rect 15514 4326 15526 4378
rect 15578 4326 15590 4378
rect 15642 4326 15654 4378
rect 15706 4326 29846 4378
rect 29898 4326 29910 4378
rect 29962 4326 29974 4378
rect 30026 4326 30038 4378
rect 30090 4326 30102 4378
rect 30154 4326 44294 4378
rect 44346 4326 44358 4378
rect 44410 4326 44422 4378
rect 44474 4326 44486 4378
rect 44538 4326 44550 4378
rect 44602 4326 58880 4378
rect 1104 4304 58880 4326
rect 3697 4267 3755 4273
rect 3697 4233 3709 4267
rect 3743 4264 3755 4267
rect 3786 4264 3792 4276
rect 3743 4236 3792 4264
rect 3743 4233 3755 4236
rect 3697 4227 3755 4233
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 10597 4267 10655 4273
rect 10597 4264 10609 4267
rect 10008 4236 10609 4264
rect 10008 4224 10014 4236
rect 10597 4233 10609 4236
rect 10643 4233 10655 4267
rect 10597 4227 10655 4233
rect 12406 4236 13400 4264
rect 2685 4199 2743 4205
rect 2685 4165 2697 4199
rect 2731 4196 2743 4199
rect 3142 4196 3148 4208
rect 2731 4168 3148 4196
rect 2731 4165 2743 4168
rect 2685 4159 2743 4165
rect 3142 4156 3148 4168
rect 3200 4156 3206 4208
rect 3234 4156 3240 4208
rect 3292 4196 3298 4208
rect 12406 4196 12434 4236
rect 13372 4205 13400 4236
rect 15286 4224 15292 4276
rect 15344 4264 15350 4276
rect 15378 4264 15384 4276
rect 15344 4236 15384 4264
rect 15344 4224 15350 4236
rect 15378 4224 15384 4236
rect 15436 4224 15442 4276
rect 15930 4224 15936 4276
rect 15988 4264 15994 4276
rect 17954 4264 17960 4276
rect 15988 4236 17960 4264
rect 15988 4224 15994 4236
rect 3292 4168 12434 4196
rect 13357 4199 13415 4205
rect 3292 4156 3298 4168
rect 13357 4165 13369 4199
rect 13403 4196 13415 4199
rect 13538 4196 13544 4208
rect 13403 4168 13544 4196
rect 13403 4165 13415 4168
rect 13357 4159 13415 4165
rect 13538 4156 13544 4168
rect 13596 4156 13602 4208
rect 16040 4205 16068 4236
rect 17954 4224 17960 4236
rect 18012 4224 18018 4276
rect 19242 4224 19248 4276
rect 19300 4224 19306 4276
rect 22738 4264 22744 4276
rect 19444 4236 22744 4264
rect 16025 4199 16083 4205
rect 15028 4168 15332 4196
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3418 4128 3424 4140
rect 2915 4100 3424 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 3786 4128 3792 4140
rect 3559 4100 3792 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 4154 4128 4160 4140
rect 4115 4100 4160 4128
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4246 4088 4252 4140
rect 4304 4128 4310 4140
rect 4413 4131 4471 4137
rect 4413 4128 4425 4131
rect 4304 4100 4425 4128
rect 4304 4088 4310 4100
rect 4413 4097 4425 4100
rect 4459 4097 4471 4131
rect 4413 4091 4471 4097
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 7282 4128 7288 4140
rect 6595 4100 7288 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 9122 4128 9128 4140
rect 7423 4100 9128 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9582 4088 9588 4140
rect 9640 4137 9646 4140
rect 9640 4128 9652 4137
rect 9858 4128 9864 4140
rect 9640 4100 9685 4128
rect 9819 4100 9864 4128
rect 9640 4091 9652 4100
rect 9640 4088 9646 4091
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 10778 4128 10784 4140
rect 10739 4100 10784 4128
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11790 4128 11796 4140
rect 11751 4100 11796 4128
rect 11790 4088 11796 4100
rect 11848 4088 11854 4140
rect 11885 4131 11943 4137
rect 11885 4097 11897 4131
rect 11931 4097 11943 4131
rect 11885 4091 11943 4097
rect 8754 4060 8760 4072
rect 6748 4032 8760 4060
rect 6748 4001 6776 4032
rect 8754 4020 8760 4032
rect 8812 4020 8818 4072
rect 10502 4020 10508 4072
rect 10560 4060 10566 4072
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10560 4032 10977 4060
rect 10560 4020 10566 4032
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 11514 4060 11520 4072
rect 11475 4032 11520 4060
rect 10965 4023 11023 4029
rect 11514 4020 11520 4032
rect 11572 4020 11578 4072
rect 11698 4020 11704 4072
rect 11756 4060 11762 4072
rect 11900 4060 11928 4091
rect 11974 4088 11980 4140
rect 12032 4128 12038 4140
rect 12032 4100 12077 4128
rect 12032 4088 12038 4100
rect 12158 4088 12164 4140
rect 12216 4128 12222 4140
rect 12216 4100 12261 4128
rect 12216 4088 12222 4100
rect 12618 4088 12624 4140
rect 12676 4128 12682 4140
rect 13081 4131 13139 4137
rect 13081 4128 13093 4131
rect 12676 4100 13093 4128
rect 12676 4088 12682 4100
rect 13081 4097 13093 4100
rect 13127 4097 13139 4131
rect 13081 4091 13139 4097
rect 11756 4032 11928 4060
rect 11756 4020 11762 4032
rect 6733 3995 6791 4001
rect 6733 3961 6745 3995
rect 6779 3961 6791 3995
rect 6733 3955 6791 3961
rect 8021 3995 8079 4001
rect 8021 3961 8033 3995
rect 8067 3992 8079 3995
rect 8846 3992 8852 4004
rect 8067 3964 8852 3992
rect 8067 3961 8079 3964
rect 8021 3955 8079 3961
rect 8846 3952 8852 3964
rect 8904 3952 8910 4004
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 12897 3995 12955 4001
rect 12897 3992 12909 3995
rect 11112 3964 12909 3992
rect 11112 3952 11118 3964
rect 12897 3961 12909 3964
rect 12943 3961 12955 3995
rect 13096 3992 13124 4091
rect 13170 4088 13176 4140
rect 13228 4128 13234 4140
rect 14645 4131 14703 4137
rect 13228 4100 13273 4128
rect 13228 4088 13234 4100
rect 14645 4097 14657 4131
rect 14691 4128 14703 4131
rect 15028 4128 15056 4168
rect 15304 4140 15332 4168
rect 16025 4165 16037 4199
rect 16071 4165 16083 4199
rect 17865 4199 17923 4205
rect 17865 4196 17877 4199
rect 16025 4159 16083 4165
rect 16684 4168 17877 4196
rect 14691 4100 15056 4128
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 15102 4088 15108 4140
rect 15160 4128 15166 4140
rect 15160 4100 15205 4128
rect 15160 4088 15166 4100
rect 15286 4088 15292 4140
rect 15344 4088 15350 4140
rect 15562 4088 15568 4140
rect 15620 4128 15626 4140
rect 15749 4131 15807 4137
rect 15749 4128 15761 4131
rect 15620 4100 15761 4128
rect 15620 4088 15626 4100
rect 15749 4097 15761 4100
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4128 15899 4131
rect 16114 4128 16120 4140
rect 15887 4100 16120 4128
rect 15887 4097 15899 4100
rect 15841 4091 15899 4097
rect 16114 4088 16120 4100
rect 16172 4128 16178 4140
rect 16482 4128 16488 4140
rect 16172 4100 16488 4128
rect 16172 4088 16178 4100
rect 16482 4088 16488 4100
rect 16540 4128 16546 4140
rect 16684 4128 16712 4168
rect 17865 4165 17877 4168
rect 17911 4165 17923 4199
rect 19260 4196 19288 4224
rect 17865 4159 17923 4165
rect 18800 4168 19288 4196
rect 18141 4131 18199 4137
rect 18141 4128 18153 4131
rect 16540 4100 16712 4128
rect 17880 4100 18153 4128
rect 16540 4088 16546 4100
rect 13188 4060 13216 4088
rect 13722 4060 13728 4072
rect 13188 4032 13728 4060
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 14001 4063 14059 4069
rect 14001 4029 14013 4063
rect 14047 4060 14059 4063
rect 16390 4060 16396 4072
rect 14047 4032 16396 4060
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 17880 4060 17908 4100
rect 18141 4097 18153 4100
rect 18187 4128 18199 4131
rect 18414 4128 18420 4140
rect 18187 4100 18420 4128
rect 18187 4097 18199 4100
rect 18141 4091 18199 4097
rect 18414 4088 18420 4100
rect 18472 4088 18478 4140
rect 18800 4137 18828 4168
rect 19334 4156 19340 4208
rect 19392 4196 19398 4208
rect 19444 4196 19472 4236
rect 22738 4224 22744 4236
rect 22796 4224 22802 4276
rect 30650 4224 30656 4276
rect 30708 4264 30714 4276
rect 31754 4264 31760 4276
rect 30708 4236 31760 4264
rect 30708 4224 30714 4236
rect 31754 4224 31760 4236
rect 31812 4264 31818 4276
rect 32582 4264 32588 4276
rect 31812 4236 32588 4264
rect 31812 4224 31818 4236
rect 32582 4224 32588 4236
rect 32640 4224 32646 4276
rect 34330 4224 34336 4276
rect 34388 4264 34394 4276
rect 34388 4236 35940 4264
rect 34388 4224 34394 4236
rect 19392 4168 19550 4196
rect 19392 4156 19398 4168
rect 23474 4156 23480 4208
rect 23532 4196 23538 4208
rect 28537 4199 28595 4205
rect 28537 4196 28549 4199
rect 23532 4168 28549 4196
rect 23532 4156 23538 4168
rect 28537 4165 28549 4168
rect 28583 4196 28595 4199
rect 28810 4196 28816 4208
rect 28583 4168 28816 4196
rect 28583 4165 28595 4168
rect 28537 4159 28595 4165
rect 28810 4156 28816 4168
rect 28868 4156 28874 4208
rect 31386 4156 31392 4208
rect 31444 4196 31450 4208
rect 35802 4196 35808 4208
rect 31444 4168 33456 4196
rect 34914 4168 35808 4196
rect 31444 4156 31450 4168
rect 33428 4140 33456 4168
rect 35802 4156 35808 4168
rect 35860 4156 35866 4208
rect 35912 4205 35940 4236
rect 39758 4224 39764 4276
rect 39816 4264 39822 4276
rect 44634 4264 44640 4276
rect 39816 4236 44640 4264
rect 39816 4224 39822 4236
rect 44634 4224 44640 4236
rect 44692 4224 44698 4276
rect 49602 4224 49608 4276
rect 49660 4264 49666 4276
rect 51077 4267 51135 4273
rect 51077 4264 51089 4267
rect 49660 4236 51089 4264
rect 49660 4224 49666 4236
rect 51077 4233 51089 4236
rect 51123 4264 51135 4267
rect 52454 4264 52460 4276
rect 51123 4236 52460 4264
rect 51123 4233 51135 4236
rect 51077 4227 51135 4233
rect 52454 4224 52460 4236
rect 52512 4224 52518 4276
rect 52638 4224 52644 4276
rect 52696 4264 52702 4276
rect 52696 4236 53144 4264
rect 52696 4224 52702 4236
rect 35897 4199 35955 4205
rect 35897 4165 35909 4199
rect 35943 4165 35955 4199
rect 49050 4196 49056 4208
rect 35897 4159 35955 4165
rect 39224 4168 40250 4196
rect 43916 4168 47886 4196
rect 49011 4168 49056 4196
rect 18785 4131 18843 4137
rect 18785 4097 18797 4131
rect 18831 4097 18843 4131
rect 18785 4091 18843 4097
rect 21174 4088 21180 4140
rect 21232 4128 21238 4140
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 21232 4100 21833 4128
rect 21232 4088 21238 4100
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 22002 4128 22008 4140
rect 21963 4100 22008 4128
rect 21821 4091 21879 4097
rect 22002 4088 22008 4100
rect 22060 4088 22066 4140
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 16546 4032 17908 4060
rect 16546 3992 16574 4032
rect 17954 4020 17960 4072
rect 18012 4060 18018 4072
rect 18322 4060 18328 4072
rect 18012 4032 18328 4060
rect 18012 4020 18018 4032
rect 18322 4020 18328 4032
rect 18380 4020 18386 4072
rect 19058 4060 19064 4072
rect 19019 4032 19064 4060
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 22112 4060 22140 4091
rect 22186 4088 22192 4140
rect 22244 4128 22250 4140
rect 23569 4131 23627 4137
rect 22244 4100 22289 4128
rect 22244 4088 22250 4100
rect 23569 4097 23581 4131
rect 23615 4128 23627 4131
rect 23842 4128 23848 4140
rect 23615 4100 23848 4128
rect 23615 4097 23627 4100
rect 23569 4091 23627 4097
rect 23842 4088 23848 4100
rect 23900 4088 23906 4140
rect 24118 4128 24124 4140
rect 24079 4100 24124 4128
rect 24118 4088 24124 4100
rect 24176 4088 24182 4140
rect 24377 4131 24435 4137
rect 24377 4128 24389 4131
rect 24228 4100 24389 4128
rect 20772 4032 22140 4060
rect 22465 4063 22523 4069
rect 20772 4020 20778 4032
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 24228 4060 24256 4100
rect 24377 4097 24389 4100
rect 24423 4097 24435 4131
rect 24377 4091 24435 4097
rect 26237 4131 26295 4137
rect 26237 4097 26249 4131
rect 26283 4128 26295 4131
rect 26326 4128 26332 4140
rect 26283 4100 26332 4128
rect 26283 4097 26295 4100
rect 26237 4091 26295 4097
rect 26326 4088 26332 4100
rect 26384 4088 26390 4140
rect 30745 4131 30803 4137
rect 30745 4097 30757 4131
rect 30791 4128 30803 4131
rect 30926 4128 30932 4140
rect 30791 4100 30932 4128
rect 30791 4097 30803 4100
rect 30745 4091 30803 4097
rect 30926 4088 30932 4100
rect 30984 4088 30990 4140
rect 32582 4128 32588 4140
rect 32543 4100 32588 4128
rect 32582 4088 32588 4100
rect 32640 4088 32646 4140
rect 33410 4128 33416 4140
rect 33371 4100 33416 4128
rect 33410 4088 33416 4100
rect 33468 4088 33474 4140
rect 37550 4088 37556 4140
rect 37608 4128 37614 4140
rect 38197 4131 38255 4137
rect 38197 4128 38209 4131
rect 37608 4100 38209 4128
rect 37608 4088 37614 4100
rect 38197 4097 38209 4100
rect 38243 4097 38255 4131
rect 39114 4128 39120 4140
rect 39027 4100 39120 4128
rect 38197 4091 38255 4097
rect 39114 4088 39120 4100
rect 39172 4088 39178 4140
rect 39224 4137 39252 4168
rect 39209 4131 39267 4137
rect 39209 4097 39221 4131
rect 39255 4097 39267 4131
rect 39209 4091 39267 4097
rect 41690 4088 41696 4140
rect 41748 4128 41754 4140
rect 42889 4131 42947 4137
rect 41748 4100 41793 4128
rect 41748 4088 41754 4100
rect 42889 4097 42901 4131
rect 42935 4128 42947 4131
rect 42978 4128 42984 4140
rect 42935 4100 42984 4128
rect 42935 4097 42947 4100
rect 42889 4091 42947 4097
rect 42978 4088 42984 4100
rect 43036 4088 43042 4140
rect 43916 4137 43944 4168
rect 49050 4156 49056 4168
rect 49108 4156 49114 4208
rect 53006 4196 53012 4208
rect 52967 4168 53012 4196
rect 53006 4156 53012 4168
rect 53064 4156 53070 4208
rect 53116 4196 53144 4236
rect 53650 4224 53656 4276
rect 53708 4264 53714 4276
rect 54754 4264 54760 4276
rect 53708 4236 54760 4264
rect 53708 4224 53714 4236
rect 54754 4224 54760 4236
rect 54812 4264 54818 4276
rect 55033 4267 55091 4273
rect 55033 4264 55045 4267
rect 54812 4236 55045 4264
rect 54812 4224 54818 4236
rect 55033 4233 55045 4236
rect 55079 4233 55091 4267
rect 55033 4227 55091 4233
rect 53116 4168 53498 4196
rect 43809 4131 43867 4137
rect 43809 4097 43821 4131
rect 43855 4097 43867 4131
rect 43809 4091 43867 4097
rect 43901 4131 43959 4137
rect 43901 4097 43913 4131
rect 43947 4097 43959 4131
rect 45738 4128 45744 4140
rect 45699 4100 45744 4128
rect 43901 4091 43959 4097
rect 30374 4060 30380 4072
rect 22511 4032 24256 4060
rect 25424 4032 30380 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 13096 3964 15332 3992
rect 12897 3955 12955 3961
rect 2133 3927 2191 3933
rect 2133 3893 2145 3927
rect 2179 3924 2191 3927
rect 3050 3924 3056 3936
rect 2179 3896 3056 3924
rect 2179 3893 2191 3896
rect 2133 3887 2191 3893
rect 3050 3884 3056 3896
rect 3108 3884 3114 3936
rect 4154 3884 4160 3936
rect 4212 3924 4218 3936
rect 5537 3927 5595 3933
rect 5537 3924 5549 3927
rect 4212 3896 5549 3924
rect 4212 3884 4218 3896
rect 5537 3893 5549 3896
rect 5583 3924 5595 3927
rect 8386 3924 8392 3936
rect 5583 3896 8392 3924
rect 5583 3893 5595 3896
rect 5537 3887 5595 3893
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 8938 3924 8944 3936
rect 8527 3896 8944 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9582 3924 9588 3936
rect 9272 3896 9588 3924
rect 9272 3884 9278 3896
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 11422 3924 11428 3936
rect 11020 3896 11428 3924
rect 11020 3884 11026 3896
rect 11422 3884 11428 3896
rect 11480 3884 11486 3936
rect 12618 3884 12624 3936
rect 12676 3924 12682 3936
rect 12986 3924 12992 3936
rect 12676 3896 12992 3924
rect 12676 3884 12682 3896
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13078 3884 13084 3936
rect 13136 3924 13142 3936
rect 13136 3896 13181 3924
rect 13136 3884 13142 3896
rect 13354 3884 13360 3936
rect 13412 3924 13418 3936
rect 15102 3924 15108 3936
rect 13412 3896 15108 3924
rect 13412 3884 13418 3896
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15304 3933 15332 3964
rect 15856 3964 16574 3992
rect 17405 3995 17463 4001
rect 15289 3927 15347 3933
rect 15289 3893 15301 3927
rect 15335 3924 15347 3927
rect 15856 3924 15884 3964
rect 17405 3961 17417 3995
rect 17451 3992 17463 3995
rect 22554 3992 22560 4004
rect 17451 3964 18000 3992
rect 17451 3961 17463 3964
rect 17405 3955 17463 3961
rect 17972 3936 18000 3964
rect 20456 3964 22560 3992
rect 15335 3896 15884 3924
rect 15933 3927 15991 3933
rect 15335 3893 15347 3896
rect 15289 3887 15347 3893
rect 15933 3893 15945 3927
rect 15979 3924 15991 3927
rect 17862 3924 17868 3936
rect 15979 3896 17868 3924
rect 15979 3893 15991 3896
rect 15933 3887 15991 3893
rect 17862 3884 17868 3896
rect 17920 3884 17926 3936
rect 17954 3884 17960 3936
rect 18012 3884 18018 3936
rect 18141 3927 18199 3933
rect 18141 3893 18153 3927
rect 18187 3924 18199 3927
rect 18230 3924 18236 3936
rect 18187 3896 18236 3924
rect 18187 3893 18199 3896
rect 18141 3887 18199 3893
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 18325 3927 18383 3933
rect 18325 3893 18337 3927
rect 18371 3924 18383 3927
rect 20456 3924 20484 3964
rect 22554 3952 22560 3964
rect 22612 3952 22618 4004
rect 18371 3896 20484 3924
rect 20533 3927 20591 3933
rect 18371 3893 18383 3896
rect 18325 3887 18383 3893
rect 20533 3893 20545 3927
rect 20579 3924 20591 3927
rect 21082 3924 21088 3936
rect 20579 3896 21088 3924
rect 20579 3893 20591 3896
rect 20533 3887 20591 3893
rect 21082 3884 21088 3896
rect 21140 3884 21146 3936
rect 21269 3927 21327 3933
rect 21269 3893 21281 3927
rect 21315 3924 21327 3927
rect 21818 3924 21824 3936
rect 21315 3896 21824 3924
rect 21315 3893 21327 3896
rect 21269 3887 21327 3893
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 23198 3884 23204 3936
rect 23256 3924 23262 3936
rect 23385 3927 23443 3933
rect 23385 3924 23397 3927
rect 23256 3896 23397 3924
rect 23256 3884 23262 3896
rect 23385 3893 23397 3896
rect 23431 3893 23443 3927
rect 23385 3887 23443 3893
rect 24302 3884 24308 3936
rect 24360 3924 24366 3936
rect 25424 3924 25452 4032
rect 30374 4020 30380 4032
rect 30432 4020 30438 4072
rect 33689 4063 33747 4069
rect 33689 4060 33701 4063
rect 31726 4032 33701 4060
rect 25498 3952 25504 4004
rect 25556 3992 25562 4004
rect 28077 3995 28135 4001
rect 25556 3964 25601 3992
rect 25556 3952 25562 3964
rect 28077 3961 28089 3995
rect 28123 3992 28135 3995
rect 29730 3992 29736 4004
rect 28123 3964 29736 3992
rect 28123 3961 28135 3964
rect 28077 3955 28135 3961
rect 29730 3952 29736 3964
rect 29788 3952 29794 4004
rect 30929 3995 30987 4001
rect 30929 3961 30941 3995
rect 30975 3992 30987 3995
rect 31726 3992 31754 4032
rect 33689 4029 33701 4032
rect 33735 4029 33747 4063
rect 33689 4023 33747 4029
rect 35894 4020 35900 4072
rect 35952 4060 35958 4072
rect 37277 4063 37335 4069
rect 37277 4060 37289 4063
rect 35952 4032 37289 4060
rect 35952 4020 35958 4032
rect 37277 4029 37289 4032
rect 37323 4029 37335 4063
rect 37277 4023 37335 4029
rect 32766 3992 32772 4004
rect 30975 3964 31754 3992
rect 32727 3964 32772 3992
rect 30975 3961 30987 3964
rect 30929 3955 30987 3961
rect 32766 3952 32772 3964
rect 32824 3952 32830 4004
rect 35618 3952 35624 4004
rect 35676 3992 35682 4004
rect 36541 3995 36599 4001
rect 36541 3992 36553 3995
rect 35676 3964 36553 3992
rect 35676 3952 35682 3964
rect 36541 3961 36553 3964
rect 36587 3961 36599 3995
rect 36541 3955 36599 3961
rect 37458 3952 37464 4004
rect 37516 3992 37522 4004
rect 37553 3995 37611 4001
rect 37553 3992 37565 3995
rect 37516 3964 37565 3992
rect 37516 3952 37522 3964
rect 37553 3961 37565 3964
rect 37599 3961 37611 3995
rect 39132 3992 39160 4088
rect 40126 4020 40132 4072
rect 40184 4060 40190 4072
rect 41417 4063 41475 4069
rect 41417 4060 41429 4063
rect 40184 4032 41429 4060
rect 40184 4020 40190 4032
rect 41417 4029 41429 4032
rect 41463 4029 41475 4063
rect 43824 4060 43852 4091
rect 45738 4088 45744 4100
rect 45796 4088 45802 4140
rect 46569 4131 46627 4137
rect 46569 4097 46581 4131
rect 46615 4097 46627 4131
rect 46569 4091 46627 4097
rect 45186 4060 45192 4072
rect 41417 4023 41475 4029
rect 42904 4032 45192 4060
rect 39132 3964 40080 3992
rect 37553 3955 37611 3961
rect 26418 3924 26424 3936
rect 24360 3896 25452 3924
rect 26379 3896 26424 3924
rect 24360 3884 24366 3896
rect 26418 3884 26424 3896
rect 26476 3884 26482 3936
rect 27157 3927 27215 3933
rect 27157 3893 27169 3927
rect 27203 3924 27215 3927
rect 27890 3924 27896 3936
rect 27203 3896 27896 3924
rect 27203 3893 27215 3896
rect 27157 3887 27215 3893
rect 27890 3884 27896 3896
rect 27948 3884 27954 3936
rect 28626 3884 28632 3936
rect 28684 3924 28690 3936
rect 29825 3927 29883 3933
rect 29825 3924 29837 3927
rect 28684 3896 29837 3924
rect 28684 3884 28690 3896
rect 29825 3893 29837 3896
rect 29871 3893 29883 3927
rect 31386 3924 31392 3936
rect 31347 3896 31392 3924
rect 29825 3887 29883 3893
rect 31386 3884 31392 3896
rect 31444 3884 31450 3936
rect 35158 3924 35164 3936
rect 35119 3896 35164 3924
rect 35158 3884 35164 3896
rect 35216 3884 35222 3936
rect 35986 3924 35992 3936
rect 35899 3896 35992 3924
rect 35986 3884 35992 3896
rect 36044 3924 36050 3936
rect 36354 3924 36360 3936
rect 36044 3896 36360 3924
rect 36044 3884 36050 3896
rect 36354 3884 36360 3896
rect 36412 3884 36418 3936
rect 37734 3924 37740 3936
rect 37695 3896 37740 3924
rect 37734 3884 37740 3896
rect 37792 3884 37798 3936
rect 39758 3884 39764 3936
rect 39816 3924 39822 3936
rect 39945 3927 40003 3933
rect 39945 3924 39957 3927
rect 39816 3896 39957 3924
rect 39816 3884 39822 3896
rect 39945 3893 39957 3896
rect 39991 3893 40003 3927
rect 40052 3924 40080 3964
rect 42904 3924 42932 4032
rect 45186 4020 45192 4032
rect 45244 4060 45250 4072
rect 46584 4060 46612 4091
rect 49326 4088 49332 4140
rect 49384 4128 49390 4140
rect 49694 4128 49700 4140
rect 49384 4100 49700 4128
rect 49384 4088 49390 4100
rect 49694 4088 49700 4100
rect 49752 4088 49758 4140
rect 49786 4088 49792 4140
rect 49844 4128 49850 4140
rect 51261 4131 51319 4137
rect 49844 4100 49889 4128
rect 49844 4088 49850 4100
rect 51261 4097 51273 4131
rect 51307 4128 51319 4131
rect 51350 4128 51356 4140
rect 51307 4100 51356 4128
rect 51307 4097 51319 4100
rect 51261 4091 51319 4097
rect 51350 4088 51356 4100
rect 51408 4088 51414 4140
rect 52178 4088 52184 4140
rect 52236 4128 52242 4140
rect 52733 4131 52791 4137
rect 52733 4128 52745 4131
rect 52236 4100 52745 4128
rect 52236 4088 52242 4100
rect 52733 4097 52745 4100
rect 52779 4097 52791 4131
rect 52733 4091 52791 4097
rect 55306 4088 55312 4140
rect 55364 4128 55370 4140
rect 55861 4131 55919 4137
rect 55861 4128 55873 4131
rect 55364 4100 55873 4128
rect 55364 4088 55370 4100
rect 55861 4097 55873 4100
rect 55907 4097 55919 4131
rect 56686 4128 56692 4140
rect 56599 4100 56692 4128
rect 55861 4091 55919 4097
rect 56686 4088 56692 4100
rect 56744 4128 56750 4140
rect 57238 4128 57244 4140
rect 56744 4100 57244 4128
rect 56744 4088 56750 4100
rect 57238 4088 57244 4100
rect 57296 4088 57302 4140
rect 45244 4032 46612 4060
rect 45244 4020 45250 4032
rect 47026 4020 47032 4072
rect 47084 4060 47090 4072
rect 49602 4060 49608 4072
rect 47084 4032 49608 4060
rect 47084 4020 47090 4032
rect 49602 4020 49608 4032
rect 49660 4060 49666 4072
rect 53650 4060 53656 4072
rect 49660 4032 53656 4060
rect 49660 4020 49666 4032
rect 53650 4020 53656 4032
rect 53708 4020 53714 4072
rect 53742 4020 53748 4072
rect 53800 4060 53806 4072
rect 55585 4063 55643 4069
rect 55585 4060 55597 4063
rect 53800 4032 55597 4060
rect 53800 4020 53806 4032
rect 55585 4029 55597 4032
rect 55631 4029 55643 4063
rect 55585 4023 55643 4029
rect 44174 3952 44180 4004
rect 44232 3992 44238 4004
rect 45097 3995 45155 4001
rect 45097 3992 45109 3995
rect 44232 3964 45109 3992
rect 44232 3952 44238 3964
rect 45097 3961 45109 3964
rect 45143 3961 45155 3995
rect 49878 3992 49884 4004
rect 49839 3964 49884 3992
rect 45097 3955 45155 3961
rect 49878 3952 49884 3964
rect 49936 3952 49942 4004
rect 49970 3952 49976 4004
rect 50028 3992 50034 4004
rect 51721 3995 51779 4001
rect 51721 3992 51733 3995
rect 50028 3964 51733 3992
rect 50028 3952 50034 3964
rect 51721 3961 51733 3964
rect 51767 3961 51779 3995
rect 55214 3992 55220 4004
rect 51721 3955 51779 3961
rect 54496 3964 55220 3992
rect 54496 3936 54524 3964
rect 55214 3952 55220 3964
rect 55272 3952 55278 4004
rect 43070 3924 43076 3936
rect 40052 3896 42932 3924
rect 43031 3896 43076 3924
rect 39945 3887 40003 3893
rect 43070 3884 43076 3896
rect 43128 3884 43134 3936
rect 43622 3884 43628 3936
rect 43680 3924 43686 3936
rect 44453 3927 44511 3933
rect 44453 3924 44465 3927
rect 43680 3896 44465 3924
rect 43680 3884 43686 3896
rect 44453 3893 44465 3896
rect 44499 3893 44511 3927
rect 45922 3924 45928 3936
rect 45883 3896 45928 3924
rect 44453 3887 44511 3893
rect 45922 3884 45928 3896
rect 45980 3884 45986 3936
rect 46658 3924 46664 3936
rect 46619 3896 46664 3924
rect 46658 3884 46664 3896
rect 46716 3884 46722 3936
rect 47578 3924 47584 3936
rect 47539 3896 47584 3924
rect 47578 3884 47584 3896
rect 47636 3884 47642 3936
rect 47762 3884 47768 3936
rect 47820 3924 47826 3936
rect 50433 3927 50491 3933
rect 50433 3924 50445 3927
rect 47820 3896 50445 3924
rect 47820 3884 47826 3896
rect 50433 3893 50445 3896
rect 50479 3893 50491 3927
rect 54478 3924 54484 3936
rect 54439 3896 54484 3924
rect 50433 3887 50491 3893
rect 54478 3884 54484 3896
rect 54536 3884 54542 3936
rect 55306 3884 55312 3936
rect 55364 3924 55370 3936
rect 55674 3924 55680 3936
rect 55364 3896 55680 3924
rect 55364 3884 55370 3896
rect 55674 3884 55680 3896
rect 55732 3924 55738 3936
rect 56318 3924 56324 3936
rect 55732 3896 56324 3924
rect 55732 3884 55738 3896
rect 56318 3884 56324 3896
rect 56376 3924 56382 3936
rect 57241 3927 57299 3933
rect 57241 3924 57253 3927
rect 56376 3896 57253 3924
rect 56376 3884 56382 3896
rect 57241 3893 57253 3896
rect 57287 3924 57299 3927
rect 57885 3927 57943 3933
rect 57885 3924 57897 3927
rect 57287 3896 57897 3924
rect 57287 3893 57299 3896
rect 57241 3887 57299 3893
rect 57885 3893 57897 3896
rect 57931 3893 57943 3927
rect 57885 3887 57943 3893
rect 1104 3834 58880 3856
rect 1104 3782 8174 3834
rect 8226 3782 8238 3834
rect 8290 3782 8302 3834
rect 8354 3782 8366 3834
rect 8418 3782 8430 3834
rect 8482 3782 22622 3834
rect 22674 3782 22686 3834
rect 22738 3782 22750 3834
rect 22802 3782 22814 3834
rect 22866 3782 22878 3834
rect 22930 3782 37070 3834
rect 37122 3782 37134 3834
rect 37186 3782 37198 3834
rect 37250 3782 37262 3834
rect 37314 3782 37326 3834
rect 37378 3782 51518 3834
rect 51570 3782 51582 3834
rect 51634 3782 51646 3834
rect 51698 3782 51710 3834
rect 51762 3782 51774 3834
rect 51826 3782 58880 3834
rect 1104 3760 58880 3782
rect 3786 3720 3792 3732
rect 3747 3692 3792 3720
rect 3786 3680 3792 3692
rect 3844 3680 3850 3732
rect 6362 3720 6368 3732
rect 6323 3692 6368 3720
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 8846 3680 8852 3732
rect 8904 3720 8910 3732
rect 9766 3720 9772 3732
rect 8904 3692 9772 3720
rect 8904 3680 8910 3692
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 11793 3723 11851 3729
rect 11793 3720 11805 3723
rect 10836 3692 11805 3720
rect 10836 3680 10842 3692
rect 11793 3689 11805 3692
rect 11839 3689 11851 3723
rect 14366 3720 14372 3732
rect 11793 3683 11851 3689
rect 13648 3692 14372 3720
rect 7650 3652 7656 3664
rect 2746 3624 7656 3652
rect 1489 3587 1547 3593
rect 1489 3553 1501 3587
rect 1535 3584 1547 3587
rect 2406 3584 2412 3596
rect 1535 3556 2412 3584
rect 1535 3553 1547 3556
rect 1489 3547 1547 3553
rect 2406 3544 2412 3556
rect 2464 3584 2470 3596
rect 2746 3584 2774 3624
rect 7650 3612 7656 3624
rect 7708 3612 7714 3664
rect 9125 3655 9183 3661
rect 9125 3621 9137 3655
rect 9171 3652 9183 3655
rect 13078 3652 13084 3664
rect 9171 3624 13084 3652
rect 9171 3621 9183 3624
rect 9125 3615 9183 3621
rect 13078 3612 13084 3624
rect 13136 3612 13142 3664
rect 2464 3556 2774 3584
rect 2884 3556 3188 3584
rect 2464 3544 2470 3556
rect 2593 3451 2651 3457
rect 2593 3417 2605 3451
rect 2639 3448 2651 3451
rect 2884 3448 2912 3556
rect 2958 3476 2964 3528
rect 3016 3518 3022 3528
rect 3053 3519 3111 3525
rect 3053 3518 3065 3519
rect 3016 3490 3065 3518
rect 3016 3476 3022 3490
rect 3053 3485 3065 3490
rect 3099 3485 3111 3519
rect 3160 3516 3188 3556
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 4212 3556 4261 3584
rect 4212 3544 4218 3556
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 4430 3584 4436 3596
rect 4391 3556 4436 3584
rect 4249 3547 4307 3553
rect 4430 3544 4436 3556
rect 4488 3544 4494 3596
rect 5442 3544 5448 3596
rect 5500 3584 5506 3596
rect 6273 3587 6331 3593
rect 5500 3556 6132 3584
rect 5500 3544 5506 3556
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 3160 3488 5273 3516
rect 3053 3479 3111 3485
rect 5261 3485 5273 3488
rect 5307 3516 5319 3519
rect 6104 3516 6132 3556
rect 6273 3553 6285 3587
rect 6319 3584 6331 3587
rect 7190 3584 7196 3596
rect 6319 3556 7196 3584
rect 6319 3553 6331 3556
rect 6273 3547 6331 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 8570 3544 8576 3596
rect 8628 3584 8634 3596
rect 8846 3584 8852 3596
rect 8628 3556 8852 3584
rect 8628 3544 8634 3556
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 9861 3587 9919 3593
rect 9861 3553 9873 3587
rect 9907 3584 9919 3587
rect 12158 3584 12164 3596
rect 9907 3556 12164 3584
rect 9907 3553 9919 3556
rect 9861 3547 9919 3553
rect 12158 3544 12164 3556
rect 12216 3544 12222 3596
rect 12342 3584 12348 3596
rect 12303 3556 12348 3584
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 6365 3519 6423 3525
rect 6365 3516 6377 3519
rect 5307 3488 6040 3516
rect 6104 3488 6377 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 2639 3420 2912 3448
rect 3068 3420 4200 3448
rect 2639 3417 2651 3420
rect 2593 3411 2651 3417
rect 2041 3383 2099 3389
rect 2041 3349 2053 3383
rect 2087 3380 2099 3383
rect 3068 3380 3096 3420
rect 2087 3352 3096 3380
rect 2087 3349 2099 3352
rect 2041 3343 2099 3349
rect 3142 3340 3148 3392
rect 3200 3380 3206 3392
rect 4172 3389 4200 3420
rect 5534 3408 5540 3460
rect 5592 3448 5598 3460
rect 5905 3451 5963 3457
rect 5905 3448 5917 3451
rect 5592 3420 5917 3448
rect 5592 3408 5598 3420
rect 5905 3417 5917 3420
rect 5951 3417 5963 3451
rect 6012 3448 6040 3488
rect 6365 3485 6377 3488
rect 6411 3516 6423 3519
rect 6638 3516 6644 3528
rect 6411 3488 6644 3516
rect 6411 3485 6423 3488
rect 6365 3479 6423 3485
rect 6638 3476 6644 3488
rect 6696 3476 6702 3528
rect 7098 3476 7104 3528
rect 7156 3476 7162 3528
rect 7742 3516 7748 3528
rect 7703 3488 7748 3516
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 10226 3516 10232 3528
rect 8435 3488 10232 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10502 3476 10508 3528
rect 10560 3516 10566 3528
rect 10597 3519 10655 3525
rect 10597 3516 10609 3519
rect 10560 3488 10609 3516
rect 10560 3476 10566 3488
rect 10597 3485 10609 3488
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 10689 3519 10747 3525
rect 10689 3485 10701 3519
rect 10735 3485 10747 3519
rect 10689 3479 10747 3485
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3516 11391 3519
rect 12986 3516 12992 3528
rect 11379 3488 12992 3516
rect 11379 3485 11391 3488
rect 11333 3479 11391 3485
rect 7116 3448 7144 3476
rect 9674 3448 9680 3460
rect 6012 3420 7144 3448
rect 9635 3420 9680 3448
rect 5905 3411 5963 3417
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 10410 3448 10416 3460
rect 10371 3420 10416 3448
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 10704 3448 10732 3479
rect 12986 3476 12992 3488
rect 13044 3476 13050 3528
rect 13648 3516 13676 3692
rect 14366 3680 14372 3692
rect 14424 3720 14430 3732
rect 14461 3723 14519 3729
rect 14461 3720 14473 3723
rect 14424 3692 14473 3720
rect 14424 3680 14430 3692
rect 14461 3689 14473 3692
rect 14507 3689 14519 3723
rect 15378 3720 15384 3732
rect 15291 3692 15384 3720
rect 14461 3683 14519 3689
rect 15378 3680 15384 3692
rect 15436 3720 15442 3732
rect 15933 3723 15991 3729
rect 15933 3720 15945 3723
rect 15436 3692 15945 3720
rect 15436 3680 15442 3692
rect 15933 3689 15945 3692
rect 15979 3689 15991 3723
rect 17586 3720 17592 3732
rect 15933 3683 15991 3689
rect 16040 3692 17592 3720
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 15396 3652 15424 3680
rect 13780 3624 15424 3652
rect 15473 3655 15531 3661
rect 13780 3612 13786 3624
rect 15473 3621 15485 3655
rect 15519 3652 15531 3655
rect 16040 3652 16068 3692
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 17862 3680 17868 3732
rect 17920 3720 17926 3732
rect 18230 3720 18236 3732
rect 17920 3692 18236 3720
rect 17920 3680 17926 3692
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 18693 3723 18751 3729
rect 18693 3689 18705 3723
rect 18739 3720 18751 3723
rect 19150 3720 19156 3732
rect 18739 3692 19156 3720
rect 18739 3689 18751 3692
rect 18693 3683 18751 3689
rect 19150 3680 19156 3692
rect 19208 3680 19214 3732
rect 22002 3720 22008 3732
rect 19812 3692 22008 3720
rect 15519 3624 16068 3652
rect 16393 3655 16451 3661
rect 15519 3621 15531 3624
rect 15473 3615 15531 3621
rect 16393 3621 16405 3655
rect 16439 3621 16451 3655
rect 16393 3615 16451 3621
rect 17773 3655 17831 3661
rect 17773 3621 17785 3655
rect 17819 3652 17831 3655
rect 19610 3652 19616 3664
rect 17819 3624 19616 3652
rect 17819 3621 17831 3624
rect 17773 3615 17831 3621
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 14251 3587 14309 3593
rect 14251 3584 14263 3587
rect 13964 3556 14263 3584
rect 13964 3544 13970 3556
rect 14251 3553 14263 3556
rect 14297 3553 14309 3587
rect 14251 3547 14309 3553
rect 15654 3544 15660 3596
rect 15712 3584 15718 3596
rect 16025 3587 16083 3593
rect 16025 3584 16037 3587
rect 15712 3556 16037 3584
rect 15712 3544 15718 3556
rect 16025 3553 16037 3556
rect 16071 3584 16083 3587
rect 16114 3584 16120 3596
rect 16071 3556 16120 3584
rect 16071 3553 16083 3556
rect 16025 3547 16083 3553
rect 16114 3544 16120 3556
rect 16172 3544 16178 3596
rect 14090 3516 14096 3528
rect 13096 3488 13676 3516
rect 14051 3488 14096 3516
rect 13096 3448 13124 3488
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 14550 3516 14556 3528
rect 14507 3488 14556 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 14550 3476 14556 3488
rect 14608 3476 14614 3528
rect 14645 3519 14703 3525
rect 14645 3485 14657 3519
rect 14691 3485 14703 3519
rect 14645 3479 14703 3485
rect 10704 3420 13124 3448
rect 13170 3408 13176 3460
rect 13228 3448 13234 3460
rect 13228 3420 13492 3448
rect 13228 3408 13234 3420
rect 4157 3383 4215 3389
rect 3200 3352 3245 3380
rect 3200 3340 3206 3352
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 4522 3380 4528 3392
rect 4203 3352 4528 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 4522 3340 4528 3352
rect 4580 3340 4586 3392
rect 5442 3380 5448 3392
rect 5403 3352 5448 3380
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 6546 3380 6552 3392
rect 6507 3352 6552 3380
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 7101 3383 7159 3389
rect 7101 3349 7113 3383
rect 7147 3380 7159 3383
rect 8294 3380 8300 3392
rect 7147 3352 8300 3380
rect 7147 3349 7159 3352
rect 7101 3343 7159 3349
rect 8294 3340 8300 3352
rect 8352 3340 8358 3392
rect 10686 3380 10692 3392
rect 10647 3352 10692 3380
rect 10686 3340 10692 3352
rect 10744 3340 10750 3392
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 12158 3380 12164 3392
rect 11664 3352 12164 3380
rect 11664 3340 11670 3352
rect 12158 3340 12164 3352
rect 12216 3340 12222 3392
rect 12250 3340 12256 3392
rect 12308 3380 12314 3392
rect 12308 3352 12353 3380
rect 12308 3340 12314 3352
rect 12618 3340 12624 3392
rect 12676 3380 12682 3392
rect 13081 3383 13139 3389
rect 13081 3380 13093 3383
rect 12676 3352 13093 3380
rect 12676 3340 12682 3352
rect 13081 3349 13093 3352
rect 13127 3349 13139 3383
rect 13464 3380 13492 3420
rect 13538 3408 13544 3460
rect 13596 3448 13602 3460
rect 14660 3448 14688 3479
rect 15102 3476 15108 3528
rect 15160 3516 15166 3528
rect 16209 3519 16267 3525
rect 16209 3516 16221 3519
rect 15160 3488 16221 3516
rect 15160 3476 15166 3488
rect 16209 3485 16221 3488
rect 16255 3485 16267 3519
rect 16209 3479 16267 3485
rect 15562 3448 15568 3460
rect 13596 3420 15568 3448
rect 13596 3408 13602 3420
rect 15562 3408 15568 3420
rect 15620 3448 15626 3460
rect 15933 3451 15991 3457
rect 15933 3448 15945 3451
rect 15620 3420 15945 3448
rect 15620 3408 15626 3420
rect 15933 3417 15945 3420
rect 15979 3417 15991 3451
rect 16408 3448 16436 3615
rect 19610 3612 19616 3624
rect 19668 3612 19674 3664
rect 17129 3587 17187 3593
rect 17129 3553 17141 3587
rect 17175 3584 17187 3587
rect 18046 3584 18052 3596
rect 17175 3556 18052 3584
rect 17175 3553 17187 3556
rect 17129 3547 17187 3553
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 18322 3584 18328 3596
rect 18283 3556 18328 3584
rect 18322 3544 18328 3556
rect 18380 3544 18386 3596
rect 19702 3584 19708 3596
rect 18432 3556 19334 3584
rect 19663 3556 19708 3584
rect 18432 3516 18460 3556
rect 17880 3488 18460 3516
rect 17880 3448 17908 3488
rect 18506 3476 18512 3528
rect 18564 3516 18570 3528
rect 19306 3516 19334 3556
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 19812 3516 19840 3692
rect 22002 3680 22008 3692
rect 22060 3680 22066 3732
rect 25314 3720 25320 3732
rect 25275 3692 25320 3720
rect 25314 3680 25320 3692
rect 25372 3680 25378 3732
rect 30926 3720 30932 3732
rect 26344 3692 29684 3720
rect 30887 3692 30932 3720
rect 20349 3655 20407 3661
rect 20349 3621 20361 3655
rect 20395 3621 20407 3655
rect 20349 3615 20407 3621
rect 18564 3488 18609 3516
rect 19306 3488 19840 3516
rect 20364 3516 20392 3615
rect 24578 3612 24584 3664
rect 24636 3652 24642 3664
rect 26344 3652 26372 3692
rect 24636 3624 26372 3652
rect 24636 3612 24642 3624
rect 26418 3612 26424 3664
rect 26476 3652 26482 3664
rect 26476 3624 27384 3652
rect 26476 3612 26482 3624
rect 21174 3584 21180 3596
rect 21135 3556 21180 3584
rect 21174 3544 21180 3556
rect 21232 3544 21238 3596
rect 24765 3587 24823 3593
rect 24765 3553 24777 3587
rect 24811 3584 24823 3587
rect 26142 3584 26148 3596
rect 24811 3556 26148 3584
rect 24811 3553 24823 3556
rect 24765 3547 24823 3553
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 26970 3544 26976 3596
rect 27028 3584 27034 3596
rect 27249 3587 27307 3593
rect 27249 3584 27261 3587
rect 27028 3556 27261 3584
rect 27028 3544 27034 3556
rect 27249 3553 27261 3556
rect 27295 3553 27307 3587
rect 27356 3584 27384 3624
rect 27525 3587 27583 3593
rect 27525 3584 27537 3587
rect 27356 3556 27537 3584
rect 27249 3547 27307 3553
rect 27525 3553 27537 3556
rect 27571 3553 27583 3587
rect 27525 3547 27583 3553
rect 20993 3519 21051 3525
rect 20993 3516 21005 3519
rect 20364 3488 21005 3516
rect 18564 3476 18570 3488
rect 20993 3485 21005 3488
rect 21039 3485 21051 3519
rect 21634 3516 21640 3528
rect 21595 3488 21640 3516
rect 20993 3479 21051 3485
rect 21634 3476 21640 3488
rect 21692 3476 21698 3528
rect 23106 3516 23112 3528
rect 23019 3488 23112 3516
rect 23106 3476 23112 3488
rect 23164 3516 23170 3528
rect 23382 3516 23388 3528
rect 23164 3488 23388 3516
rect 23164 3476 23170 3488
rect 23382 3476 23388 3488
rect 23440 3476 23446 3528
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3516 23903 3519
rect 24670 3516 24676 3528
rect 23891 3488 24676 3516
rect 23891 3485 23903 3488
rect 23845 3479 23903 3485
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 24949 3519 25007 3525
rect 24949 3485 24961 3519
rect 24995 3516 25007 3519
rect 26050 3516 26056 3528
rect 24995 3488 26056 3516
rect 24995 3485 25007 3488
rect 24949 3479 25007 3485
rect 26050 3476 26056 3488
rect 26108 3476 26114 3528
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 26789 3519 26847 3525
rect 26789 3516 26801 3519
rect 26752 3488 26801 3516
rect 26752 3476 26758 3488
rect 26789 3485 26801 3488
rect 26835 3485 26847 3519
rect 26789 3479 26847 3485
rect 28994 3476 29000 3528
rect 29052 3516 29058 3528
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 29052 3488 29561 3516
rect 29052 3476 29058 3488
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 29656 3516 29684 3692
rect 30926 3680 30932 3692
rect 30984 3680 30990 3732
rect 35434 3720 35440 3732
rect 35395 3692 35440 3720
rect 35434 3680 35440 3692
rect 35492 3680 35498 3732
rect 39206 3680 39212 3732
rect 39264 3720 39270 3732
rect 40037 3723 40095 3729
rect 39264 3692 39988 3720
rect 39264 3680 39270 3692
rect 35158 3652 35164 3664
rect 30576 3624 35164 3652
rect 30374 3584 30380 3596
rect 30335 3556 30380 3584
rect 30374 3544 30380 3556
rect 30432 3544 30438 3596
rect 30576 3525 30604 3624
rect 35158 3612 35164 3624
rect 35216 3612 35222 3664
rect 39960 3652 39988 3692
rect 40037 3689 40049 3723
rect 40083 3720 40095 3723
rect 40126 3720 40132 3732
rect 40083 3692 40132 3720
rect 40083 3689 40095 3692
rect 40037 3683 40095 3689
rect 40126 3680 40132 3692
rect 40184 3680 40190 3732
rect 40218 3680 40224 3732
rect 40276 3720 40282 3732
rect 41141 3723 41199 3729
rect 41141 3720 41153 3723
rect 40276 3692 41153 3720
rect 40276 3680 40282 3692
rect 41141 3689 41153 3692
rect 41187 3689 41199 3723
rect 41141 3683 41199 3689
rect 42242 3680 42248 3732
rect 42300 3720 42306 3732
rect 43901 3723 43959 3729
rect 43901 3720 43913 3723
rect 42300 3692 43913 3720
rect 42300 3680 42306 3692
rect 43901 3689 43913 3692
rect 43947 3689 43959 3723
rect 45738 3720 45744 3732
rect 45699 3692 45744 3720
rect 43901 3683 43959 3689
rect 45738 3680 45744 3692
rect 45796 3680 45802 3732
rect 46937 3723 46995 3729
rect 46937 3689 46949 3723
rect 46983 3720 46995 3723
rect 47026 3720 47032 3732
rect 46983 3692 47032 3720
rect 46983 3689 46995 3692
rect 46937 3683 46995 3689
rect 47026 3680 47032 3692
rect 47084 3680 47090 3732
rect 48038 3680 48044 3732
rect 48096 3720 48102 3732
rect 51629 3723 51687 3729
rect 51629 3720 51641 3723
rect 48096 3692 51641 3720
rect 48096 3680 48102 3692
rect 51629 3689 51641 3692
rect 51675 3689 51687 3723
rect 51629 3683 51687 3689
rect 51736 3692 53604 3720
rect 43441 3655 43499 3661
rect 39960 3624 41920 3652
rect 31202 3544 31208 3596
rect 31260 3584 31266 3596
rect 35342 3584 35348 3596
rect 31260 3556 35348 3584
rect 31260 3544 31266 3556
rect 35342 3544 35348 3556
rect 35400 3544 35406 3596
rect 35986 3584 35992 3596
rect 35947 3556 35992 3584
rect 35986 3544 35992 3556
rect 36044 3544 36050 3596
rect 36906 3544 36912 3596
rect 36964 3584 36970 3596
rect 37737 3587 37795 3593
rect 37737 3584 37749 3587
rect 36964 3556 37749 3584
rect 36964 3544 36970 3556
rect 37737 3553 37749 3556
rect 37783 3553 37795 3587
rect 38654 3584 38660 3596
rect 38615 3556 38660 3584
rect 37737 3547 37795 3553
rect 38654 3544 38660 3556
rect 38712 3544 38718 3596
rect 41598 3584 41604 3596
rect 38948 3556 41604 3584
rect 30561 3519 30619 3525
rect 30561 3516 30573 3519
rect 29656 3488 30573 3516
rect 29549 3479 29607 3485
rect 30561 3485 30573 3488
rect 30607 3485 30619 3519
rect 30561 3479 30619 3485
rect 31389 3519 31447 3525
rect 31389 3485 31401 3519
rect 31435 3516 31447 3519
rect 31570 3516 31576 3528
rect 31435 3488 31576 3516
rect 31435 3485 31447 3488
rect 31389 3479 31447 3485
rect 31570 3476 31576 3488
rect 31628 3476 31634 3528
rect 32309 3519 32367 3525
rect 32309 3485 32321 3519
rect 32355 3485 32367 3519
rect 32309 3479 32367 3485
rect 16408 3420 17908 3448
rect 15933 3411 15991 3417
rect 18138 3408 18144 3460
rect 18196 3448 18202 3460
rect 18233 3451 18291 3457
rect 18233 3448 18245 3451
rect 18196 3420 18245 3448
rect 18196 3408 18202 3420
rect 18233 3417 18245 3420
rect 18279 3417 18291 3451
rect 18233 3411 18291 3417
rect 18322 3408 18328 3460
rect 18380 3448 18386 3460
rect 20809 3451 20867 3457
rect 20809 3448 20821 3451
rect 18380 3420 20821 3448
rect 18380 3408 18386 3420
rect 20809 3417 20821 3420
rect 20855 3417 20867 3451
rect 20809 3411 20867 3417
rect 21082 3408 21088 3460
rect 21140 3448 21146 3460
rect 24854 3448 24860 3460
rect 21140 3420 24860 3448
rect 21140 3408 21146 3420
rect 24854 3408 24860 3420
rect 24912 3408 24918 3460
rect 32217 3451 32275 3457
rect 32217 3448 32229 3451
rect 28750 3420 32229 3448
rect 32217 3417 32229 3420
rect 32263 3417 32275 3451
rect 32324 3448 32352 3479
rect 32582 3476 32588 3528
rect 32640 3516 32646 3528
rect 32769 3519 32827 3525
rect 32769 3516 32781 3519
rect 32640 3488 32781 3516
rect 32640 3476 32646 3488
rect 32769 3485 32781 3488
rect 32815 3485 32827 3519
rect 32769 3479 32827 3485
rect 33134 3476 33140 3528
rect 33192 3516 33198 3528
rect 33413 3519 33471 3525
rect 33413 3516 33425 3519
rect 33192 3488 33425 3516
rect 33192 3476 33198 3488
rect 33413 3485 33425 3488
rect 33459 3485 33471 3519
rect 33413 3479 33471 3485
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 33652 3488 33916 3516
rect 33652 3476 33658 3488
rect 33778 3448 33784 3460
rect 32324 3420 33784 3448
rect 32217 3411 32275 3417
rect 33778 3408 33784 3420
rect 33836 3408 33842 3460
rect 33888 3448 33916 3488
rect 33962 3476 33968 3528
rect 34020 3516 34026 3528
rect 34701 3519 34759 3525
rect 34701 3516 34713 3519
rect 34020 3488 34713 3516
rect 34020 3476 34026 3488
rect 34701 3485 34713 3488
rect 34747 3485 34759 3519
rect 34701 3479 34759 3485
rect 36170 3476 36176 3528
rect 36228 3516 36234 3528
rect 37093 3519 37151 3525
rect 37093 3516 37105 3519
rect 36228 3488 37105 3516
rect 36228 3476 36234 3488
rect 37093 3485 37105 3488
rect 37139 3485 37151 3519
rect 37093 3479 37151 3485
rect 38746 3476 38752 3528
rect 38804 3516 38810 3528
rect 38948 3525 38976 3556
rect 41598 3544 41604 3556
rect 41656 3544 41662 3596
rect 38933 3519 38991 3525
rect 38933 3516 38945 3519
rect 38804 3488 38945 3516
rect 38804 3476 38810 3488
rect 38933 3485 38945 3488
rect 38979 3485 38991 3519
rect 39853 3519 39911 3525
rect 39853 3516 39865 3519
rect 38933 3479 38991 3485
rect 39040 3488 39865 3516
rect 36446 3448 36452 3460
rect 33888 3420 36452 3448
rect 36446 3408 36452 3420
rect 36504 3408 36510 3460
rect 38194 3408 38200 3460
rect 38252 3448 38258 3460
rect 38838 3448 38844 3460
rect 38252 3420 38844 3448
rect 38252 3408 38258 3420
rect 38838 3408 38844 3420
rect 38896 3408 38902 3460
rect 17862 3380 17868 3392
rect 13464 3352 17868 3380
rect 13081 3343 13139 3349
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 19794 3340 19800 3392
rect 19852 3380 19858 3392
rect 19889 3383 19947 3389
rect 19889 3380 19901 3383
rect 19852 3352 19901 3380
rect 19852 3340 19858 3352
rect 19889 3349 19901 3352
rect 19935 3349 19947 3383
rect 19889 3343 19947 3349
rect 19978 3340 19984 3392
rect 20036 3380 20042 3392
rect 20036 3352 20081 3380
rect 20036 3340 20042 3352
rect 21726 3340 21732 3392
rect 21784 3380 21790 3392
rect 21821 3383 21879 3389
rect 21821 3380 21833 3383
rect 21784 3352 21833 3380
rect 21784 3340 21790 3352
rect 21821 3349 21833 3352
rect 21867 3349 21879 3383
rect 21821 3343 21879 3349
rect 22925 3383 22983 3389
rect 22925 3349 22937 3383
rect 22971 3380 22983 3383
rect 23566 3380 23572 3392
rect 22971 3352 23572 3380
rect 22971 3349 22983 3352
rect 22925 3343 22983 3349
rect 23566 3340 23572 3352
rect 23624 3340 23630 3392
rect 23661 3383 23719 3389
rect 23661 3349 23673 3383
rect 23707 3380 23719 3383
rect 24302 3380 24308 3392
rect 23707 3352 24308 3380
rect 23707 3349 23719 3352
rect 23661 3343 23719 3349
rect 24302 3340 24308 3352
rect 24360 3340 24366 3392
rect 25682 3340 25688 3392
rect 25740 3380 25746 3392
rect 25869 3383 25927 3389
rect 25869 3380 25881 3383
rect 25740 3352 25881 3380
rect 25740 3340 25746 3352
rect 25869 3349 25881 3352
rect 25915 3349 25927 3383
rect 25869 3343 25927 3349
rect 26234 3340 26240 3392
rect 26292 3380 26298 3392
rect 26605 3383 26663 3389
rect 26605 3380 26617 3383
rect 26292 3352 26617 3380
rect 26292 3340 26298 3352
rect 26605 3349 26617 3352
rect 26651 3349 26663 3383
rect 26605 3343 26663 3349
rect 28997 3383 29055 3389
rect 28997 3349 29009 3383
rect 29043 3380 29055 3383
rect 29086 3380 29092 3392
rect 29043 3352 29092 3380
rect 29043 3349 29055 3352
rect 28997 3343 29055 3349
rect 29086 3340 29092 3352
rect 29144 3340 29150 3392
rect 30466 3380 30472 3392
rect 30427 3352 30472 3380
rect 30466 3340 30472 3352
rect 30524 3340 30530 3392
rect 31573 3383 31631 3389
rect 31573 3349 31585 3383
rect 31619 3380 31631 3383
rect 33870 3380 33876 3392
rect 31619 3352 33876 3380
rect 31619 3349 31631 3352
rect 31573 3343 31631 3349
rect 33870 3340 33876 3352
rect 33928 3340 33934 3392
rect 34054 3380 34060 3392
rect 34015 3352 34060 3380
rect 34054 3340 34060 3352
rect 34112 3340 34118 3392
rect 36078 3340 36084 3392
rect 36136 3380 36142 3392
rect 36173 3383 36231 3389
rect 36173 3380 36185 3383
rect 36136 3352 36185 3380
rect 36136 3340 36142 3352
rect 36173 3349 36185 3352
rect 36219 3349 36231 3383
rect 36173 3343 36231 3349
rect 36262 3340 36268 3392
rect 36320 3380 36326 3392
rect 36633 3383 36691 3389
rect 36320 3352 36365 3380
rect 36320 3340 36326 3352
rect 36633 3349 36645 3383
rect 36679 3380 36691 3383
rect 39040 3380 39068 3488
rect 39853 3485 39865 3488
rect 39899 3485 39911 3519
rect 39853 3479 39911 3485
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40497 3519 40555 3525
rect 40497 3516 40509 3519
rect 40000 3488 40509 3516
rect 40000 3476 40006 3488
rect 40497 3485 40509 3488
rect 40543 3485 40555 3519
rect 41892 3516 41920 3624
rect 43441 3621 43453 3655
rect 43487 3652 43499 3655
rect 44266 3652 44272 3664
rect 43487 3624 44272 3652
rect 43487 3621 43499 3624
rect 43441 3615 43499 3621
rect 44266 3612 44272 3624
rect 44324 3612 44330 3664
rect 50154 3652 50160 3664
rect 50115 3624 50160 3652
rect 50154 3612 50160 3624
rect 50212 3612 50218 3664
rect 51166 3612 51172 3664
rect 51224 3652 51230 3664
rect 51736 3652 51764 3692
rect 51224 3624 51764 3652
rect 53576 3652 53604 3692
rect 55214 3680 55220 3732
rect 55272 3720 55278 3732
rect 56042 3720 56048 3732
rect 55272 3692 56048 3720
rect 55272 3680 55278 3692
rect 56042 3680 56048 3692
rect 56100 3680 56106 3732
rect 55309 3655 55367 3661
rect 53576 3624 55214 3652
rect 51224 3612 51230 3624
rect 44634 3544 44640 3596
rect 44692 3584 44698 3596
rect 45186 3584 45192 3596
rect 44692 3556 45192 3584
rect 44692 3544 44698 3556
rect 45186 3544 45192 3556
rect 45244 3544 45250 3596
rect 45922 3544 45928 3596
rect 45980 3584 45986 3596
rect 49053 3587 49111 3593
rect 49053 3584 49065 3587
rect 45980 3556 49065 3584
rect 45980 3544 45986 3556
rect 49053 3553 49065 3556
rect 49099 3553 49111 3587
rect 49326 3584 49332 3596
rect 49287 3556 49332 3584
rect 49053 3547 49111 3553
rect 49326 3544 49332 3556
rect 49384 3544 49390 3596
rect 52178 3544 52184 3596
rect 52236 3584 52242 3596
rect 52273 3587 52331 3593
rect 52273 3584 52285 3587
rect 52236 3556 52285 3584
rect 52236 3544 52242 3556
rect 52273 3553 52285 3556
rect 52319 3553 52331 3587
rect 52546 3584 52552 3596
rect 52507 3556 52552 3584
rect 52273 3547 52331 3553
rect 52546 3544 52552 3556
rect 52604 3544 52610 3596
rect 52638 3544 52644 3596
rect 52696 3584 52702 3596
rect 52696 3556 54708 3584
rect 52696 3544 52702 3556
rect 42426 3516 42432 3528
rect 41892 3488 42432 3516
rect 40497 3479 40555 3485
rect 42426 3476 42432 3488
rect 42484 3476 42490 3528
rect 42521 3519 42579 3525
rect 42521 3485 42533 3519
rect 42567 3516 42579 3519
rect 42610 3516 42616 3528
rect 42567 3488 42616 3516
rect 42567 3485 42579 3488
rect 42521 3479 42579 3485
rect 42610 3476 42616 3488
rect 42668 3476 42674 3528
rect 42797 3519 42855 3525
rect 42797 3485 42809 3519
rect 42843 3516 42855 3519
rect 42886 3516 42892 3528
rect 42843 3488 42892 3516
rect 42843 3485 42855 3488
rect 42797 3479 42855 3485
rect 42886 3476 42892 3488
rect 42944 3476 42950 3528
rect 43257 3519 43315 3525
rect 43257 3485 43269 3519
rect 43303 3485 43315 3519
rect 43257 3479 43315 3485
rect 43272 3448 43300 3479
rect 45370 3476 45376 3528
rect 45428 3476 45434 3528
rect 46566 3516 46572 3528
rect 46527 3488 46572 3516
rect 46566 3476 46572 3488
rect 46624 3476 46630 3528
rect 46658 3476 46664 3528
rect 46716 3516 46722 3528
rect 46716 3488 47978 3516
rect 46716 3476 46722 3488
rect 49418 3476 49424 3528
rect 49476 3516 49482 3528
rect 50706 3516 50712 3528
rect 49476 3488 50712 3516
rect 49476 3476 49482 3488
rect 50706 3476 50712 3488
rect 50764 3476 50770 3528
rect 50890 3516 50896 3528
rect 50851 3488 50896 3516
rect 50890 3476 50896 3488
rect 50948 3476 50954 3528
rect 51166 3516 51172 3528
rect 51127 3488 51172 3516
rect 51166 3476 51172 3488
rect 51224 3476 51230 3528
rect 39316 3420 40540 3448
rect 39316 3389 39344 3420
rect 36679 3352 39068 3380
rect 39301 3383 39359 3389
rect 36679 3349 36691 3352
rect 36633 3343 36691 3349
rect 39301 3349 39313 3383
rect 39347 3349 39359 3383
rect 39301 3343 39359 3349
rect 39482 3340 39488 3392
rect 39540 3380 39546 3392
rect 40218 3380 40224 3392
rect 39540 3352 40224 3380
rect 39540 3340 39546 3352
rect 40218 3340 40224 3352
rect 40276 3340 40282 3392
rect 40512 3380 40540 3420
rect 41386 3420 43300 3448
rect 45281 3451 45339 3457
rect 41386 3380 41414 3420
rect 45281 3417 45293 3451
rect 45327 3448 45339 3451
rect 45388 3448 45416 3476
rect 47026 3448 47032 3460
rect 45327 3420 47032 3448
rect 45327 3417 45339 3420
rect 45281 3411 45339 3417
rect 47026 3408 47032 3420
rect 47084 3408 47090 3460
rect 49326 3408 49332 3460
rect 49384 3448 49390 3460
rect 52196 3448 52224 3544
rect 54573 3519 54631 3525
rect 54573 3516 54585 3519
rect 53852 3488 54585 3516
rect 49384 3420 52224 3448
rect 49384 3408 49390 3420
rect 52822 3408 52828 3460
rect 52880 3448 52886 3460
rect 52880 3420 53038 3448
rect 52880 3408 52886 3420
rect 41782 3380 41788 3392
rect 40512 3352 41414 3380
rect 41743 3352 41788 3380
rect 41782 3340 41788 3352
rect 41840 3340 41846 3392
rect 45373 3383 45431 3389
rect 45373 3349 45385 3383
rect 45419 3380 45431 3383
rect 45462 3380 45468 3392
rect 45419 3352 45468 3380
rect 45419 3349 45431 3352
rect 45373 3343 45431 3349
rect 45462 3340 45468 3352
rect 45520 3340 45526 3392
rect 46934 3380 46940 3392
rect 46895 3352 46940 3380
rect 46934 3340 46940 3352
rect 46992 3340 46998 3392
rect 47118 3380 47124 3392
rect 47079 3352 47124 3380
rect 47118 3340 47124 3352
rect 47176 3340 47182 3392
rect 47578 3380 47584 3392
rect 47539 3352 47584 3380
rect 47578 3340 47584 3352
rect 47636 3340 47642 3392
rect 48866 3340 48872 3392
rect 48924 3380 48930 3392
rect 53852 3380 53880 3488
rect 54573 3485 54585 3488
rect 54619 3485 54631 3519
rect 54573 3479 54631 3485
rect 54680 3448 54708 3556
rect 55186 3516 55214 3624
rect 55309 3621 55321 3655
rect 55355 3621 55367 3655
rect 55309 3615 55367 3621
rect 55324 3584 55352 3615
rect 55490 3612 55496 3664
rect 55548 3652 55554 3664
rect 57793 3655 57851 3661
rect 57793 3652 57805 3655
rect 55548 3624 57805 3652
rect 55548 3612 55554 3624
rect 57793 3621 57805 3624
rect 57839 3621 57851 3655
rect 57793 3615 57851 3621
rect 55398 3584 55404 3596
rect 55324 3556 55404 3584
rect 55398 3544 55404 3556
rect 55456 3544 55462 3596
rect 55858 3584 55864 3596
rect 55819 3556 55864 3584
rect 55858 3544 55864 3556
rect 55916 3584 55922 3596
rect 56226 3584 56232 3596
rect 55916 3556 56232 3584
rect 55916 3544 55922 3556
rect 56226 3544 56232 3556
rect 56284 3544 56290 3596
rect 56505 3519 56563 3525
rect 56505 3516 56517 3519
rect 55186 3488 56517 3516
rect 56505 3485 56517 3488
rect 56551 3485 56563 3519
rect 56505 3479 56563 3485
rect 57333 3519 57391 3525
rect 57333 3485 57345 3519
rect 57379 3485 57391 3519
rect 57333 3479 57391 3485
rect 57348 3448 57376 3479
rect 57422 3476 57428 3528
rect 57480 3516 57486 3528
rect 57977 3519 58035 3525
rect 57977 3516 57989 3519
rect 57480 3488 57989 3516
rect 57480 3476 57486 3488
rect 57977 3485 57989 3488
rect 58023 3485 58035 3519
rect 57977 3479 58035 3485
rect 54680 3420 57376 3448
rect 48924 3352 53880 3380
rect 48924 3340 48930 3352
rect 54018 3340 54024 3392
rect 54076 3380 54082 3392
rect 55306 3380 55312 3392
rect 54076 3352 55312 3380
rect 54076 3340 54082 3352
rect 55306 3340 55312 3352
rect 55364 3340 55370 3392
rect 55674 3380 55680 3392
rect 55635 3352 55680 3380
rect 55674 3340 55680 3352
rect 55732 3340 55738 3392
rect 55766 3340 55772 3392
rect 55824 3380 55830 3392
rect 55824 3352 55869 3380
rect 55824 3340 55830 3352
rect 55950 3340 55956 3392
rect 56008 3380 56014 3392
rect 57149 3383 57207 3389
rect 57149 3380 57161 3383
rect 56008 3352 57161 3380
rect 56008 3340 56014 3352
rect 57149 3349 57161 3352
rect 57195 3349 57207 3383
rect 57149 3343 57207 3349
rect 1104 3290 58880 3312
rect 1104 3238 15398 3290
rect 15450 3238 15462 3290
rect 15514 3238 15526 3290
rect 15578 3238 15590 3290
rect 15642 3238 15654 3290
rect 15706 3238 29846 3290
rect 29898 3238 29910 3290
rect 29962 3238 29974 3290
rect 30026 3238 30038 3290
rect 30090 3238 30102 3290
rect 30154 3238 44294 3290
rect 44346 3238 44358 3290
rect 44410 3238 44422 3290
rect 44474 3238 44486 3290
rect 44538 3238 44550 3290
rect 44602 3238 58880 3290
rect 1104 3216 58880 3238
rect 2961 3179 3019 3185
rect 2961 3145 2973 3179
rect 3007 3176 3019 3179
rect 3007 3148 6776 3176
rect 3007 3145 3019 3148
rect 2961 3139 3019 3145
rect 3436 3080 5488 3108
rect 3436 3049 3464 3080
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3040 1915 3043
rect 3421 3043 3479 3049
rect 3421 3040 3433 3043
rect 1903 3012 3433 3040
rect 1903 3009 1915 3012
rect 1857 3003 1915 3009
rect 3421 3009 3433 3012
rect 3467 3009 3479 3043
rect 4341 3043 4399 3049
rect 3421 3003 3479 3009
rect 3620 3012 4292 3040
rect 3620 2913 3648 3012
rect 3605 2907 3663 2913
rect 3605 2873 3617 2907
rect 3651 2873 3663 2907
rect 4264 2904 4292 3012
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4430 3040 4436 3052
rect 4387 3012 4436 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 4430 3000 4436 3012
rect 4488 3000 4494 3052
rect 4614 3040 4620 3052
rect 4575 3012 4620 3040
rect 4614 3000 4620 3012
rect 4672 3040 4678 3052
rect 5261 3043 5319 3049
rect 5261 3040 5273 3043
rect 4672 3012 5273 3040
rect 4672 3000 4678 3012
rect 5261 3009 5273 3012
rect 5307 3009 5319 3043
rect 5261 3003 5319 3009
rect 4525 2975 4583 2981
rect 4525 2941 4537 2975
rect 4571 2972 4583 2975
rect 5074 2972 5080 2984
rect 4571 2944 5080 2972
rect 4571 2941 4583 2944
rect 4525 2935 4583 2941
rect 5074 2932 5080 2944
rect 5132 2972 5138 2984
rect 5169 2975 5227 2981
rect 5169 2972 5181 2975
rect 5132 2944 5181 2972
rect 5132 2932 5138 2944
rect 5169 2941 5181 2944
rect 5215 2941 5227 2975
rect 5169 2935 5227 2941
rect 4982 2904 4988 2916
rect 4264 2876 4988 2904
rect 3605 2867 3663 2873
rect 4982 2864 4988 2876
rect 5040 2864 5046 2916
rect 5276 2904 5304 3003
rect 5460 2972 5488 3080
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 6748 3108 6776 3148
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 6880 3148 6925 3176
rect 6880 3136 6886 3148
rect 7282 3136 7288 3188
rect 7340 3176 7346 3188
rect 10134 3176 10140 3188
rect 7340 3148 10140 3176
rect 7340 3136 7346 3148
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 11606 3176 11612 3188
rect 11567 3148 11612 3176
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 13354 3176 13360 3188
rect 12176 3148 13360 3176
rect 7374 3108 7380 3120
rect 5592 3080 6500 3108
rect 6748 3080 7380 3108
rect 5592 3068 5598 3080
rect 5626 3000 5632 3052
rect 5684 3040 5690 3052
rect 6472 3049 6500 3080
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 7742 3068 7748 3120
rect 7800 3108 7806 3120
rect 11698 3108 11704 3120
rect 7800 3080 11704 3108
rect 7800 3068 7806 3080
rect 11698 3068 11704 3080
rect 11756 3068 11762 3120
rect 6457 3043 6515 3049
rect 5684 3012 5729 3040
rect 5684 3000 5690 3012
rect 6457 3009 6469 3043
rect 6503 3009 6515 3043
rect 6638 3040 6644 3052
rect 6599 3012 6644 3040
rect 6457 3003 6515 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 7190 3040 7196 3052
rect 7055 3012 7196 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 7190 3000 7196 3012
rect 7248 3000 7254 3052
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3009 7895 3043
rect 8754 3040 8760 3052
rect 8715 3012 8760 3040
rect 7837 3003 7895 3009
rect 7558 2972 7564 2984
rect 5460 2944 7564 2972
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 7852 2972 7880 3003
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3040 9735 3043
rect 12176 3040 12204 3148
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 13449 3179 13507 3185
rect 13449 3145 13461 3179
rect 13495 3176 13507 3179
rect 13538 3176 13544 3188
rect 13495 3148 13544 3176
rect 13495 3145 13507 3148
rect 13449 3139 13507 3145
rect 13538 3136 13544 3148
rect 13596 3136 13602 3188
rect 13722 3136 13728 3188
rect 13780 3176 13786 3188
rect 14737 3179 14795 3185
rect 14737 3176 14749 3179
rect 13780 3148 14749 3176
rect 13780 3136 13786 3148
rect 14737 3145 14749 3148
rect 14783 3145 14795 3179
rect 15654 3176 15660 3188
rect 14737 3139 14795 3145
rect 15120 3148 15660 3176
rect 15120 3108 15148 3148
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 15838 3136 15844 3188
rect 15896 3176 15902 3188
rect 16390 3176 16396 3188
rect 15896 3148 16396 3176
rect 15896 3136 15902 3148
rect 16390 3136 16396 3148
rect 16448 3136 16454 3188
rect 17681 3179 17739 3185
rect 17681 3145 17693 3179
rect 17727 3145 17739 3179
rect 17681 3139 17739 3145
rect 12268 3080 15148 3108
rect 12268 3049 12296 3080
rect 15194 3068 15200 3120
rect 15252 3108 15258 3120
rect 17696 3108 17724 3139
rect 18046 3136 18052 3188
rect 18104 3176 18110 3188
rect 18506 3176 18512 3188
rect 18104 3148 18512 3176
rect 18104 3136 18110 3148
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 19794 3136 19800 3188
rect 19852 3176 19858 3188
rect 20809 3179 20867 3185
rect 20809 3176 20821 3179
rect 19852 3148 20821 3176
rect 19852 3136 19858 3148
rect 20809 3145 20821 3148
rect 20855 3145 20867 3179
rect 20809 3139 20867 3145
rect 23845 3179 23903 3185
rect 23845 3145 23857 3179
rect 23891 3176 23903 3179
rect 24118 3176 24124 3188
rect 23891 3148 24124 3176
rect 23891 3145 23903 3148
rect 23845 3139 23903 3145
rect 24118 3136 24124 3148
rect 24176 3136 24182 3188
rect 24670 3136 24676 3188
rect 24728 3176 24734 3188
rect 31202 3176 31208 3188
rect 24728 3148 31208 3176
rect 24728 3136 24734 3148
rect 31202 3136 31208 3148
rect 31260 3136 31266 3188
rect 31570 3176 31576 3188
rect 31531 3148 31576 3176
rect 31570 3136 31576 3148
rect 31628 3136 31634 3188
rect 32306 3136 32312 3188
rect 32364 3176 32370 3188
rect 34790 3176 34796 3188
rect 32364 3148 34796 3176
rect 32364 3136 32370 3148
rect 34790 3136 34796 3148
rect 34848 3136 34854 3188
rect 35250 3136 35256 3188
rect 35308 3176 35314 3188
rect 35308 3148 37964 3176
rect 35308 3136 35314 3148
rect 19674 3111 19732 3117
rect 19674 3108 19686 3111
rect 15252 3080 15976 3108
rect 17696 3080 19686 3108
rect 15252 3068 15258 3080
rect 9723 3012 12204 3040
rect 12253 3043 12311 3049
rect 9723 3009 9735 3012
rect 9677 3003 9735 3009
rect 12253 3009 12265 3043
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 12526 3000 12532 3052
rect 12584 3040 12590 3052
rect 12710 3040 12716 3052
rect 12584 3012 12716 3040
rect 12584 3000 12590 3012
rect 12710 3000 12716 3012
rect 12768 3040 12774 3052
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 12768 3012 12817 3040
rect 12768 3000 12774 3012
rect 12805 3009 12817 3012
rect 12851 3009 12863 3043
rect 12805 3003 12863 3009
rect 12894 3000 12900 3052
rect 12952 3040 12958 3052
rect 13262 3040 13268 3052
rect 12952 3012 12997 3040
rect 13223 3012 13268 3040
rect 12952 3000 12958 3012
rect 13262 3000 13268 3012
rect 13320 3000 13326 3052
rect 13354 3000 13360 3052
rect 13412 3040 13418 3052
rect 13538 3040 13544 3052
rect 13412 3012 13544 3040
rect 13412 3000 13418 3012
rect 13538 3000 13544 3012
rect 13596 3000 13602 3052
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14369 3043 14427 3049
rect 14369 3040 14381 3043
rect 14056 3012 14381 3040
rect 14056 3000 14062 3012
rect 14369 3009 14381 3012
rect 14415 3009 14427 3043
rect 14369 3003 14427 3009
rect 15565 3043 15623 3049
rect 15565 3009 15577 3043
rect 15611 3040 15623 3043
rect 15746 3040 15752 3052
rect 15611 3012 15752 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 15948 3049 15976 3080
rect 19674 3077 19686 3080
rect 19720 3077 19732 3111
rect 25133 3111 25191 3117
rect 19674 3071 19732 3077
rect 22204 3080 24716 3108
rect 15933 3043 15991 3049
rect 15933 3009 15945 3043
rect 15979 3009 15991 3043
rect 15933 3003 15991 3009
rect 16025 3043 16083 3049
rect 16025 3009 16037 3043
rect 16071 3040 16083 3043
rect 16298 3040 16304 3052
rect 16071 3012 16304 3040
rect 16071 3009 16083 3012
rect 16025 3003 16083 3009
rect 16298 3000 16304 3012
rect 16356 3000 16362 3052
rect 17497 3043 17555 3049
rect 17497 3009 17509 3043
rect 17543 3040 17555 3043
rect 18322 3040 18328 3052
rect 17543 3012 18328 3040
rect 17543 3009 17555 3012
rect 17497 3003 17555 3009
rect 18322 3000 18328 3012
rect 18380 3000 18386 3052
rect 19242 3000 19248 3052
rect 19300 3040 19306 3052
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 19300 3012 19441 3040
rect 19300 3000 19306 3012
rect 19429 3009 19441 3012
rect 19475 3009 19487 3043
rect 20438 3040 20444 3052
rect 19429 3003 19487 3009
rect 19536 3012 20444 3040
rect 8294 2972 8300 2984
rect 7852 2944 8300 2972
rect 8294 2932 8300 2944
rect 8352 2972 8358 2984
rect 9398 2972 9404 2984
rect 8352 2944 9404 2972
rect 8352 2932 8358 2944
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 10226 2932 10232 2984
rect 10284 2972 10290 2984
rect 12342 2972 12348 2984
rect 10284 2944 12348 2972
rect 10284 2932 10290 2944
rect 12342 2932 12348 2944
rect 12400 2932 12406 2984
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 13630 2972 13636 2984
rect 13044 2944 13636 2972
rect 13044 2932 13050 2944
rect 13630 2932 13636 2944
rect 13688 2932 13694 2984
rect 13814 2932 13820 2984
rect 13872 2972 13878 2984
rect 14461 2975 14519 2981
rect 14461 2972 14473 2975
rect 13872 2944 14473 2972
rect 13872 2932 13878 2944
rect 14461 2941 14473 2944
rect 14507 2972 14519 2975
rect 14550 2972 14556 2984
rect 14507 2944 14556 2972
rect 14507 2941 14519 2944
rect 14461 2935 14519 2941
rect 14550 2932 14556 2944
rect 14608 2932 14614 2984
rect 15286 2932 15292 2984
rect 15344 2972 15350 2984
rect 16390 2972 16396 2984
rect 15344 2944 16396 2972
rect 15344 2932 15350 2944
rect 16390 2932 16396 2944
rect 16448 2932 16454 2984
rect 19536 2972 19564 3012
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 22204 3049 22232 3080
rect 24688 3052 24716 3080
rect 25133 3077 25145 3111
rect 25179 3108 25191 3111
rect 28626 3108 28632 3120
rect 25179 3080 28632 3108
rect 25179 3077 25191 3080
rect 25133 3071 25191 3077
rect 28626 3068 28632 3080
rect 28684 3068 28690 3120
rect 30377 3111 30435 3117
rect 30377 3077 30389 3111
rect 30423 3108 30435 3111
rect 31386 3108 31392 3120
rect 30423 3080 31392 3108
rect 30423 3077 30435 3080
rect 30377 3071 30435 3077
rect 31386 3068 31392 3080
rect 31444 3068 31450 3120
rect 33870 3108 33876 3120
rect 33831 3080 33876 3108
rect 33870 3068 33876 3080
rect 33928 3068 33934 3120
rect 35098 3080 37504 3108
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3009 22247 3043
rect 22189 3003 22247 3009
rect 22925 3043 22983 3049
rect 22925 3009 22937 3043
rect 22971 3040 22983 3043
rect 22971 3012 24532 3040
rect 22971 3009 22983 3012
rect 22925 3003 22983 3009
rect 24504 2984 24532 3012
rect 24670 3000 24676 3052
rect 24728 3000 24734 3052
rect 24854 3000 24860 3052
rect 24912 3040 24918 3052
rect 26053 3043 26111 3049
rect 26053 3040 26065 3043
rect 24912 3012 26065 3040
rect 24912 3000 24918 3012
rect 26053 3009 26065 3012
rect 26099 3009 26111 3043
rect 26053 3003 26111 3009
rect 26602 3000 26608 3052
rect 26660 3040 26666 3052
rect 27249 3043 27307 3049
rect 27249 3040 27261 3043
rect 26660 3012 27261 3040
rect 26660 3000 26666 3012
rect 27249 3009 27261 3012
rect 27295 3040 27307 3043
rect 27338 3040 27344 3052
rect 27295 3012 27344 3040
rect 27295 3009 27307 3012
rect 27249 3003 27307 3009
rect 27338 3000 27344 3012
rect 27396 3000 27402 3052
rect 29086 3000 29092 3052
rect 29144 3040 29150 3052
rect 31113 3043 31171 3049
rect 31113 3040 31125 3043
rect 29144 3012 31125 3040
rect 29144 3000 29150 3012
rect 31113 3009 31125 3012
rect 31159 3009 31171 3043
rect 32766 3040 32772 3052
rect 31113 3003 31171 3009
rect 31220 3012 32772 3040
rect 18340 2944 19564 2972
rect 5534 2904 5540 2916
rect 5276 2876 5540 2904
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 5644 2876 6408 2904
rect 2409 2839 2467 2845
rect 2409 2805 2421 2839
rect 2455 2836 2467 2839
rect 2774 2836 2780 2848
rect 2455 2808 2780 2836
rect 2455 2805 2467 2808
rect 2409 2799 2467 2805
rect 2774 2796 2780 2808
rect 2832 2836 2838 2848
rect 2958 2836 2964 2848
rect 2832 2808 2964 2836
rect 2832 2796 2838 2808
rect 2958 2796 2964 2808
rect 3016 2796 3022 2848
rect 4062 2796 4068 2848
rect 4120 2836 4126 2848
rect 4157 2839 4215 2845
rect 4157 2836 4169 2839
rect 4120 2808 4169 2836
rect 4120 2796 4126 2808
rect 4157 2805 4169 2808
rect 4203 2805 4215 2839
rect 4338 2836 4344 2848
rect 4299 2808 4344 2836
rect 4157 2799 4215 2805
rect 4338 2796 4344 2808
rect 4396 2796 4402 2848
rect 4430 2796 4436 2848
rect 4488 2836 4494 2848
rect 5258 2836 5264 2848
rect 4488 2808 5264 2836
rect 4488 2796 4494 2808
rect 5258 2796 5264 2808
rect 5316 2796 5322 2848
rect 5350 2796 5356 2848
rect 5408 2836 5414 2848
rect 5644 2845 5672 2876
rect 6380 2848 6408 2876
rect 8938 2864 8944 2916
rect 8996 2904 9002 2916
rect 9214 2904 9220 2916
rect 8996 2876 9220 2904
rect 8996 2864 9002 2876
rect 9214 2864 9220 2876
rect 9272 2904 9278 2916
rect 10965 2907 11023 2913
rect 9272 2876 10916 2904
rect 9272 2864 9278 2876
rect 5629 2839 5687 2845
rect 5629 2836 5641 2839
rect 5408 2808 5641 2836
rect 5408 2796 5414 2808
rect 5629 2805 5641 2808
rect 5675 2805 5687 2839
rect 5810 2836 5816 2848
rect 5771 2808 5816 2836
rect 5629 2799 5687 2805
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 6420 2808 6561 2836
rect 6420 2796 6426 2808
rect 6549 2805 6561 2808
rect 6595 2805 6607 2839
rect 6549 2799 6607 2805
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 7653 2839 7711 2845
rect 7653 2836 7665 2839
rect 7524 2808 7665 2836
rect 7524 2796 7530 2808
rect 7653 2805 7665 2808
rect 7699 2805 7711 2839
rect 8570 2836 8576 2848
rect 8531 2808 8576 2836
rect 7653 2799 7711 2805
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 10321 2839 10379 2845
rect 10321 2805 10333 2839
rect 10367 2836 10379 2839
rect 10778 2836 10784 2848
rect 10367 2808 10784 2836
rect 10367 2805 10379 2808
rect 10321 2799 10379 2805
rect 10778 2796 10784 2808
rect 10836 2796 10842 2848
rect 10888 2836 10916 2876
rect 10965 2873 10977 2907
rect 11011 2904 11023 2907
rect 13906 2904 13912 2916
rect 11011 2876 13912 2904
rect 11011 2873 11023 2876
rect 10965 2867 11023 2873
rect 13906 2864 13912 2876
rect 13964 2864 13970 2916
rect 18340 2913 18368 2944
rect 24486 2932 24492 2984
rect 24544 2972 24550 2984
rect 29104 2972 29132 3000
rect 24544 2944 29132 2972
rect 24544 2932 24550 2944
rect 30374 2932 30380 2984
rect 30432 2972 30438 2984
rect 30929 2975 30987 2981
rect 30929 2972 30941 2975
rect 30432 2944 30941 2972
rect 30432 2932 30438 2944
rect 30929 2941 30941 2944
rect 30975 2972 30987 2975
rect 31220 2972 31248 3012
rect 32766 3000 32772 3012
rect 32824 3000 32830 3052
rect 33502 3000 33508 3052
rect 33560 3040 33566 3052
rect 33597 3043 33655 3049
rect 33597 3040 33609 3043
rect 33560 3012 33609 3040
rect 33560 3000 33566 3012
rect 33597 3009 33609 3012
rect 33643 3009 33655 3043
rect 33597 3003 33655 3009
rect 35158 3000 35164 3052
rect 35216 3040 35222 3052
rect 37277 3043 37335 3049
rect 37277 3040 37289 3043
rect 35216 3012 37289 3040
rect 35216 3000 35222 3012
rect 37277 3009 37289 3012
rect 37323 3009 37335 3043
rect 37277 3003 37335 3009
rect 30975 2944 31248 2972
rect 30975 2941 30987 2944
rect 30929 2935 30987 2941
rect 31754 2932 31760 2984
rect 31812 2972 31818 2984
rect 34514 2972 34520 2984
rect 31812 2944 34520 2972
rect 31812 2932 31818 2944
rect 34514 2932 34520 2944
rect 34572 2932 34578 2984
rect 34606 2932 34612 2984
rect 34664 2972 34670 2984
rect 36814 2972 36820 2984
rect 34664 2944 36820 2972
rect 34664 2932 34670 2944
rect 36814 2932 36820 2944
rect 36872 2932 36878 2984
rect 37476 2972 37504 3080
rect 37936 3049 37964 3148
rect 38930 3136 38936 3188
rect 38988 3176 38994 3188
rect 39850 3176 39856 3188
rect 38988 3148 39856 3176
rect 38988 3136 38994 3148
rect 39850 3136 39856 3148
rect 39908 3136 39914 3188
rect 41690 3136 41696 3188
rect 41748 3176 41754 3188
rect 41748 3148 41920 3176
rect 41748 3136 41754 3148
rect 39945 3111 40003 3117
rect 39945 3108 39957 3111
rect 38028 3080 39957 3108
rect 37921 3043 37979 3049
rect 37921 3009 37933 3043
rect 37967 3009 37979 3043
rect 37921 3003 37979 3009
rect 38028 2972 38056 3080
rect 39945 3077 39957 3080
rect 39991 3077 40003 3111
rect 39945 3071 40003 3077
rect 40586 3068 40592 3120
rect 40644 3068 40650 3120
rect 41598 3068 41604 3120
rect 41656 3108 41662 3120
rect 41785 3111 41843 3117
rect 41785 3108 41797 3111
rect 41656 3080 41797 3108
rect 41656 3068 41662 3080
rect 41785 3077 41797 3080
rect 41831 3077 41843 3111
rect 41892 3108 41920 3148
rect 42518 3136 42524 3188
rect 42576 3176 42582 3188
rect 45002 3176 45008 3188
rect 42576 3148 45008 3176
rect 42576 3136 42582 3148
rect 45002 3136 45008 3148
rect 45060 3136 45066 3188
rect 45112 3148 45784 3176
rect 43070 3108 43076 3120
rect 41892 3080 43076 3108
rect 41785 3071 41843 3077
rect 43070 3068 43076 3080
rect 43128 3068 43134 3120
rect 43162 3068 43168 3120
rect 43220 3108 43226 3120
rect 45112 3108 45140 3148
rect 43220 3080 45140 3108
rect 45756 3108 45784 3148
rect 46106 3136 46112 3188
rect 46164 3176 46170 3188
rect 49418 3176 49424 3188
rect 46164 3148 49424 3176
rect 46164 3136 46170 3148
rect 49418 3136 49424 3148
rect 49476 3136 49482 3188
rect 49602 3136 49608 3188
rect 49660 3176 49666 3188
rect 50270 3179 50328 3185
rect 50270 3176 50282 3179
rect 49660 3148 50282 3176
rect 49660 3136 49666 3148
rect 50270 3145 50282 3148
rect 50316 3145 50328 3179
rect 50270 3139 50328 3145
rect 50433 3179 50491 3185
rect 50433 3145 50445 3179
rect 50479 3176 50491 3179
rect 52638 3176 52644 3188
rect 50479 3148 52644 3176
rect 50479 3145 50491 3148
rect 50433 3139 50491 3145
rect 52638 3136 52644 3148
rect 52696 3136 52702 3188
rect 53944 3148 57928 3176
rect 47026 3108 47032 3120
rect 45756 3080 46336 3108
rect 46987 3080 47032 3108
rect 43220 3068 43226 3080
rect 40037 3043 40095 3049
rect 40037 3009 40049 3043
rect 40083 3040 40095 3043
rect 40126 3040 40132 3052
rect 40083 3012 40132 3040
rect 40083 3009 40095 3012
rect 40037 3003 40095 3009
rect 40126 3000 40132 3012
rect 40184 3040 40190 3052
rect 40604 3040 40632 3068
rect 43717 3043 43775 3049
rect 43717 3040 43729 3043
rect 40184 3012 40632 3040
rect 41386 3012 43729 3040
rect 40184 3000 40190 3012
rect 37476 2944 38056 2972
rect 38102 2932 38108 2984
rect 38160 2972 38166 2984
rect 40497 2975 40555 2981
rect 40497 2972 40509 2975
rect 38160 2944 40509 2972
rect 38160 2932 38166 2944
rect 40497 2941 40509 2944
rect 40543 2941 40555 2975
rect 40497 2935 40555 2941
rect 40586 2932 40592 2984
rect 40644 2972 40650 2984
rect 41386 2972 41414 3012
rect 43717 3009 43729 3012
rect 43763 3009 43775 3043
rect 43717 3003 43775 3009
rect 43898 3000 43904 3052
rect 43956 3040 43962 3052
rect 43956 3012 45140 3040
rect 43956 3000 43962 3012
rect 44361 2975 44419 2981
rect 44361 2972 44373 2975
rect 40644 2944 41414 2972
rect 41524 2944 44373 2972
rect 40644 2932 40650 2944
rect 15381 2907 15439 2913
rect 15381 2904 15393 2907
rect 14384 2876 15393 2904
rect 14384 2848 14412 2876
rect 15381 2873 15393 2876
rect 15427 2873 15439 2907
rect 15381 2867 15439 2873
rect 18325 2907 18383 2913
rect 18325 2873 18337 2907
rect 18371 2873 18383 2907
rect 19334 2904 19340 2916
rect 18325 2867 18383 2873
rect 18892 2876 19340 2904
rect 12250 2836 12256 2848
rect 10888 2808 12256 2836
rect 12250 2796 12256 2808
rect 12308 2796 12314 2848
rect 12618 2796 12624 2848
rect 12676 2836 12682 2848
rect 13265 2839 13323 2845
rect 13265 2836 13277 2839
rect 12676 2808 13277 2836
rect 12676 2796 12682 2808
rect 13265 2805 13277 2808
rect 13311 2836 13323 2839
rect 13354 2836 13360 2848
rect 13311 2808 13360 2836
rect 13311 2805 13323 2808
rect 13265 2799 13323 2805
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 14366 2836 14372 2848
rect 14327 2808 14372 2836
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 15562 2836 15568 2848
rect 15523 2808 15568 2836
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 17037 2839 17095 2845
rect 17037 2805 17049 2839
rect 17083 2836 17095 2839
rect 18892 2836 18920 2876
rect 19334 2864 19340 2876
rect 19392 2864 19398 2916
rect 20990 2904 20996 2916
rect 20732 2876 20996 2904
rect 17083 2808 18920 2836
rect 18969 2839 19027 2845
rect 17083 2805 17095 2808
rect 17037 2799 17095 2805
rect 18969 2805 18981 2839
rect 19015 2836 19027 2839
rect 20732 2836 20760 2876
rect 20990 2864 20996 2876
rect 21048 2864 21054 2916
rect 22005 2907 22063 2913
rect 22005 2873 22017 2907
rect 22051 2904 22063 2907
rect 23750 2904 23756 2916
rect 22051 2876 23756 2904
rect 22051 2873 22063 2876
rect 22005 2867 22063 2873
rect 23750 2864 23756 2876
rect 23808 2864 23814 2916
rect 23842 2864 23848 2916
rect 23900 2904 23906 2916
rect 26878 2904 26884 2916
rect 23900 2876 26884 2904
rect 23900 2864 23906 2876
rect 26878 2864 26884 2876
rect 26936 2864 26942 2916
rect 31478 2864 31484 2916
rect 31536 2904 31542 2916
rect 32769 2907 32827 2913
rect 32769 2904 32781 2907
rect 31536 2876 32781 2904
rect 31536 2864 31542 2876
rect 32769 2873 32781 2876
rect 32815 2873 32827 2907
rect 35805 2907 35863 2913
rect 35805 2904 35817 2907
rect 32769 2867 32827 2873
rect 34900 2876 35817 2904
rect 19015 2808 20760 2836
rect 22741 2839 22799 2845
rect 19015 2805 19027 2808
rect 18969 2799 19027 2805
rect 22741 2805 22753 2839
rect 22787 2836 22799 2839
rect 24026 2836 24032 2848
rect 22787 2808 24032 2836
rect 22787 2805 22799 2808
rect 22741 2799 22799 2805
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 25958 2796 25964 2848
rect 26016 2836 26022 2848
rect 26237 2839 26295 2845
rect 26237 2836 26249 2839
rect 26016 2808 26249 2836
rect 26016 2796 26022 2808
rect 26237 2805 26249 2808
rect 26283 2805 26295 2839
rect 26237 2799 26295 2805
rect 26510 2796 26516 2848
rect 26568 2836 26574 2848
rect 27065 2839 27123 2845
rect 27065 2836 27077 2839
rect 26568 2808 27077 2836
rect 26568 2796 26574 2808
rect 27065 2805 27077 2808
rect 27111 2805 27123 2839
rect 27065 2799 27123 2805
rect 28169 2839 28227 2845
rect 28169 2805 28181 2839
rect 28215 2836 28227 2839
rect 29546 2836 29552 2848
rect 28215 2808 29552 2836
rect 28215 2805 28227 2808
rect 28169 2799 28227 2805
rect 29546 2796 29552 2808
rect 29604 2796 29610 2848
rect 30190 2796 30196 2848
rect 30248 2836 30254 2848
rect 32125 2839 32183 2845
rect 32125 2836 32137 2839
rect 30248 2808 32137 2836
rect 30248 2796 30254 2808
rect 32125 2805 32137 2808
rect 32171 2805 32183 2839
rect 32125 2799 32183 2805
rect 34238 2796 34244 2848
rect 34296 2836 34302 2848
rect 34900 2836 34928 2876
rect 35805 2873 35817 2876
rect 35851 2873 35863 2907
rect 36446 2904 36452 2916
rect 36407 2876 36452 2904
rect 35805 2867 35863 2873
rect 36446 2864 36452 2876
rect 36504 2864 36510 2916
rect 36538 2864 36544 2916
rect 36596 2904 36602 2916
rect 38565 2907 38623 2913
rect 38565 2904 38577 2907
rect 36596 2876 38577 2904
rect 36596 2864 36602 2876
rect 38565 2873 38577 2876
rect 38611 2873 38623 2907
rect 38565 2867 38623 2873
rect 38654 2864 38660 2916
rect 38712 2904 38718 2916
rect 38712 2876 39344 2904
rect 38712 2864 38718 2876
rect 35342 2836 35348 2848
rect 34296 2808 34928 2836
rect 35303 2808 35348 2836
rect 34296 2796 34302 2808
rect 35342 2796 35348 2808
rect 35400 2796 35406 2848
rect 36722 2796 36728 2848
rect 36780 2836 36786 2848
rect 39209 2839 39267 2845
rect 39209 2836 39221 2839
rect 36780 2808 39221 2836
rect 36780 2796 36786 2808
rect 39209 2805 39221 2808
rect 39255 2805 39267 2839
rect 39316 2836 39344 2876
rect 41230 2864 41236 2916
rect 41288 2904 41294 2916
rect 41524 2904 41552 2944
rect 44361 2941 44373 2944
rect 44407 2941 44419 2975
rect 44361 2935 44419 2941
rect 43070 2904 43076 2916
rect 41288 2876 41552 2904
rect 43031 2876 43076 2904
rect 41288 2864 41294 2876
rect 43070 2864 43076 2876
rect 43128 2864 43134 2916
rect 44266 2904 44272 2916
rect 43180 2876 44272 2904
rect 41141 2839 41199 2845
rect 41141 2836 41153 2839
rect 39316 2808 41153 2836
rect 39209 2799 39267 2805
rect 41141 2805 41153 2808
rect 41187 2805 41199 2839
rect 42426 2836 42432 2848
rect 42387 2808 42432 2836
rect 41141 2799 41199 2805
rect 42426 2796 42432 2808
rect 42484 2796 42490 2848
rect 42794 2796 42800 2848
rect 42852 2836 42858 2848
rect 43180 2836 43208 2876
rect 44266 2864 44272 2876
rect 44324 2864 44330 2916
rect 42852 2808 43208 2836
rect 42852 2796 42858 2808
rect 43254 2796 43260 2848
rect 43312 2836 43318 2848
rect 45005 2839 45063 2845
rect 45005 2836 45017 2839
rect 43312 2808 45017 2836
rect 43312 2796 43318 2808
rect 45005 2805 45017 2808
rect 45051 2805 45063 2839
rect 45112 2836 45140 3012
rect 45186 3000 45192 3052
rect 45244 3040 45250 3052
rect 46308 3049 46336 3080
rect 47026 3068 47032 3080
rect 47084 3068 47090 3120
rect 49513 3111 49571 3117
rect 49513 3108 49525 3111
rect 47136 3080 49525 3108
rect 45649 3043 45707 3049
rect 45649 3040 45661 3043
rect 45244 3012 45661 3040
rect 45244 3000 45250 3012
rect 45649 3009 45661 3012
rect 45695 3009 45707 3043
rect 45649 3003 45707 3009
rect 46293 3043 46351 3049
rect 46293 3009 46305 3043
rect 46339 3009 46351 3043
rect 46293 3003 46351 3009
rect 46566 3000 46572 3052
rect 46624 3040 46630 3052
rect 47136 3040 47164 3080
rect 49513 3077 49525 3080
rect 49559 3108 49571 3111
rect 49878 3108 49884 3120
rect 49559 3080 49884 3108
rect 49559 3077 49571 3080
rect 49513 3071 49571 3077
rect 49878 3068 49884 3080
rect 49936 3068 49942 3120
rect 50062 3108 50068 3120
rect 50023 3080 50068 3108
rect 50062 3068 50068 3080
rect 50120 3068 50126 3120
rect 50706 3068 50712 3120
rect 50764 3108 50770 3120
rect 50764 3080 50936 3108
rect 50764 3068 50770 3080
rect 46624 3012 47164 3040
rect 46624 3000 46630 3012
rect 47210 3000 47216 3052
rect 47268 3040 47274 3052
rect 50798 3040 50804 3052
rect 47268 3012 50804 3040
rect 47268 3000 47274 3012
rect 50798 3000 50804 3012
rect 50856 3000 50862 3052
rect 50908 3049 50936 3080
rect 52454 3068 52460 3120
rect 52512 3108 52518 3120
rect 53944 3108 53972 3148
rect 55858 3108 55864 3120
rect 52512 3080 53972 3108
rect 54036 3080 55864 3108
rect 52512 3068 52518 3080
rect 50893 3043 50951 3049
rect 50893 3009 50905 3043
rect 50939 3009 50951 3043
rect 50893 3003 50951 3009
rect 51350 3000 51356 3052
rect 51408 3040 51414 3052
rect 54036 3040 54064 3080
rect 55858 3068 55864 3080
rect 55916 3068 55922 3120
rect 56042 3108 56048 3120
rect 56003 3080 56048 3108
rect 56042 3068 56048 3080
rect 56100 3068 56106 3120
rect 56137 3111 56195 3117
rect 56137 3077 56149 3111
rect 56183 3108 56195 3111
rect 56183 3080 56272 3108
rect 56183 3077 56195 3080
rect 56137 3071 56195 3077
rect 51408 3012 54064 3040
rect 54941 3043 54999 3049
rect 51408 3000 51414 3012
rect 54941 3009 54953 3043
rect 54987 3040 54999 3043
rect 55950 3040 55956 3052
rect 54987 3012 55956 3040
rect 54987 3009 54999 3012
rect 54941 3003 54999 3009
rect 55950 3000 55956 3012
rect 56008 3000 56014 3052
rect 56244 3040 56272 3080
rect 56318 3040 56324 3052
rect 56244 3012 56324 3040
rect 56318 3000 56324 3012
rect 56376 3000 56382 3052
rect 57900 3049 57928 3148
rect 57885 3043 57943 3049
rect 57885 3009 57897 3043
rect 57931 3009 57943 3043
rect 57885 3003 57943 3009
rect 45554 2932 45560 2984
rect 45612 2972 45618 2984
rect 48869 2975 48927 2981
rect 48869 2972 48881 2975
rect 45612 2944 48881 2972
rect 45612 2932 45618 2944
rect 48869 2941 48881 2944
rect 48915 2941 48927 2975
rect 53377 2975 53435 2981
rect 53377 2972 53389 2975
rect 48869 2935 48927 2941
rect 48976 2944 53389 2972
rect 45278 2864 45284 2916
rect 45336 2904 45342 2916
rect 48225 2907 48283 2913
rect 48225 2904 48237 2907
rect 45336 2876 48237 2904
rect 45336 2864 45342 2876
rect 48225 2873 48237 2876
rect 48271 2873 48283 2907
rect 48225 2867 48283 2873
rect 48590 2864 48596 2916
rect 48648 2904 48654 2916
rect 48976 2904 49004 2944
rect 53377 2941 53389 2944
rect 53423 2941 53435 2975
rect 53377 2935 53435 2941
rect 55217 2975 55275 2981
rect 55217 2941 55229 2975
rect 55263 2972 55275 2975
rect 55490 2972 55496 2984
rect 55263 2944 55496 2972
rect 55263 2941 55275 2944
rect 55217 2935 55275 2941
rect 55490 2932 55496 2944
rect 55548 2932 55554 2984
rect 56226 2932 56232 2984
rect 56284 2972 56290 2984
rect 56284 2944 56329 2972
rect 56284 2932 56290 2944
rect 48648 2876 49004 2904
rect 49160 2876 50936 2904
rect 48648 2864 48654 2876
rect 47581 2839 47639 2845
rect 47581 2836 47593 2839
rect 45112 2808 47593 2836
rect 45005 2799 45063 2805
rect 47581 2805 47593 2808
rect 47627 2805 47639 2839
rect 47581 2799 47639 2805
rect 47670 2796 47676 2848
rect 47728 2836 47734 2848
rect 49160 2836 49188 2876
rect 47728 2808 49188 2836
rect 47728 2796 47734 2808
rect 49878 2796 49884 2848
rect 49936 2836 49942 2848
rect 50249 2839 50307 2845
rect 50249 2836 50261 2839
rect 49936 2808 50261 2836
rect 49936 2796 49942 2808
rect 50249 2805 50261 2808
rect 50295 2836 50307 2839
rect 50430 2836 50436 2848
rect 50295 2808 50436 2836
rect 50295 2805 50307 2808
rect 50249 2799 50307 2805
rect 50430 2796 50436 2808
rect 50488 2796 50494 2848
rect 50908 2836 50936 2876
rect 50982 2864 50988 2916
rect 51040 2904 51046 2916
rect 51537 2907 51595 2913
rect 51537 2904 51549 2907
rect 51040 2876 51549 2904
rect 51040 2864 51046 2876
rect 51537 2873 51549 2876
rect 51583 2873 51595 2907
rect 51537 2867 51595 2873
rect 52362 2864 52368 2916
rect 52420 2904 52426 2916
rect 56873 2907 56931 2913
rect 56873 2904 56885 2907
rect 52420 2876 54340 2904
rect 52420 2864 52426 2876
rect 52733 2839 52791 2845
rect 52733 2836 52745 2839
rect 50908 2808 52745 2836
rect 52733 2805 52745 2808
rect 52779 2805 52791 2839
rect 54202 2836 54208 2848
rect 54163 2808 54208 2836
rect 52733 2799 52791 2805
rect 54202 2796 54208 2808
rect 54260 2796 54266 2848
rect 54312 2836 54340 2876
rect 55186 2876 56885 2904
rect 55186 2836 55214 2876
rect 56873 2873 56885 2876
rect 56919 2873 56931 2907
rect 56873 2867 56931 2873
rect 54312 2808 55214 2836
rect 55582 2796 55588 2848
rect 55640 2836 55646 2848
rect 55677 2839 55735 2845
rect 55677 2836 55689 2839
rect 55640 2808 55689 2836
rect 55640 2796 55646 2808
rect 55677 2805 55689 2808
rect 55723 2805 55735 2839
rect 55677 2799 55735 2805
rect 55766 2796 55772 2848
rect 55824 2836 55830 2848
rect 56594 2836 56600 2848
rect 55824 2808 56600 2836
rect 55824 2796 55830 2808
rect 56594 2796 56600 2808
rect 56652 2796 56658 2848
rect 1104 2746 58880 2768
rect 1104 2694 8174 2746
rect 8226 2694 8238 2746
rect 8290 2694 8302 2746
rect 8354 2694 8366 2746
rect 8418 2694 8430 2746
rect 8482 2694 22622 2746
rect 22674 2694 22686 2746
rect 22738 2694 22750 2746
rect 22802 2694 22814 2746
rect 22866 2694 22878 2746
rect 22930 2694 37070 2746
rect 37122 2694 37134 2746
rect 37186 2694 37198 2746
rect 37250 2694 37262 2746
rect 37314 2694 37326 2746
rect 37378 2694 51518 2746
rect 51570 2694 51582 2746
rect 51634 2694 51646 2746
rect 51698 2694 51710 2746
rect 51762 2694 51774 2746
rect 51826 2694 58880 2746
rect 1104 2672 58880 2694
rect 4065 2635 4123 2641
rect 4065 2601 4077 2635
rect 4111 2632 4123 2635
rect 4614 2632 4620 2644
rect 4111 2604 4620 2632
rect 4111 2601 4123 2604
rect 4065 2595 4123 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 5074 2592 5080 2644
rect 5132 2632 5138 2644
rect 5534 2632 5540 2644
rect 5132 2604 5540 2632
rect 5132 2592 5138 2604
rect 5534 2592 5540 2604
rect 5592 2632 5598 2644
rect 7282 2632 7288 2644
rect 5592 2604 7288 2632
rect 5592 2592 5598 2604
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 7484 2604 9674 2632
rect 2593 2567 2651 2573
rect 2593 2533 2605 2567
rect 2639 2533 2651 2567
rect 5442 2564 5448 2576
rect 2593 2527 2651 2533
rect 2746 2536 5448 2564
rect 2608 2496 2636 2527
rect 2746 2496 2774 2536
rect 5442 2524 5448 2536
rect 5500 2524 5506 2576
rect 5813 2567 5871 2573
rect 5813 2533 5825 2567
rect 5859 2564 5871 2567
rect 7098 2564 7104 2576
rect 5859 2536 7104 2564
rect 5859 2533 5871 2536
rect 5813 2527 5871 2533
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 2608 2468 2774 2496
rect 2866 2456 2872 2508
rect 2924 2496 2930 2508
rect 5169 2499 5227 2505
rect 2924 2468 4936 2496
rect 2924 2456 2930 2468
rect 2406 2428 2412 2440
rect 2367 2400 2412 2428
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 3050 2428 3056 2440
rect 3011 2400 3056 2428
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3878 2428 3884 2440
rect 3839 2400 3884 2428
rect 3878 2388 3884 2400
rect 3936 2388 3942 2440
rect 4706 2428 4712 2440
rect 4667 2400 4712 2428
rect 4706 2388 4712 2400
rect 4764 2388 4770 2440
rect 1949 2363 2007 2369
rect 1949 2329 1961 2363
rect 1995 2360 2007 2363
rect 3896 2360 3924 2388
rect 1995 2332 3924 2360
rect 4908 2360 4936 2468
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5258 2496 5264 2508
rect 5215 2468 5264 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 5626 2456 5632 2508
rect 5684 2505 5690 2508
rect 5684 2499 5712 2505
rect 5700 2465 5712 2499
rect 5684 2459 5712 2465
rect 6641 2499 6699 2505
rect 6641 2465 6653 2499
rect 6687 2496 6699 2499
rect 7484 2496 7512 2604
rect 9646 2564 9674 2604
rect 10410 2592 10416 2644
rect 10468 2632 10474 2644
rect 11517 2635 11575 2641
rect 11517 2632 11529 2635
rect 10468 2604 11529 2632
rect 10468 2592 10474 2604
rect 10502 2564 10508 2576
rect 9646 2536 10508 2564
rect 10502 2524 10508 2536
rect 10560 2524 10566 2576
rect 6687 2468 7512 2496
rect 6687 2465 6699 2468
rect 6641 2459 6699 2465
rect 5684 2456 5690 2459
rect 8846 2456 8852 2508
rect 8904 2496 8910 2508
rect 10888 2496 10916 2604
rect 11517 2601 11529 2604
rect 11563 2601 11575 2635
rect 11517 2595 11575 2601
rect 11606 2592 11612 2644
rect 11664 2632 11670 2644
rect 13173 2635 13231 2641
rect 11664 2604 13124 2632
rect 11664 2592 11670 2604
rect 10965 2567 11023 2573
rect 10965 2533 10977 2567
rect 11011 2564 11023 2567
rect 13096 2564 13124 2604
rect 13173 2601 13185 2635
rect 13219 2632 13231 2635
rect 13262 2632 13268 2644
rect 13219 2604 13268 2632
rect 13219 2601 13231 2604
rect 13173 2595 13231 2601
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 14056 2604 14197 2632
rect 14056 2592 14062 2604
rect 14185 2601 14197 2604
rect 14231 2632 14243 2635
rect 16482 2632 16488 2644
rect 14231 2604 16488 2632
rect 14231 2601 14243 2604
rect 14185 2595 14243 2601
rect 16482 2592 16488 2604
rect 16540 2592 16546 2644
rect 17405 2635 17463 2641
rect 17405 2601 17417 2635
rect 17451 2632 17463 2635
rect 20714 2632 20720 2644
rect 17451 2604 20720 2632
rect 17451 2601 17463 2604
rect 17405 2595 17463 2601
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 22189 2635 22247 2641
rect 22189 2601 22201 2635
rect 22235 2632 22247 2635
rect 24578 2632 24584 2644
rect 22235 2604 24584 2632
rect 22235 2601 22247 2604
rect 22189 2595 22247 2601
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 25777 2635 25835 2641
rect 25777 2601 25789 2635
rect 25823 2632 25835 2635
rect 26694 2632 26700 2644
rect 25823 2604 26700 2632
rect 25823 2601 25835 2604
rect 25777 2595 25835 2601
rect 26694 2592 26700 2604
rect 26752 2592 26758 2644
rect 33870 2592 33876 2644
rect 33928 2632 33934 2644
rect 34057 2635 34115 2641
rect 34057 2632 34069 2635
rect 33928 2604 34069 2632
rect 33928 2592 33934 2604
rect 34057 2601 34069 2604
rect 34103 2601 34115 2635
rect 34057 2595 34115 2601
rect 34514 2592 34520 2644
rect 34572 2632 34578 2644
rect 34701 2635 34759 2641
rect 34701 2632 34713 2635
rect 34572 2604 34713 2632
rect 34572 2592 34578 2604
rect 34701 2601 34713 2604
rect 34747 2601 34759 2635
rect 34701 2595 34759 2601
rect 34790 2592 34796 2644
rect 34848 2632 34854 2644
rect 35345 2635 35403 2641
rect 35345 2632 35357 2635
rect 34848 2604 35357 2632
rect 34848 2592 34854 2604
rect 35345 2601 35357 2604
rect 35391 2601 35403 2635
rect 35345 2595 35403 2601
rect 36814 2592 36820 2644
rect 36872 2632 36878 2644
rect 37921 2635 37979 2641
rect 37921 2632 37933 2635
rect 36872 2604 37933 2632
rect 36872 2592 36878 2604
rect 37921 2601 37933 2604
rect 37967 2601 37979 2635
rect 37921 2595 37979 2601
rect 38010 2592 38016 2644
rect 38068 2632 38074 2644
rect 38838 2632 38844 2644
rect 38068 2604 38844 2632
rect 38068 2592 38074 2604
rect 38838 2592 38844 2604
rect 38896 2632 38902 2644
rect 39209 2635 39267 2641
rect 39209 2632 39221 2635
rect 38896 2604 39221 2632
rect 38896 2592 38902 2604
rect 39209 2601 39221 2604
rect 39255 2601 39267 2635
rect 39209 2595 39267 2601
rect 40310 2592 40316 2644
rect 40368 2632 40374 2644
rect 43717 2635 43775 2641
rect 43717 2632 43729 2635
rect 40368 2604 43729 2632
rect 40368 2592 40374 2604
rect 43717 2601 43729 2604
rect 43763 2601 43775 2635
rect 43717 2595 43775 2601
rect 44266 2592 44272 2644
rect 44324 2632 44330 2644
rect 47581 2635 47639 2641
rect 47581 2632 47593 2635
rect 44324 2604 47593 2632
rect 44324 2592 44330 2604
rect 47581 2601 47593 2604
rect 47627 2601 47639 2635
rect 49510 2632 49516 2644
rect 49471 2604 49516 2632
rect 47581 2595 47639 2601
rect 49510 2592 49516 2604
rect 49568 2592 49574 2644
rect 49602 2592 49608 2644
rect 49660 2632 49666 2644
rect 53377 2635 53435 2641
rect 53377 2632 53389 2635
rect 49660 2604 53389 2632
rect 49660 2592 49666 2604
rect 53377 2601 53389 2604
rect 53423 2601 53435 2635
rect 55585 2635 55643 2641
rect 55585 2632 55597 2635
rect 53377 2595 53435 2601
rect 55186 2604 55597 2632
rect 14090 2564 14096 2576
rect 11011 2536 13032 2564
rect 13096 2536 14096 2564
rect 11011 2533 11023 2536
rect 10965 2527 11023 2533
rect 12618 2496 12624 2508
rect 8904 2468 9720 2496
rect 10888 2468 12624 2496
rect 8904 2456 8910 2468
rect 4982 2388 4988 2440
rect 5040 2428 5046 2440
rect 6549 2431 6607 2437
rect 6549 2430 6561 2431
rect 6472 2428 6561 2430
rect 5040 2402 6561 2428
rect 5040 2400 6500 2402
rect 5040 2388 5046 2400
rect 6549 2397 6561 2402
rect 6595 2397 6607 2431
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6549 2391 6607 2397
rect 6656 2400 6745 2428
rect 4908 2332 5672 2360
rect 1995 2329 2007 2332
rect 1949 2323 2007 2329
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 4338 2292 4344 2304
rect 3283 2264 4344 2292
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 4338 2252 4344 2264
rect 4396 2292 4402 2304
rect 5350 2292 5356 2304
rect 4396 2264 5356 2292
rect 4396 2252 4402 2264
rect 5350 2252 5356 2264
rect 5408 2292 5414 2304
rect 5445 2295 5503 2301
rect 5445 2292 5457 2295
rect 5408 2264 5457 2292
rect 5408 2252 5414 2264
rect 5445 2261 5457 2264
rect 5491 2261 5503 2295
rect 5644 2292 5672 2332
rect 5718 2320 5724 2372
rect 5776 2360 5782 2372
rect 6656 2360 6684 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 7374 2388 7380 2440
rect 7432 2428 7438 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7432 2400 7481 2428
rect 7432 2388 7438 2400
rect 7469 2397 7481 2400
rect 7515 2397 7527 2431
rect 9214 2428 9220 2440
rect 9175 2400 9220 2428
rect 7469 2391 7527 2397
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 9692 2437 9720 2468
rect 12618 2456 12624 2468
rect 12676 2456 12682 2508
rect 13004 2496 13032 2536
rect 14090 2524 14096 2536
rect 14148 2524 14154 2576
rect 15473 2567 15531 2573
rect 15473 2533 15485 2567
rect 15519 2564 15531 2567
rect 19058 2564 19064 2576
rect 15519 2536 19064 2564
rect 15519 2533 15531 2536
rect 15473 2527 15531 2533
rect 19058 2524 19064 2536
rect 19116 2524 19122 2576
rect 20625 2567 20683 2573
rect 20625 2533 20637 2567
rect 20671 2564 20683 2567
rect 22646 2564 22652 2576
rect 20671 2536 22652 2564
rect 20671 2533 20683 2536
rect 20625 2527 20683 2533
rect 22646 2524 22652 2536
rect 22704 2524 22710 2576
rect 23753 2567 23811 2573
rect 23753 2533 23765 2567
rect 23799 2564 23811 2567
rect 25130 2564 25136 2576
rect 23799 2536 25136 2564
rect 23799 2533 23811 2536
rect 23753 2527 23811 2533
rect 25130 2524 25136 2536
rect 25188 2524 25194 2576
rect 26145 2567 26203 2573
rect 26145 2533 26157 2567
rect 26191 2564 26203 2567
rect 26602 2564 26608 2576
rect 26191 2536 26608 2564
rect 26191 2533 26203 2536
rect 26145 2527 26203 2533
rect 26602 2524 26608 2536
rect 26660 2524 26666 2576
rect 28997 2567 29055 2573
rect 28997 2533 29009 2567
rect 29043 2564 29055 2567
rect 30374 2564 30380 2576
rect 29043 2536 30380 2564
rect 29043 2533 29055 2536
rect 28997 2527 29055 2533
rect 30374 2524 30380 2536
rect 30432 2524 30438 2576
rect 32030 2524 32036 2576
rect 32088 2564 32094 2576
rect 33413 2567 33471 2573
rect 33413 2564 33425 2567
rect 32088 2536 33425 2564
rect 32088 2524 32094 2536
rect 33413 2533 33425 2536
rect 33459 2533 33471 2567
rect 33413 2527 33471 2533
rect 33686 2524 33692 2576
rect 33744 2564 33750 2576
rect 37277 2567 37335 2573
rect 37277 2564 37289 2567
rect 33744 2536 37289 2564
rect 33744 2524 33750 2536
rect 37277 2533 37289 2536
rect 37323 2533 37335 2567
rect 37277 2527 37335 2533
rect 37826 2524 37832 2576
rect 37884 2564 37890 2576
rect 41141 2567 41199 2573
rect 41141 2564 41153 2567
rect 37884 2536 41153 2564
rect 37884 2524 37890 2536
rect 41141 2533 41153 2536
rect 41187 2533 41199 2567
rect 45005 2567 45063 2573
rect 45005 2564 45017 2567
rect 41141 2527 41199 2533
rect 41248 2536 45017 2564
rect 15562 2496 15568 2508
rect 13004 2468 15568 2496
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 18049 2499 18107 2505
rect 18049 2465 18061 2499
rect 18095 2496 18107 2499
rect 18414 2496 18420 2508
rect 18095 2468 18420 2496
rect 18095 2465 18107 2468
rect 18049 2459 18107 2465
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 18693 2499 18751 2505
rect 18693 2465 18705 2499
rect 18739 2465 18751 2499
rect 18693 2459 18751 2465
rect 19981 2499 20039 2505
rect 19981 2465 19993 2499
rect 20027 2496 20039 2499
rect 21269 2499 21327 2505
rect 20027 2468 21036 2496
rect 20027 2465 20039 2468
rect 19981 2459 20039 2465
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 10781 2431 10839 2437
rect 10781 2397 10793 2431
rect 10827 2397 10839 2431
rect 12250 2428 12256 2440
rect 12211 2400 12256 2428
rect 10781 2391 10839 2397
rect 5776 2332 6684 2360
rect 5776 2320 5782 2332
rect 7098 2320 7104 2372
rect 7156 2360 7162 2372
rect 10796 2360 10824 2391
rect 12250 2388 12256 2400
rect 12308 2388 12314 2440
rect 12710 2428 12716 2440
rect 12671 2400 12716 2428
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 12952 2400 13093 2428
rect 12952 2388 12958 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13354 2428 13360 2440
rect 13315 2400 13360 2428
rect 13081 2391 13139 2397
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2428 16175 2431
rect 18322 2428 18328 2440
rect 16163 2400 18328 2428
rect 16163 2397 16175 2400
rect 16117 2391 16175 2397
rect 13998 2360 14004 2372
rect 7156 2332 9996 2360
rect 10796 2332 14004 2360
rect 7156 2320 7162 2332
rect 7742 2301 7748 2304
rect 7699 2295 7748 2301
rect 7699 2292 7711 2295
rect 5644 2264 7711 2292
rect 5445 2255 5503 2261
rect 7699 2261 7711 2264
rect 7745 2261 7748 2295
rect 7699 2255 7748 2261
rect 7742 2252 7748 2255
rect 7800 2292 7806 2304
rect 7800 2264 7847 2292
rect 7800 2252 7806 2264
rect 8754 2252 8760 2304
rect 8812 2292 8818 2304
rect 9033 2295 9091 2301
rect 9033 2292 9045 2295
rect 8812 2264 9045 2292
rect 8812 2252 8818 2264
rect 9033 2261 9045 2264
rect 9079 2261 9091 2295
rect 9033 2255 9091 2261
rect 9214 2252 9220 2304
rect 9272 2292 9278 2304
rect 9861 2295 9919 2301
rect 9861 2292 9873 2295
rect 9272 2264 9873 2292
rect 9272 2252 9278 2264
rect 9861 2261 9873 2264
rect 9907 2261 9919 2295
rect 9968 2292 9996 2332
rect 13998 2320 14004 2332
rect 14056 2320 14062 2372
rect 11606 2292 11612 2304
rect 9968 2264 11612 2292
rect 9861 2255 9919 2261
rect 11606 2252 11612 2264
rect 11664 2252 11670 2304
rect 12897 2295 12955 2301
rect 12897 2261 12909 2295
rect 12943 2292 12955 2295
rect 13170 2292 13176 2304
rect 12943 2264 13176 2292
rect 12943 2261 12955 2264
rect 12897 2255 12955 2261
rect 13170 2252 13176 2264
rect 13228 2252 13234 2304
rect 14844 2292 14872 2391
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 18708 2360 18736 2459
rect 21008 2428 21036 2468
rect 21269 2465 21281 2499
rect 21315 2496 21327 2499
rect 22922 2496 22928 2508
rect 21315 2468 22928 2496
rect 21315 2465 21327 2468
rect 21269 2459 21327 2465
rect 22922 2456 22928 2468
rect 22980 2456 22986 2508
rect 23032 2468 23612 2496
rect 22278 2428 22284 2440
rect 21008 2400 22284 2428
rect 22278 2388 22284 2400
rect 22336 2388 22342 2440
rect 22373 2431 22431 2437
rect 22373 2397 22385 2431
rect 22419 2428 22431 2431
rect 22462 2428 22468 2440
rect 22419 2400 22468 2428
rect 22419 2397 22431 2400
rect 22373 2391 22431 2397
rect 22462 2388 22468 2400
rect 22520 2388 22526 2440
rect 23032 2428 23060 2468
rect 22848 2400 23060 2428
rect 23109 2431 23167 2437
rect 22094 2360 22100 2372
rect 18708 2332 22100 2360
rect 22094 2320 22100 2332
rect 22152 2320 22158 2372
rect 18782 2292 18788 2304
rect 14844 2264 18788 2292
rect 18782 2252 18788 2264
rect 18840 2252 18846 2304
rect 19337 2295 19395 2301
rect 19337 2261 19349 2295
rect 19383 2292 19395 2295
rect 22848 2292 22876 2400
rect 23109 2397 23121 2431
rect 23155 2428 23167 2431
rect 23290 2428 23296 2440
rect 23155 2400 23296 2428
rect 23155 2397 23167 2400
rect 23109 2391 23167 2397
rect 23290 2388 23296 2400
rect 23348 2388 23354 2440
rect 23584 2437 23612 2468
rect 24210 2456 24216 2508
rect 24268 2496 24274 2508
rect 24489 2499 24547 2505
rect 24489 2496 24501 2499
rect 24268 2468 24501 2496
rect 24268 2456 24274 2468
rect 24489 2465 24501 2468
rect 24535 2465 24547 2499
rect 24670 2496 24676 2508
rect 24631 2468 24676 2496
rect 24489 2459 24547 2465
rect 24670 2456 24676 2468
rect 24728 2456 24734 2508
rect 24762 2456 24768 2508
rect 24820 2496 24826 2508
rect 26970 2496 26976 2508
rect 24820 2468 26234 2496
rect 26931 2468 26976 2496
rect 24820 2456 24826 2468
rect 23569 2431 23627 2437
rect 23569 2397 23581 2431
rect 23615 2428 23627 2431
rect 23658 2428 23664 2440
rect 23615 2400 23664 2428
rect 23615 2397 23627 2400
rect 23569 2391 23627 2397
rect 23658 2388 23664 2400
rect 23716 2388 23722 2440
rect 26206 2428 26234 2468
rect 26970 2456 26976 2468
rect 27028 2456 27034 2508
rect 29270 2456 29276 2508
rect 29328 2496 29334 2508
rect 30285 2499 30343 2505
rect 30285 2496 30297 2499
rect 29328 2468 30297 2496
rect 29328 2456 29334 2468
rect 30285 2465 30297 2468
rect 30331 2465 30343 2499
rect 30285 2459 30343 2465
rect 30650 2456 30656 2508
rect 30708 2496 30714 2508
rect 32125 2499 32183 2505
rect 32125 2496 32137 2499
rect 30708 2468 32137 2496
rect 30708 2456 30714 2468
rect 32125 2465 32137 2468
rect 32171 2465 32183 2499
rect 36262 2496 36268 2508
rect 32125 2459 32183 2465
rect 32876 2468 36268 2496
rect 27229 2431 27287 2437
rect 27229 2428 27241 2431
rect 26206 2400 27241 2428
rect 27229 2397 27241 2400
rect 27275 2397 27287 2431
rect 27229 2391 27287 2397
rect 29825 2431 29883 2437
rect 29825 2397 29837 2431
rect 29871 2397 29883 2431
rect 29825 2391 29883 2397
rect 24854 2360 24860 2372
rect 22940 2332 24860 2360
rect 22940 2301 22968 2332
rect 24854 2320 24860 2332
rect 24912 2320 24918 2372
rect 26326 2360 26332 2372
rect 25148 2332 26332 2360
rect 19383 2264 22876 2292
rect 22925 2295 22983 2301
rect 19383 2261 19395 2264
rect 19337 2255 19395 2261
rect 22925 2261 22937 2295
rect 22971 2261 22983 2295
rect 22925 2255 22983 2261
rect 24486 2252 24492 2304
rect 24544 2292 24550 2304
rect 25148 2301 25176 2332
rect 26326 2320 26332 2332
rect 26384 2320 26390 2372
rect 27522 2320 27528 2372
rect 27580 2360 27586 2372
rect 29840 2360 29868 2391
rect 30926 2388 30932 2440
rect 30984 2428 30990 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30984 2400 31033 2428
rect 30984 2388 30990 2400
rect 31021 2397 31033 2400
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 31202 2388 31208 2440
rect 31260 2428 31266 2440
rect 32769 2431 32827 2437
rect 32769 2428 32781 2431
rect 31260 2400 32781 2428
rect 31260 2388 31266 2400
rect 32769 2397 32781 2400
rect 32815 2397 32827 2431
rect 32769 2391 32827 2397
rect 32876 2360 32904 2468
rect 36262 2456 36268 2468
rect 36320 2496 36326 2508
rect 36320 2468 36768 2496
rect 36320 2456 36326 2468
rect 32950 2388 32956 2440
rect 33008 2428 33014 2440
rect 36740 2437 36768 2468
rect 37366 2456 37372 2508
rect 37424 2496 37430 2508
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 37424 2468 40509 2496
rect 37424 2456 37430 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 40497 2459 40555 2465
rect 40862 2456 40868 2508
rect 40920 2496 40926 2508
rect 41248 2496 41276 2536
rect 45005 2533 45017 2536
rect 45051 2533 45063 2567
rect 45005 2527 45063 2533
rect 45186 2524 45192 2576
rect 45244 2564 45250 2576
rect 45649 2567 45707 2573
rect 45649 2564 45661 2567
rect 45244 2536 45661 2564
rect 45244 2524 45250 2536
rect 45649 2533 45661 2536
rect 45695 2533 45707 2567
rect 45649 2527 45707 2533
rect 45830 2524 45836 2576
rect 45888 2564 45894 2576
rect 50157 2567 50215 2573
rect 50157 2564 50169 2567
rect 45888 2536 50169 2564
rect 45888 2524 45894 2536
rect 50157 2533 50169 2536
rect 50203 2533 50215 2567
rect 50157 2527 50215 2533
rect 50430 2524 50436 2576
rect 50488 2564 50494 2576
rect 54665 2567 54723 2573
rect 54665 2564 54677 2567
rect 50488 2536 54677 2564
rect 50488 2524 50494 2536
rect 54665 2533 54677 2536
rect 54711 2564 54723 2567
rect 55186 2564 55214 2604
rect 55585 2601 55597 2604
rect 55631 2632 55643 2635
rect 55769 2635 55827 2641
rect 55631 2604 55720 2632
rect 55631 2601 55643 2604
rect 55585 2595 55643 2601
rect 54711 2536 55214 2564
rect 54711 2533 54723 2536
rect 54665 2527 54723 2533
rect 40920 2468 41276 2496
rect 44453 2499 44511 2505
rect 40920 2456 40926 2468
rect 44453 2465 44465 2499
rect 44499 2496 44511 2499
rect 44542 2496 44548 2508
rect 44499 2468 44548 2496
rect 44499 2465 44511 2468
rect 44453 2459 44511 2465
rect 44542 2456 44548 2468
rect 44600 2456 44606 2508
rect 44634 2456 44640 2508
rect 44692 2496 44698 2508
rect 48225 2499 48283 2505
rect 48225 2496 48237 2499
rect 44692 2468 48237 2496
rect 44692 2456 44698 2468
rect 48225 2465 48237 2468
rect 48271 2465 48283 2499
rect 48225 2459 48283 2465
rect 49694 2456 49700 2508
rect 49752 2496 49758 2508
rect 54021 2499 54079 2505
rect 54021 2496 54033 2499
rect 49752 2468 54033 2496
rect 49752 2456 49758 2468
rect 54021 2465 54033 2468
rect 54067 2465 54079 2499
rect 55692 2496 55720 2604
rect 55769 2601 55781 2635
rect 55815 2632 55827 2635
rect 57422 2632 57428 2644
rect 55815 2604 57428 2632
rect 55815 2601 55827 2604
rect 55769 2595 55827 2601
rect 57422 2592 57428 2604
rect 57480 2592 57486 2644
rect 55858 2524 55864 2576
rect 55916 2564 55922 2576
rect 57885 2567 57943 2573
rect 57885 2564 57897 2567
rect 55916 2536 57897 2564
rect 55916 2524 55922 2536
rect 57885 2533 57897 2536
rect 57931 2533 57943 2567
rect 57885 2527 57943 2533
rect 56686 2496 56692 2508
rect 55692 2468 56692 2496
rect 54021 2459 54079 2465
rect 56686 2456 56692 2468
rect 56744 2456 56750 2508
rect 35989 2431 36047 2437
rect 35989 2428 36001 2431
rect 33008 2400 36001 2428
rect 33008 2388 33014 2400
rect 35989 2397 36001 2400
rect 36035 2397 36047 2431
rect 35989 2391 36047 2397
rect 36725 2431 36783 2437
rect 36725 2397 36737 2431
rect 36771 2428 36783 2431
rect 38010 2428 38016 2440
rect 36771 2400 38016 2428
rect 36771 2397 36783 2400
rect 36725 2391 36783 2397
rect 38010 2388 38016 2400
rect 38068 2388 38074 2440
rect 38565 2431 38623 2437
rect 38565 2397 38577 2431
rect 38611 2397 38623 2431
rect 39853 2431 39911 2437
rect 39853 2428 39865 2431
rect 38565 2391 38623 2397
rect 38672 2400 39865 2428
rect 27580 2332 29684 2360
rect 29840 2332 32904 2360
rect 27580 2320 27586 2332
rect 24765 2295 24823 2301
rect 24765 2292 24777 2295
rect 24544 2264 24777 2292
rect 24544 2252 24550 2264
rect 24765 2261 24777 2264
rect 24811 2261 24823 2295
rect 24765 2255 24823 2261
rect 25133 2295 25191 2301
rect 25133 2261 25145 2295
rect 25179 2261 25191 2295
rect 25590 2292 25596 2304
rect 25551 2264 25596 2292
rect 25133 2255 25191 2261
rect 25590 2252 25596 2264
rect 25648 2252 25654 2304
rect 25774 2292 25780 2304
rect 25735 2264 25780 2292
rect 25774 2252 25780 2264
rect 25832 2252 25838 2304
rect 28350 2292 28356 2304
rect 28311 2264 28356 2292
rect 28350 2252 28356 2264
rect 28408 2252 28414 2304
rect 29656 2301 29684 2332
rect 35434 2320 35440 2372
rect 35492 2360 35498 2372
rect 38580 2360 38608 2391
rect 35492 2332 38608 2360
rect 35492 2320 35498 2332
rect 29641 2295 29699 2301
rect 29641 2261 29653 2295
rect 29687 2261 29699 2295
rect 29641 2255 29699 2261
rect 33870 2252 33876 2304
rect 33928 2292 33934 2304
rect 36998 2292 37004 2304
rect 33928 2264 37004 2292
rect 33928 2252 33934 2264
rect 36998 2252 37004 2264
rect 37056 2252 37062 2304
rect 37090 2252 37096 2304
rect 37148 2292 37154 2304
rect 38672 2292 38700 2400
rect 39853 2397 39865 2400
rect 39899 2397 39911 2431
rect 39853 2391 39911 2397
rect 39942 2388 39948 2440
rect 40000 2428 40006 2440
rect 42429 2431 42487 2437
rect 42429 2428 42441 2431
rect 40000 2400 42441 2428
rect 40000 2388 40006 2400
rect 42429 2397 42441 2400
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 43073 2431 43131 2437
rect 43073 2397 43085 2431
rect 43119 2397 43131 2431
rect 46293 2431 46351 2437
rect 46293 2428 46305 2431
rect 43073 2391 43131 2397
rect 43272 2400 46305 2428
rect 39758 2320 39764 2372
rect 39816 2360 39822 2372
rect 43088 2360 43116 2391
rect 39816 2332 43116 2360
rect 39816 2320 39822 2332
rect 37148 2264 38700 2292
rect 37148 2252 37154 2264
rect 40126 2252 40132 2304
rect 40184 2292 40190 2304
rect 41785 2295 41843 2301
rect 41785 2292 41797 2295
rect 40184 2264 41797 2292
rect 40184 2252 40190 2264
rect 41785 2261 41797 2264
rect 41831 2261 41843 2295
rect 41785 2255 41843 2261
rect 41966 2252 41972 2304
rect 42024 2292 42030 2304
rect 43272 2292 43300 2400
rect 46293 2397 46305 2400
rect 46339 2397 46351 2431
rect 46293 2391 46351 2397
rect 46842 2388 46848 2440
rect 46900 2428 46906 2440
rect 48869 2431 48927 2437
rect 48869 2428 48881 2431
rect 46900 2400 48881 2428
rect 46900 2388 46906 2400
rect 48869 2397 48881 2400
rect 48915 2397 48927 2431
rect 48869 2391 48927 2397
rect 50801 2431 50859 2437
rect 50801 2397 50813 2431
rect 50847 2397 50859 2431
rect 51442 2428 51448 2440
rect 51403 2400 51448 2428
rect 50801 2391 50859 2397
rect 45278 2320 45284 2372
rect 45336 2360 45342 2372
rect 50816 2360 50844 2391
rect 51442 2388 51448 2400
rect 51500 2388 51506 2440
rect 52730 2428 52736 2440
rect 52691 2400 52736 2428
rect 52730 2388 52736 2400
rect 52788 2388 52794 2440
rect 54754 2388 54760 2440
rect 54812 2428 54818 2440
rect 55309 2431 55367 2437
rect 55309 2428 55321 2431
rect 54812 2400 55321 2428
rect 54812 2388 54818 2400
rect 55309 2397 55321 2400
rect 55355 2397 55367 2431
rect 56226 2428 56232 2440
rect 56187 2400 56232 2428
rect 55309 2391 55367 2397
rect 56226 2388 56232 2400
rect 56284 2388 56290 2440
rect 56873 2431 56931 2437
rect 56873 2397 56885 2431
rect 56919 2397 56931 2431
rect 56873 2391 56931 2397
rect 56888 2360 56916 2391
rect 45336 2332 50844 2360
rect 50908 2332 56916 2360
rect 45336 2320 45342 2332
rect 42024 2264 43300 2292
rect 42024 2252 42030 2264
rect 44818 2252 44824 2304
rect 44876 2292 44882 2304
rect 45462 2292 45468 2304
rect 44876 2264 45468 2292
rect 44876 2252 44882 2264
rect 45462 2252 45468 2264
rect 45520 2292 45526 2304
rect 47029 2295 47087 2301
rect 47029 2292 47041 2295
rect 45520 2264 47041 2292
rect 45520 2252 45526 2264
rect 47029 2261 47041 2264
rect 47075 2292 47087 2295
rect 47578 2292 47584 2304
rect 47075 2264 47584 2292
rect 47075 2261 47087 2264
rect 47029 2255 47087 2261
rect 47578 2252 47584 2264
rect 47636 2252 47642 2304
rect 50798 2252 50804 2304
rect 50856 2292 50862 2304
rect 50908 2292 50936 2332
rect 50856 2264 50936 2292
rect 50856 2252 50862 2264
rect 51166 2252 51172 2304
rect 51224 2292 51230 2304
rect 52089 2295 52147 2301
rect 52089 2292 52101 2295
rect 51224 2264 52101 2292
rect 51224 2252 51230 2264
rect 52089 2261 52101 2264
rect 52135 2261 52147 2295
rect 52089 2255 52147 2261
rect 1104 2202 58880 2224
rect 1104 2150 15398 2202
rect 15450 2150 15462 2202
rect 15514 2150 15526 2202
rect 15578 2150 15590 2202
rect 15642 2150 15654 2202
rect 15706 2150 29846 2202
rect 29898 2150 29910 2202
rect 29962 2150 29974 2202
rect 30026 2150 30038 2202
rect 30090 2150 30102 2202
rect 30154 2150 44294 2202
rect 44346 2150 44358 2202
rect 44410 2150 44422 2202
rect 44474 2150 44486 2202
rect 44538 2150 44550 2202
rect 44602 2150 58880 2202
rect 1104 2128 58880 2150
rect 3878 2048 3884 2100
rect 3936 2088 3942 2100
rect 8938 2088 8944 2100
rect 3936 2060 8944 2088
rect 3936 2048 3942 2060
rect 8938 2048 8944 2060
rect 8996 2048 9002 2100
rect 10502 2048 10508 2100
rect 10560 2088 10566 2100
rect 10560 2060 11284 2088
rect 10560 2048 10566 2060
rect 4706 1980 4712 2032
rect 4764 2020 4770 2032
rect 11146 2020 11152 2032
rect 4764 1992 11152 2020
rect 4764 1980 4770 1992
rect 11146 1980 11152 1992
rect 11204 1980 11210 2032
rect 11256 2020 11284 2060
rect 12250 2048 12256 2100
rect 12308 2088 12314 2100
rect 18230 2088 18236 2100
rect 12308 2060 18236 2088
rect 12308 2048 12314 2060
rect 18230 2048 18236 2060
rect 18288 2048 18294 2100
rect 18414 2048 18420 2100
rect 18472 2088 18478 2100
rect 21542 2088 21548 2100
rect 18472 2060 21548 2088
rect 18472 2048 18478 2060
rect 21542 2048 21548 2060
rect 21600 2048 21606 2100
rect 36998 2048 37004 2100
rect 37056 2088 37062 2100
rect 40126 2088 40132 2100
rect 37056 2060 40132 2088
rect 37056 2048 37062 2060
rect 40126 2048 40132 2060
rect 40184 2048 40190 2100
rect 41414 2048 41420 2100
rect 41472 2088 41478 2100
rect 45186 2088 45192 2100
rect 41472 2060 45192 2088
rect 41472 2048 41478 2060
rect 45186 2048 45192 2060
rect 45244 2048 45250 2100
rect 46382 2048 46388 2100
rect 46440 2088 46446 2100
rect 51442 2088 51448 2100
rect 46440 2060 51448 2088
rect 46440 2048 46446 2060
rect 51442 2048 51448 2060
rect 51500 2048 51506 2100
rect 13814 2020 13820 2032
rect 11256 1992 13820 2020
rect 13814 1980 13820 1992
rect 13872 1980 13878 2032
rect 18322 1980 18328 2032
rect 18380 2020 18386 2032
rect 20162 2020 20168 2032
rect 18380 1992 20168 2020
rect 18380 1980 18386 1992
rect 20162 1980 20168 1992
rect 20220 1980 20226 2032
rect 23290 1980 23296 2032
rect 23348 2020 23354 2032
rect 45370 2020 45376 2032
rect 23348 1992 45376 2020
rect 23348 1980 23354 1992
rect 45370 1980 45376 1992
rect 45428 1980 45434 2032
rect 46934 1980 46940 2032
rect 46992 2020 46998 2032
rect 52730 2020 52736 2032
rect 46992 1992 52736 2020
rect 46992 1980 46998 1992
rect 52730 1980 52736 1992
rect 52788 1980 52794 2032
rect 4522 1912 4528 1964
rect 4580 1952 4586 1964
rect 25590 1952 25596 1964
rect 4580 1924 25596 1952
rect 4580 1912 4586 1924
rect 25590 1912 25596 1924
rect 25648 1952 25654 1964
rect 30466 1952 30472 1964
rect 25648 1924 30472 1952
rect 25648 1912 25654 1924
rect 30466 1912 30472 1924
rect 30524 1912 30530 1964
rect 41598 1912 41604 1964
rect 41656 1952 41662 1964
rect 41656 1924 45554 1952
rect 41656 1912 41662 1924
rect 7742 1844 7748 1896
rect 7800 1884 7806 1896
rect 12434 1884 12440 1896
rect 7800 1856 12440 1884
rect 7800 1844 7806 1856
rect 12434 1844 12440 1856
rect 12492 1844 12498 1896
rect 12618 1844 12624 1896
rect 12676 1884 12682 1896
rect 18598 1884 18604 1896
rect 12676 1856 18604 1884
rect 12676 1844 12682 1856
rect 18598 1844 18604 1856
rect 18656 1844 18662 1896
rect 23106 1844 23112 1896
rect 23164 1884 23170 1896
rect 41782 1884 41788 1896
rect 23164 1856 41788 1884
rect 23164 1844 23170 1856
rect 41782 1844 41788 1856
rect 41840 1844 41846 1896
rect 45526 1884 45554 1924
rect 49418 1912 49424 1964
rect 49476 1952 49482 1964
rect 56226 1952 56232 1964
rect 49476 1924 56232 1952
rect 49476 1912 49482 1924
rect 56226 1912 56232 1924
rect 56284 1912 56290 1964
rect 54202 1884 54208 1896
rect 45526 1856 54208 1884
rect 54202 1844 54208 1856
rect 54260 1844 54266 1896
rect 3050 1776 3056 1828
rect 3108 1816 3114 1828
rect 8202 1816 8208 1828
rect 3108 1788 8208 1816
rect 3108 1776 3114 1788
rect 8202 1776 8208 1788
rect 8260 1776 8266 1828
rect 10686 1776 10692 1828
rect 10744 1816 10750 1828
rect 24762 1816 24768 1828
rect 10744 1788 24768 1816
rect 10744 1776 10750 1788
rect 24762 1776 24768 1788
rect 24820 1776 24826 1828
rect 26206 1788 47072 1816
rect 6546 1708 6552 1760
rect 6604 1748 6610 1760
rect 18138 1748 18144 1760
rect 6604 1720 18144 1748
rect 6604 1708 6610 1720
rect 18138 1708 18144 1720
rect 18196 1708 18202 1760
rect 22462 1708 22468 1760
rect 22520 1748 22526 1760
rect 26206 1748 26234 1788
rect 22520 1720 26234 1748
rect 22520 1708 22526 1720
rect 40034 1708 40040 1760
rect 40092 1748 40098 1760
rect 43070 1748 43076 1760
rect 40092 1720 43076 1748
rect 40092 1708 40098 1720
rect 43070 1708 43076 1720
rect 43128 1708 43134 1760
rect 44726 1708 44732 1760
rect 44784 1748 44790 1760
rect 46842 1748 46848 1760
rect 44784 1720 46848 1748
rect 44784 1708 44790 1720
rect 46842 1708 46848 1720
rect 46900 1708 46906 1760
rect 47044 1748 47072 1788
rect 47118 1776 47124 1828
rect 47176 1816 47182 1828
rect 55766 1816 55772 1828
rect 47176 1788 55772 1816
rect 47176 1776 47182 1788
rect 55766 1776 55772 1788
rect 55824 1776 55830 1828
rect 54018 1748 54024 1760
rect 47044 1720 54024 1748
rect 54018 1708 54024 1720
rect 54076 1708 54082 1760
rect 12434 1640 12440 1692
rect 12492 1680 12498 1692
rect 21634 1680 21640 1692
rect 12492 1652 21640 1680
rect 12492 1640 12498 1652
rect 21634 1640 21640 1652
rect 21692 1640 21698 1692
rect 23658 1640 23664 1692
rect 23716 1680 23722 1692
rect 44818 1680 44824 1692
rect 23716 1652 44824 1680
rect 23716 1640 23722 1652
rect 44818 1640 44824 1652
rect 44876 1640 44882 1692
rect 7190 1436 7196 1488
rect 7248 1476 7254 1488
rect 7926 1476 7932 1488
rect 7248 1448 7932 1476
rect 7248 1436 7254 1448
rect 7926 1436 7932 1448
rect 7984 1436 7990 1488
rect 7006 1368 7012 1420
rect 7064 1408 7070 1420
rect 7742 1408 7748 1420
rect 7064 1380 7748 1408
rect 7064 1368 7070 1380
rect 7742 1368 7748 1380
rect 7800 1368 7806 1420
rect 9214 1408 9220 1420
rect 8036 1380 9220 1408
rect 8036 1352 8064 1380
rect 9214 1368 9220 1380
rect 9272 1368 9278 1420
rect 25406 1368 25412 1420
rect 25464 1408 25470 1420
rect 27522 1408 27528 1420
rect 25464 1380 27528 1408
rect 25464 1368 25470 1380
rect 27522 1368 27528 1380
rect 27580 1368 27586 1420
rect 35894 1368 35900 1420
rect 35952 1408 35958 1420
rect 37090 1408 37096 1420
rect 35952 1380 37096 1408
rect 35952 1368 35958 1380
rect 37090 1368 37096 1380
rect 37148 1368 37154 1420
rect 38378 1368 38384 1420
rect 38436 1408 38442 1420
rect 39942 1408 39948 1420
rect 38436 1380 39948 1408
rect 38436 1368 38442 1380
rect 39942 1368 39948 1380
rect 40000 1368 40006 1420
rect 48314 1368 48320 1420
rect 48372 1408 48378 1420
rect 49602 1408 49608 1420
rect 48372 1380 49608 1408
rect 48372 1368 48378 1380
rect 49602 1368 49608 1380
rect 49660 1368 49666 1420
rect 8018 1300 8024 1352
rect 8076 1300 8082 1352
<< via1 >>
rect 15398 7590 15450 7642
rect 15462 7590 15514 7642
rect 15526 7590 15578 7642
rect 15590 7590 15642 7642
rect 15654 7590 15706 7642
rect 29846 7590 29898 7642
rect 29910 7590 29962 7642
rect 29974 7590 30026 7642
rect 30038 7590 30090 7642
rect 30102 7590 30154 7642
rect 44294 7590 44346 7642
rect 44358 7590 44410 7642
rect 44422 7590 44474 7642
rect 44486 7590 44538 7642
rect 44550 7590 44602 7642
rect 4436 7352 4488 7404
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 5816 7395 5868 7404
rect 5816 7361 5825 7395
rect 5825 7361 5859 7395
rect 5859 7361 5868 7395
rect 5816 7352 5868 7361
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 7564 7395 7616 7404
rect 7564 7361 7573 7395
rect 7573 7361 7607 7395
rect 7607 7361 7616 7395
rect 7564 7352 7616 7361
rect 8392 7395 8444 7404
rect 8392 7361 8401 7395
rect 8401 7361 8435 7395
rect 8435 7361 8444 7395
rect 8392 7352 8444 7361
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9956 7352 10008 7404
rect 10416 7352 10468 7404
rect 11888 7395 11940 7404
rect 11888 7361 11897 7395
rect 11897 7361 11931 7395
rect 11931 7361 11940 7395
rect 11888 7352 11940 7361
rect 12624 7395 12676 7404
rect 12624 7361 12633 7395
rect 12633 7361 12667 7395
rect 12667 7361 12676 7395
rect 12624 7352 12676 7361
rect 13268 7395 13320 7404
rect 13268 7361 13277 7395
rect 13277 7361 13311 7395
rect 13311 7361 13320 7395
rect 13268 7352 13320 7361
rect 14648 7395 14700 7404
rect 14648 7361 14657 7395
rect 14657 7361 14691 7395
rect 14691 7361 14700 7395
rect 14648 7352 14700 7361
rect 15292 7352 15344 7404
rect 15936 7395 15988 7404
rect 15936 7361 15945 7395
rect 15945 7361 15979 7395
rect 15979 7361 15988 7395
rect 15936 7352 15988 7361
rect 17224 7395 17276 7404
rect 17224 7361 17233 7395
rect 17233 7361 17267 7395
rect 17267 7361 17276 7395
rect 17224 7352 17276 7361
rect 18052 7395 18104 7404
rect 18052 7361 18061 7395
rect 18061 7361 18095 7395
rect 18095 7361 18104 7395
rect 18052 7352 18104 7361
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 19524 7395 19576 7404
rect 19524 7361 19533 7395
rect 19533 7361 19567 7395
rect 19567 7361 19576 7395
rect 19524 7352 19576 7361
rect 20168 7395 20220 7404
rect 20168 7361 20177 7395
rect 20177 7361 20211 7395
rect 20211 7361 20220 7395
rect 20168 7352 20220 7361
rect 21272 7395 21324 7404
rect 21272 7361 21281 7395
rect 21281 7361 21315 7395
rect 21315 7361 21324 7395
rect 21272 7352 21324 7361
rect 22376 7352 22428 7404
rect 22928 7395 22980 7404
rect 22928 7361 22937 7395
rect 22937 7361 22971 7395
rect 22971 7361 22980 7395
rect 22928 7352 22980 7361
rect 23664 7395 23716 7404
rect 23664 7361 23673 7395
rect 23673 7361 23707 7395
rect 23707 7361 23716 7395
rect 23664 7352 23716 7361
rect 25136 7395 25188 7404
rect 25136 7361 25145 7395
rect 25145 7361 25179 7395
rect 25179 7361 25188 7395
rect 25136 7352 25188 7361
rect 25596 7395 25648 7404
rect 25596 7361 25605 7395
rect 25605 7361 25639 7395
rect 25639 7361 25648 7395
rect 25596 7352 25648 7361
rect 26424 7395 26476 7404
rect 26424 7361 26433 7395
rect 26433 7361 26467 7395
rect 26467 7361 26476 7395
rect 26424 7352 26476 7361
rect 27712 7395 27764 7404
rect 27712 7361 27721 7395
rect 27721 7361 27755 7395
rect 27755 7361 27764 7395
rect 27712 7352 27764 7361
rect 28356 7395 28408 7404
rect 28356 7361 28365 7395
rect 28365 7361 28399 7395
rect 28399 7361 28408 7395
rect 28356 7352 28408 7361
rect 29000 7395 29052 7404
rect 29000 7361 29009 7395
rect 29009 7361 29043 7395
rect 29043 7361 29052 7395
rect 29000 7352 29052 7361
rect 29736 7352 29788 7404
rect 30564 7395 30616 7404
rect 30564 7361 30573 7395
rect 30573 7361 30607 7395
rect 30607 7361 30616 7395
rect 30564 7352 30616 7361
rect 31208 7395 31260 7404
rect 31208 7361 31217 7395
rect 31217 7361 31251 7395
rect 31251 7361 31260 7395
rect 31208 7352 31260 7361
rect 32128 7395 32180 7404
rect 32128 7361 32137 7395
rect 32137 7361 32171 7395
rect 32171 7361 32180 7395
rect 32128 7352 32180 7361
rect 32772 7395 32824 7404
rect 32772 7361 32781 7395
rect 32781 7361 32815 7395
rect 32815 7361 32824 7395
rect 32772 7352 32824 7361
rect 33416 7352 33468 7404
rect 33876 7352 33928 7404
rect 34796 7352 34848 7404
rect 36636 7352 36688 7404
rect 37556 7352 37608 7404
rect 38016 7352 38068 7404
rect 38936 7352 38988 7404
rect 40500 7395 40552 7404
rect 40500 7361 40509 7395
rect 40509 7361 40543 7395
rect 40543 7361 40552 7395
rect 40500 7352 40552 7361
rect 41144 7395 41196 7404
rect 41144 7361 41153 7395
rect 41153 7361 41187 7395
rect 41187 7361 41196 7395
rect 41144 7352 41196 7361
rect 41696 7352 41748 7404
rect 43076 7352 43128 7404
rect 44640 7352 44692 7404
rect 45192 7352 45244 7404
rect 45836 7352 45888 7404
rect 47584 7395 47636 7404
rect 47584 7361 47593 7395
rect 47593 7361 47627 7395
rect 47627 7361 47636 7395
rect 47584 7352 47636 7361
rect 47676 7352 47728 7404
rect 48872 7395 48924 7404
rect 48872 7361 48881 7395
rect 48881 7361 48915 7395
rect 48915 7361 48924 7395
rect 48872 7352 48924 7361
rect 50160 7395 50212 7404
rect 50160 7361 50169 7395
rect 50169 7361 50203 7395
rect 50203 7361 50212 7395
rect 50160 7352 50212 7361
rect 50436 7352 50488 7404
rect 51448 7395 51500 7404
rect 51448 7361 51457 7395
rect 51457 7361 51491 7395
rect 51491 7361 51500 7395
rect 51448 7352 51500 7361
rect 52184 7352 52236 7404
rect 53104 7352 53156 7404
rect 53472 7352 53524 7404
rect 55220 7352 55272 7404
rect 55496 7352 55548 7404
rect 56232 7352 56284 7404
rect 35256 7284 35308 7336
rect 42432 7216 42484 7268
rect 8174 7046 8226 7098
rect 8238 7046 8290 7098
rect 8302 7046 8354 7098
rect 8366 7046 8418 7098
rect 8430 7046 8482 7098
rect 22622 7046 22674 7098
rect 22686 7046 22738 7098
rect 22750 7046 22802 7098
rect 22814 7046 22866 7098
rect 22878 7046 22930 7098
rect 37070 7046 37122 7098
rect 37134 7046 37186 7098
rect 37198 7046 37250 7098
rect 37262 7046 37314 7098
rect 37326 7046 37378 7098
rect 51518 7046 51570 7098
rect 51582 7046 51634 7098
rect 51646 7046 51698 7098
rect 51710 7046 51762 7098
rect 51774 7046 51826 7098
rect 6368 6851 6420 6860
rect 6368 6817 6377 6851
rect 6377 6817 6411 6851
rect 6411 6817 6420 6851
rect 6368 6808 6420 6817
rect 11428 6851 11480 6860
rect 11428 6817 11437 6851
rect 11437 6817 11471 6851
rect 11471 6817 11480 6851
rect 11428 6808 11480 6817
rect 14096 6808 14148 6860
rect 16948 6851 17000 6860
rect 16948 6817 16957 6851
rect 16957 6817 16991 6851
rect 16991 6817 17000 6851
rect 16948 6808 17000 6817
rect 20996 6808 21048 6860
rect 24400 6851 24452 6860
rect 24400 6817 24409 6851
rect 24409 6817 24443 6851
rect 24443 6817 24452 6851
rect 24400 6808 24452 6817
rect 26976 6808 27028 6860
rect 36268 6851 36320 6860
rect 36268 6817 36277 6851
rect 36277 6817 36311 6851
rect 36311 6817 36320 6851
rect 36268 6808 36320 6817
rect 39396 6808 39448 6860
rect 43628 6851 43680 6860
rect 43628 6817 43637 6851
rect 43637 6817 43671 6851
rect 43671 6817 43680 6851
rect 43628 6808 43680 6817
rect 46296 6808 46348 6860
rect 49056 6808 49108 6860
rect 54208 6851 54260 6860
rect 54208 6817 54217 6851
rect 54217 6817 54251 6851
rect 54251 6817 54260 6851
rect 54208 6808 54260 6817
rect 27344 6672 27396 6724
rect 47032 6672 47084 6724
rect 48136 6672 48188 6724
rect 9864 6604 9916 6656
rect 33508 6647 33560 6656
rect 33508 6613 33517 6647
rect 33517 6613 33551 6647
rect 33551 6613 33560 6647
rect 33508 6604 33560 6613
rect 52184 6647 52236 6656
rect 52184 6613 52193 6647
rect 52193 6613 52227 6647
rect 52227 6613 52236 6647
rect 52184 6604 52236 6613
rect 15398 6502 15450 6554
rect 15462 6502 15514 6554
rect 15526 6502 15578 6554
rect 15590 6502 15642 6554
rect 15654 6502 15706 6554
rect 29846 6502 29898 6554
rect 29910 6502 29962 6554
rect 29974 6502 30026 6554
rect 30038 6502 30090 6554
rect 30102 6502 30154 6554
rect 44294 6502 44346 6554
rect 44358 6502 44410 6554
rect 44422 6502 44474 6554
rect 44486 6502 44538 6554
rect 44550 6502 44602 6554
rect 8668 6196 8720 6248
rect 20812 6196 20864 6248
rect 30288 6196 30340 6248
rect 9864 6128 9916 6180
rect 8760 6103 8812 6112
rect 8760 6069 8769 6103
rect 8769 6069 8803 6103
rect 8803 6069 8812 6103
rect 8760 6060 8812 6069
rect 9312 6103 9364 6112
rect 9312 6069 9321 6103
rect 9321 6069 9355 6103
rect 9355 6069 9364 6103
rect 9312 6060 9364 6069
rect 9496 6060 9548 6112
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 20720 6060 20772 6112
rect 23296 6103 23348 6112
rect 23296 6069 23305 6103
rect 23305 6069 23339 6103
rect 23339 6069 23348 6103
rect 23296 6060 23348 6069
rect 25136 6060 25188 6112
rect 26976 6103 27028 6112
rect 26976 6069 26985 6103
rect 26985 6069 27019 6103
rect 27019 6069 27028 6103
rect 26976 6060 27028 6069
rect 28264 6060 28316 6112
rect 30472 6103 30524 6112
rect 30472 6069 30481 6103
rect 30481 6069 30515 6103
rect 30515 6069 30524 6103
rect 30472 6060 30524 6069
rect 31760 6060 31812 6112
rect 33232 6103 33284 6112
rect 33232 6069 33241 6103
rect 33241 6069 33275 6103
rect 33275 6069 33284 6103
rect 33232 6060 33284 6069
rect 38384 6196 38436 6248
rect 42984 6196 43036 6248
rect 33508 6128 33560 6180
rect 40040 6128 40092 6180
rect 50896 6128 50948 6180
rect 34612 6103 34664 6112
rect 34612 6069 34621 6103
rect 34621 6069 34655 6103
rect 34655 6069 34664 6103
rect 34612 6060 34664 6069
rect 35072 6103 35124 6112
rect 35072 6069 35081 6103
rect 35081 6069 35115 6103
rect 35115 6069 35124 6103
rect 35072 6060 35124 6069
rect 35716 6103 35768 6112
rect 35716 6069 35725 6103
rect 35725 6069 35759 6103
rect 35759 6069 35768 6103
rect 35716 6060 35768 6069
rect 35808 6060 35860 6112
rect 36268 6060 36320 6112
rect 39764 6060 39816 6112
rect 45560 6103 45612 6112
rect 45560 6069 45569 6103
rect 45569 6069 45603 6103
rect 45603 6069 45612 6103
rect 45560 6060 45612 6069
rect 46940 6060 46992 6112
rect 51356 6060 51408 6112
rect 52000 6060 52052 6112
rect 8174 5958 8226 6010
rect 8238 5958 8290 6010
rect 8302 5958 8354 6010
rect 8366 5958 8418 6010
rect 8430 5958 8482 6010
rect 22622 5958 22674 6010
rect 22686 5958 22738 6010
rect 22750 5958 22802 6010
rect 22814 5958 22866 6010
rect 22878 5958 22930 6010
rect 37070 5958 37122 6010
rect 37134 5958 37186 6010
rect 37198 5958 37250 6010
rect 37262 5958 37314 6010
rect 37326 5958 37378 6010
rect 51518 5958 51570 6010
rect 51582 5958 51634 6010
rect 51646 5958 51698 6010
rect 51710 5958 51762 6010
rect 51774 5958 51826 6010
rect 5448 5856 5500 5908
rect 10508 5856 10560 5908
rect 20812 5856 20864 5908
rect 31852 5856 31904 5908
rect 33048 5856 33100 5908
rect 34704 5899 34756 5908
rect 34704 5865 34713 5899
rect 34713 5865 34747 5899
rect 34747 5865 34756 5899
rect 34704 5856 34756 5865
rect 35532 5856 35584 5908
rect 35716 5856 35768 5908
rect 41696 5856 41748 5908
rect 42984 5856 43036 5908
rect 49792 5856 49844 5908
rect 52184 5856 52236 5908
rect 4344 5788 4396 5840
rect 7840 5720 7892 5772
rect 8024 5652 8076 5704
rect 9312 5652 9364 5704
rect 10048 5652 10100 5704
rect 10876 5652 10928 5704
rect 12072 5695 12124 5704
rect 12072 5661 12081 5695
rect 12081 5661 12115 5695
rect 12115 5661 12124 5695
rect 12072 5652 12124 5661
rect 4160 5584 4212 5636
rect 9864 5584 9916 5636
rect 27712 5788 27764 5840
rect 27620 5720 27672 5772
rect 31024 5831 31076 5840
rect 31024 5797 31033 5831
rect 31033 5797 31067 5831
rect 31067 5797 31076 5831
rect 31024 5788 31076 5797
rect 34612 5788 34664 5840
rect 48136 5831 48188 5840
rect 31668 5763 31720 5772
rect 12808 5652 12860 5704
rect 14740 5652 14792 5704
rect 16212 5652 16264 5704
rect 16948 5652 17000 5704
rect 26792 5652 26844 5704
rect 29736 5652 29788 5704
rect 22744 5584 22796 5636
rect 31668 5729 31677 5763
rect 31677 5729 31711 5763
rect 31711 5729 31720 5763
rect 31668 5720 31720 5729
rect 7748 5516 7800 5568
rect 12900 5516 12952 5568
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 16304 5559 16356 5568
rect 16304 5525 16313 5559
rect 16313 5525 16347 5559
rect 16347 5525 16356 5559
rect 16304 5516 16356 5525
rect 19984 5516 20036 5568
rect 20720 5559 20772 5568
rect 20720 5525 20729 5559
rect 20729 5525 20763 5559
rect 20763 5525 20772 5559
rect 20720 5516 20772 5525
rect 21640 5516 21692 5568
rect 22468 5516 22520 5568
rect 23020 5516 23072 5568
rect 23480 5559 23532 5568
rect 23480 5525 23489 5559
rect 23489 5525 23523 5559
rect 23523 5525 23532 5559
rect 23480 5516 23532 5525
rect 24768 5516 24820 5568
rect 25136 5559 25188 5568
rect 25136 5525 25145 5559
rect 25145 5525 25179 5559
rect 25179 5525 25188 5559
rect 25136 5516 25188 5525
rect 25228 5516 25280 5568
rect 26700 5516 26752 5568
rect 26884 5516 26936 5568
rect 28816 5559 28868 5568
rect 28816 5525 28825 5559
rect 28825 5525 28859 5559
rect 28859 5525 28868 5559
rect 28816 5516 28868 5525
rect 29460 5516 29512 5568
rect 30380 5559 30432 5568
rect 30380 5525 30389 5559
rect 30389 5525 30423 5559
rect 30423 5525 30432 5559
rect 30380 5516 30432 5525
rect 31852 5584 31904 5636
rect 32128 5627 32180 5636
rect 32128 5593 32137 5627
rect 32137 5593 32171 5627
rect 32171 5593 32180 5627
rect 32128 5584 32180 5593
rect 33048 5720 33100 5772
rect 34888 5763 34940 5772
rect 34888 5729 34897 5763
rect 34897 5729 34931 5763
rect 34931 5729 34940 5763
rect 34888 5720 34940 5729
rect 32864 5652 32916 5704
rect 34152 5652 34204 5704
rect 35808 5720 35860 5772
rect 32036 5516 32088 5568
rect 33416 5559 33468 5568
rect 33416 5525 33425 5559
rect 33425 5525 33459 5559
rect 33459 5525 33468 5559
rect 33416 5516 33468 5525
rect 35532 5652 35584 5704
rect 36268 5695 36320 5704
rect 36268 5661 36277 5695
rect 36277 5661 36311 5695
rect 36311 5661 36320 5695
rect 36268 5652 36320 5661
rect 36452 5695 36504 5704
rect 36452 5661 36461 5695
rect 36461 5661 36495 5695
rect 36495 5661 36504 5695
rect 36452 5652 36504 5661
rect 40132 5720 40184 5772
rect 48136 5797 48145 5831
rect 48145 5797 48179 5831
rect 48179 5797 48188 5831
rect 48136 5788 48188 5797
rect 35348 5584 35400 5636
rect 42800 5652 42852 5704
rect 52276 5720 52328 5772
rect 39856 5584 39908 5636
rect 40040 5584 40092 5636
rect 40500 5584 40552 5636
rect 45560 5652 45612 5704
rect 50252 5652 50304 5704
rect 50528 5652 50580 5704
rect 51448 5652 51500 5704
rect 51908 5652 51960 5704
rect 43076 5516 43128 5568
rect 45192 5516 45244 5568
rect 46020 5516 46072 5568
rect 49700 5584 49752 5636
rect 54760 5584 54812 5636
rect 46940 5516 46992 5568
rect 49792 5516 49844 5568
rect 55220 5516 55272 5568
rect 15398 5414 15450 5466
rect 15462 5414 15514 5466
rect 15526 5414 15578 5466
rect 15590 5414 15642 5466
rect 15654 5414 15706 5466
rect 29846 5414 29898 5466
rect 29910 5414 29962 5466
rect 29974 5414 30026 5466
rect 30038 5414 30090 5466
rect 30102 5414 30154 5466
rect 44294 5414 44346 5466
rect 44358 5414 44410 5466
rect 44422 5414 44474 5466
rect 44486 5414 44538 5466
rect 44550 5414 44602 5466
rect 4344 5355 4396 5364
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 5448 5312 5500 5364
rect 9864 5312 9916 5364
rect 19248 5312 19300 5364
rect 20720 5355 20772 5364
rect 20720 5321 20729 5355
rect 20729 5321 20763 5355
rect 20763 5321 20772 5355
rect 20720 5312 20772 5321
rect 24124 5312 24176 5364
rect 25136 5312 25188 5364
rect 25780 5312 25832 5364
rect 29552 5312 29604 5364
rect 31024 5312 31076 5364
rect 6276 5244 6328 5296
rect 6552 5244 6604 5296
rect 12716 5244 12768 5296
rect 13452 5287 13504 5296
rect 13452 5253 13461 5287
rect 13461 5253 13495 5287
rect 13495 5253 13504 5287
rect 13452 5244 13504 5253
rect 18328 5244 18380 5296
rect 20812 5244 20864 5296
rect 21180 5287 21232 5296
rect 21180 5253 21189 5287
rect 21189 5253 21223 5287
rect 21223 5253 21232 5287
rect 21180 5244 21232 5253
rect 22744 5287 22796 5296
rect 22744 5253 22753 5287
rect 22753 5253 22787 5287
rect 22787 5253 22796 5287
rect 22744 5244 22796 5253
rect 23388 5244 23440 5296
rect 25228 5244 25280 5296
rect 4620 5176 4672 5228
rect 5172 5219 5224 5228
rect 5172 5185 5181 5219
rect 5181 5185 5215 5219
rect 5215 5185 5224 5219
rect 5172 5176 5224 5185
rect 4068 5151 4120 5160
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 4068 5108 4120 5117
rect 4436 5108 4488 5160
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 7012 5176 7064 5228
rect 7840 5176 7892 5228
rect 8668 5176 8720 5228
rect 8760 5176 8812 5228
rect 9220 5176 9272 5228
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 11796 5176 11848 5228
rect 16764 5176 16816 5228
rect 17960 5176 18012 5228
rect 3424 4972 3476 5024
rect 7196 5040 7248 5092
rect 12348 5108 12400 5160
rect 12624 5151 12676 5160
rect 12624 5117 12633 5151
rect 12633 5117 12667 5151
rect 12667 5117 12676 5151
rect 12624 5108 12676 5117
rect 16488 5108 16540 5160
rect 25320 5176 25372 5228
rect 28172 5244 28224 5296
rect 26976 5219 27028 5228
rect 26976 5185 26985 5219
rect 26985 5185 27019 5219
rect 27019 5185 27028 5219
rect 26976 5176 27028 5185
rect 22192 5108 22244 5160
rect 24768 5108 24820 5160
rect 25044 5108 25096 5160
rect 31668 5176 31720 5228
rect 32128 5219 32180 5228
rect 32128 5185 32137 5219
rect 32137 5185 32171 5219
rect 32171 5185 32180 5219
rect 32128 5176 32180 5185
rect 33416 5244 33468 5296
rect 41696 5355 41748 5364
rect 33232 5176 33284 5228
rect 33876 5176 33928 5228
rect 34152 5219 34204 5228
rect 34152 5185 34161 5219
rect 34161 5185 34195 5219
rect 34195 5185 34204 5219
rect 34152 5176 34204 5185
rect 35348 5176 35400 5228
rect 36728 5219 36780 5228
rect 36728 5185 36737 5219
rect 36737 5185 36771 5219
rect 36771 5185 36780 5219
rect 36728 5176 36780 5185
rect 38660 5176 38712 5228
rect 38752 5176 38804 5228
rect 39488 5219 39540 5228
rect 39488 5185 39497 5219
rect 39497 5185 39531 5219
rect 39531 5185 39540 5219
rect 41696 5321 41705 5355
rect 41705 5321 41739 5355
rect 41739 5321 41748 5355
rect 41696 5312 41748 5321
rect 42616 5355 42668 5364
rect 42616 5321 42625 5355
rect 42625 5321 42659 5355
rect 42659 5321 42668 5355
rect 42616 5312 42668 5321
rect 39488 5176 39540 5185
rect 29460 5108 29512 5160
rect 30288 5108 30340 5160
rect 32864 5108 32916 5160
rect 33968 5151 34020 5160
rect 33968 5117 33977 5151
rect 33977 5117 34011 5151
rect 34011 5117 34020 5151
rect 33968 5108 34020 5117
rect 12440 5040 12492 5092
rect 16028 5040 16080 5092
rect 17592 5040 17644 5092
rect 19156 5040 19208 5092
rect 24584 5040 24636 5092
rect 29736 5040 29788 5092
rect 4712 4972 4764 5024
rect 7104 5015 7156 5024
rect 7104 4981 7113 5015
rect 7113 4981 7147 5015
rect 7147 4981 7156 5015
rect 7104 4972 7156 4981
rect 10232 4972 10284 5024
rect 10600 4972 10652 5024
rect 10968 5015 11020 5024
rect 10968 4981 10977 5015
rect 10977 4981 11011 5015
rect 11011 4981 11020 5015
rect 10968 4972 11020 4981
rect 14464 4972 14516 5024
rect 15016 4972 15068 5024
rect 15752 4972 15804 5024
rect 16764 5015 16816 5024
rect 16764 4981 16773 5015
rect 16773 4981 16807 5015
rect 16807 4981 16816 5015
rect 16764 4972 16816 4981
rect 17132 4972 17184 5024
rect 18972 5015 19024 5024
rect 18972 4981 18981 5015
rect 18981 4981 19015 5015
rect 19015 4981 19024 5015
rect 18972 4972 19024 4981
rect 19892 4972 19944 5024
rect 22100 4972 22152 5024
rect 23020 4972 23072 5024
rect 23848 4972 23900 5024
rect 24952 5015 25004 5024
rect 24952 4981 24961 5015
rect 24961 4981 24995 5015
rect 24995 4981 25004 5015
rect 24952 4972 25004 4981
rect 27160 4972 27212 5024
rect 28448 4972 28500 5024
rect 31668 4972 31720 5024
rect 34888 5108 34940 5160
rect 35808 5151 35860 5160
rect 35808 5117 35817 5151
rect 35817 5117 35851 5151
rect 35851 5117 35860 5151
rect 35808 5108 35860 5117
rect 42432 5244 42484 5296
rect 40132 5219 40184 5228
rect 40132 5185 40178 5219
rect 40178 5185 40184 5219
rect 40500 5219 40552 5228
rect 40132 5176 40184 5185
rect 40500 5185 40509 5219
rect 40509 5185 40543 5219
rect 40543 5185 40552 5219
rect 40500 5176 40552 5185
rect 41052 5219 41104 5228
rect 41052 5185 41061 5219
rect 41061 5185 41095 5219
rect 41095 5185 41104 5219
rect 41052 5176 41104 5185
rect 41236 5219 41288 5228
rect 41236 5185 41245 5219
rect 41245 5185 41279 5219
rect 41279 5185 41288 5219
rect 43444 5219 43496 5228
rect 41236 5176 41288 5185
rect 43444 5185 43453 5219
rect 43453 5185 43487 5219
rect 43487 5185 43496 5219
rect 43444 5176 43496 5185
rect 44548 5219 44600 5228
rect 44548 5185 44557 5219
rect 44557 5185 44591 5219
rect 44591 5185 44600 5219
rect 44548 5176 44600 5185
rect 44732 5219 44784 5228
rect 44732 5185 44741 5219
rect 44741 5185 44775 5219
rect 44775 5185 44784 5219
rect 44732 5176 44784 5185
rect 45192 5219 45244 5228
rect 45192 5185 45201 5219
rect 45201 5185 45235 5219
rect 45235 5185 45244 5219
rect 45192 5176 45244 5185
rect 54024 5312 54076 5364
rect 48320 5287 48372 5296
rect 48320 5253 48329 5287
rect 48329 5253 48363 5287
rect 48363 5253 48372 5287
rect 48320 5244 48372 5253
rect 51172 5244 51224 5296
rect 46388 5176 46440 5228
rect 40684 5108 40736 5160
rect 42800 5151 42852 5160
rect 42800 5117 42809 5151
rect 42809 5117 42843 5151
rect 42843 5117 42852 5151
rect 42800 5108 42852 5117
rect 34336 5015 34388 5024
rect 34336 4981 34345 5015
rect 34345 4981 34379 5015
rect 34379 4981 34388 5015
rect 34336 4972 34388 4981
rect 35440 4972 35492 5024
rect 37556 5015 37608 5024
rect 37556 4981 37565 5015
rect 37565 4981 37599 5015
rect 37599 4981 37608 5015
rect 37556 4972 37608 4981
rect 38200 5015 38252 5024
rect 38200 4981 38209 5015
rect 38209 4981 38243 5015
rect 38243 4981 38252 5015
rect 38200 4972 38252 4981
rect 40224 5083 40276 5092
rect 40224 5049 40233 5083
rect 40233 5049 40267 5083
rect 40267 5049 40276 5083
rect 40224 5040 40276 5049
rect 39212 4972 39264 5024
rect 39764 4972 39816 5024
rect 42432 4972 42484 5024
rect 44548 5040 44600 5092
rect 43444 5015 43496 5024
rect 43444 4981 43453 5015
rect 43453 4981 43487 5015
rect 43487 4981 43496 5015
rect 43444 4972 43496 4981
rect 44640 4972 44692 5024
rect 50896 5219 50948 5228
rect 50896 5185 50905 5219
rect 50905 5185 50939 5219
rect 50939 5185 50948 5219
rect 50896 5176 50948 5185
rect 55404 5244 55456 5296
rect 52000 5219 52052 5228
rect 52000 5185 52009 5219
rect 52009 5185 52043 5219
rect 52043 5185 52052 5219
rect 52000 5176 52052 5185
rect 45376 5040 45428 5092
rect 47124 5040 47176 5092
rect 49332 5108 49384 5160
rect 51264 5108 51316 5160
rect 55680 5176 55732 5228
rect 55588 5108 55640 5160
rect 46296 4972 46348 5024
rect 46756 4972 46808 5024
rect 50160 5040 50212 5092
rect 52552 5040 52604 5092
rect 52736 5040 52788 5092
rect 49608 4972 49660 5024
rect 52644 4972 52696 5024
rect 52828 5015 52880 5024
rect 52828 4981 52837 5015
rect 52837 4981 52871 5015
rect 52871 4981 52880 5015
rect 52828 4972 52880 4981
rect 53012 4972 53064 5024
rect 55312 5015 55364 5024
rect 55312 4981 55321 5015
rect 55321 4981 55355 5015
rect 55355 4981 55364 5015
rect 55312 4972 55364 4981
rect 55772 5015 55824 5024
rect 55772 4981 55781 5015
rect 55781 4981 55815 5015
rect 55815 4981 55824 5015
rect 55772 4972 55824 4981
rect 8174 4870 8226 4922
rect 8238 4870 8290 4922
rect 8302 4870 8354 4922
rect 8366 4870 8418 4922
rect 8430 4870 8482 4922
rect 22622 4870 22674 4922
rect 22686 4870 22738 4922
rect 22750 4870 22802 4922
rect 22814 4870 22866 4922
rect 22878 4870 22930 4922
rect 37070 4870 37122 4922
rect 37134 4870 37186 4922
rect 37198 4870 37250 4922
rect 37262 4870 37314 4922
rect 37326 4870 37378 4922
rect 51518 4870 51570 4922
rect 51582 4870 51634 4922
rect 51646 4870 51698 4922
rect 51710 4870 51762 4922
rect 51774 4870 51826 4922
rect 4252 4768 4304 4820
rect 4620 4768 4672 4820
rect 11704 4768 11756 4820
rect 13084 4768 13136 4820
rect 18144 4811 18196 4820
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 18972 4768 19024 4820
rect 10324 4700 10376 4752
rect 11796 4743 11848 4752
rect 11796 4709 11805 4743
rect 11805 4709 11839 4743
rect 11839 4709 11848 4743
rect 11796 4700 11848 4709
rect 12992 4700 13044 4752
rect 16120 4700 16172 4752
rect 8300 4632 8352 4684
rect 9404 4632 9456 4684
rect 9864 4632 9916 4684
rect 13176 4632 13228 4684
rect 16672 4632 16724 4684
rect 17408 4632 17460 4684
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3792 4607 3844 4616
rect 3240 4564 3292 4573
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 4160 4564 4212 4616
rect 4712 4607 4764 4616
rect 4712 4573 4746 4607
rect 4746 4573 4764 4607
rect 4712 4564 4764 4573
rect 5816 4564 5868 4616
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7104 4564 7156 4616
rect 7748 4607 7800 4616
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 9956 4607 10008 4616
rect 9956 4573 9965 4607
rect 9965 4573 9999 4607
rect 9999 4573 10008 4607
rect 9956 4564 10008 4573
rect 10232 4564 10284 4616
rect 4068 4496 4120 4548
rect 6276 4539 6328 4548
rect 6276 4505 6285 4539
rect 6285 4505 6319 4539
rect 6319 4505 6328 4539
rect 6276 4496 6328 4505
rect 4252 4428 4304 4480
rect 5172 4428 5224 4480
rect 9680 4496 9732 4548
rect 11520 4496 11572 4548
rect 7288 4428 7340 4480
rect 7656 4471 7708 4480
rect 7656 4437 7665 4471
rect 7665 4437 7699 4471
rect 7699 4437 7708 4471
rect 7656 4428 7708 4437
rect 9588 4428 9640 4480
rect 11980 4428 12032 4480
rect 12716 4607 12768 4616
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 14188 4564 14240 4616
rect 14372 4564 14424 4616
rect 12624 4496 12676 4548
rect 15384 4564 15436 4616
rect 17592 4607 17644 4616
rect 17592 4573 17601 4607
rect 17601 4573 17635 4607
rect 17635 4573 17644 4607
rect 17592 4564 17644 4573
rect 18052 4700 18104 4752
rect 18328 4675 18380 4684
rect 15844 4496 15896 4548
rect 16120 4496 16172 4548
rect 18328 4641 18337 4675
rect 18337 4641 18371 4675
rect 18371 4641 18380 4675
rect 18328 4632 18380 4641
rect 18420 4607 18472 4616
rect 18420 4573 18429 4607
rect 18429 4573 18463 4607
rect 18463 4573 18472 4607
rect 18420 4564 18472 4573
rect 22100 4700 22152 4752
rect 19248 4675 19300 4684
rect 19248 4641 19257 4675
rect 19257 4641 19291 4675
rect 19291 4641 19300 4675
rect 19248 4632 19300 4641
rect 21272 4564 21324 4616
rect 17960 4496 18012 4548
rect 22560 4607 22612 4616
rect 22560 4573 22569 4607
rect 22569 4573 22603 4607
rect 22603 4573 22612 4607
rect 22560 4564 22612 4573
rect 22744 4607 22796 4616
rect 22744 4573 22753 4607
rect 22753 4573 22787 4607
rect 22787 4573 22796 4607
rect 23388 4700 23440 4752
rect 25044 4743 25096 4752
rect 25044 4709 25053 4743
rect 25053 4709 25087 4743
rect 25087 4709 25096 4743
rect 25044 4700 25096 4709
rect 22744 4564 22796 4573
rect 24216 4564 24268 4616
rect 25136 4632 25188 4684
rect 26884 4632 26936 4684
rect 30288 4768 30340 4820
rect 29460 4700 29512 4752
rect 32128 4700 32180 4752
rect 29552 4675 29604 4684
rect 24584 4607 24636 4616
rect 24584 4573 24593 4607
rect 24593 4573 24627 4607
rect 24627 4573 24636 4607
rect 24584 4564 24636 4573
rect 12716 4428 12768 4480
rect 15200 4428 15252 4480
rect 15936 4471 15988 4480
rect 15936 4437 15945 4471
rect 15945 4437 15979 4471
rect 15979 4437 15988 4471
rect 15936 4428 15988 4437
rect 25780 4564 25832 4616
rect 28264 4607 28316 4616
rect 28264 4573 28273 4607
rect 28273 4573 28307 4607
rect 28307 4573 28316 4607
rect 28264 4564 28316 4573
rect 29552 4641 29561 4675
rect 29561 4641 29595 4675
rect 29595 4641 29604 4675
rect 29552 4632 29604 4641
rect 35624 4768 35676 4820
rect 35808 4768 35860 4820
rect 38752 4768 38804 4820
rect 39488 4768 39540 4820
rect 41236 4768 41288 4820
rect 38660 4700 38712 4752
rect 39120 4700 39172 4752
rect 39212 4700 39264 4752
rect 42432 4768 42484 4820
rect 43444 4768 43496 4820
rect 44364 4768 44416 4820
rect 48320 4768 48372 4820
rect 51172 4811 51224 4820
rect 51172 4777 51181 4811
rect 51181 4777 51215 4811
rect 51215 4777 51224 4811
rect 51172 4768 51224 4777
rect 52460 4768 52512 4820
rect 55680 4811 55732 4820
rect 42892 4700 42944 4752
rect 48596 4743 48648 4752
rect 48596 4709 48605 4743
rect 48605 4709 48639 4743
rect 48639 4709 48648 4743
rect 48596 4700 48648 4709
rect 49608 4700 49660 4752
rect 35440 4675 35492 4684
rect 35440 4641 35449 4675
rect 35449 4641 35483 4675
rect 35483 4641 35492 4675
rect 35440 4632 35492 4641
rect 38752 4632 38804 4684
rect 41052 4632 41104 4684
rect 41788 4632 41840 4684
rect 46020 4675 46072 4684
rect 46020 4641 46029 4675
rect 46029 4641 46063 4675
rect 46063 4641 46072 4675
rect 46020 4632 46072 4641
rect 46296 4675 46348 4684
rect 46296 4641 46305 4675
rect 46305 4641 46339 4675
rect 46339 4641 46348 4675
rect 46296 4632 46348 4641
rect 46388 4632 46440 4684
rect 28724 4564 28776 4616
rect 30656 4564 30708 4616
rect 31392 4564 31444 4616
rect 33876 4607 33928 4616
rect 33876 4573 33885 4607
rect 33885 4573 33919 4607
rect 33919 4573 33928 4607
rect 33876 4564 33928 4573
rect 35072 4564 35124 4616
rect 26148 4428 26200 4480
rect 34428 4496 34480 4548
rect 37556 4564 37608 4616
rect 37648 4607 37700 4616
rect 37648 4573 37657 4607
rect 37657 4573 37691 4607
rect 37691 4573 37700 4607
rect 38384 4607 38436 4616
rect 37648 4564 37700 4573
rect 38384 4573 38393 4607
rect 38393 4573 38427 4607
rect 38427 4573 38436 4607
rect 38384 4564 38436 4573
rect 35716 4496 35768 4548
rect 32588 4428 32640 4480
rect 35808 4428 35860 4480
rect 43352 4564 43404 4616
rect 44364 4564 44416 4616
rect 44640 4564 44692 4616
rect 45192 4607 45244 4616
rect 45192 4573 45201 4607
rect 45201 4573 45235 4607
rect 45235 4573 45244 4607
rect 45192 4564 45244 4573
rect 49608 4607 49660 4616
rect 49608 4573 49617 4607
rect 49617 4573 49651 4607
rect 49651 4573 49660 4607
rect 49608 4564 49660 4573
rect 50160 4607 50212 4616
rect 50160 4573 50169 4607
rect 50169 4573 50203 4607
rect 50203 4573 50212 4607
rect 50160 4564 50212 4573
rect 55680 4777 55689 4811
rect 55689 4777 55723 4811
rect 55723 4777 55732 4811
rect 55680 4768 55732 4777
rect 53748 4675 53800 4684
rect 53748 4641 53757 4675
rect 53757 4641 53791 4675
rect 53791 4641 53800 4675
rect 53748 4632 53800 4641
rect 54024 4607 54076 4616
rect 38936 4471 38988 4480
rect 38936 4437 38945 4471
rect 38945 4437 38979 4471
rect 38979 4437 38988 4471
rect 38936 4428 38988 4437
rect 40592 4471 40644 4480
rect 40592 4437 40601 4471
rect 40601 4437 40635 4471
rect 40635 4437 40644 4471
rect 40592 4428 40644 4437
rect 49884 4496 49936 4548
rect 45560 4428 45612 4480
rect 50896 4428 50948 4480
rect 52092 4471 52144 4480
rect 52092 4437 52101 4471
rect 52101 4437 52135 4471
rect 52135 4437 52144 4471
rect 52092 4428 52144 4437
rect 54024 4573 54033 4607
rect 54033 4573 54067 4607
rect 54067 4573 54076 4607
rect 54024 4564 54076 4573
rect 55496 4607 55548 4616
rect 55496 4573 55505 4607
rect 55505 4573 55539 4607
rect 55539 4573 55548 4607
rect 55496 4564 55548 4573
rect 54760 4471 54812 4480
rect 54760 4437 54769 4471
rect 54769 4437 54803 4471
rect 54803 4437 54812 4471
rect 54760 4428 54812 4437
rect 56600 4428 56652 4480
rect 57244 4471 57296 4480
rect 57244 4437 57253 4471
rect 57253 4437 57287 4471
rect 57287 4437 57296 4471
rect 57244 4428 57296 4437
rect 15398 4326 15450 4378
rect 15462 4326 15514 4378
rect 15526 4326 15578 4378
rect 15590 4326 15642 4378
rect 15654 4326 15706 4378
rect 29846 4326 29898 4378
rect 29910 4326 29962 4378
rect 29974 4326 30026 4378
rect 30038 4326 30090 4378
rect 30102 4326 30154 4378
rect 44294 4326 44346 4378
rect 44358 4326 44410 4378
rect 44422 4326 44474 4378
rect 44486 4326 44538 4378
rect 44550 4326 44602 4378
rect 3792 4224 3844 4276
rect 9956 4224 10008 4276
rect 3148 4156 3200 4208
rect 3240 4156 3292 4208
rect 15292 4224 15344 4276
rect 15384 4224 15436 4276
rect 15936 4224 15988 4276
rect 13544 4156 13596 4208
rect 17960 4224 18012 4276
rect 19248 4224 19300 4276
rect 3424 4131 3476 4140
rect 3424 4097 3433 4131
rect 3433 4097 3467 4131
rect 3467 4097 3476 4131
rect 3424 4088 3476 4097
rect 3792 4088 3844 4140
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 4252 4088 4304 4140
rect 7288 4088 7340 4140
rect 9128 4088 9180 4140
rect 9588 4131 9640 4140
rect 9588 4097 9606 4131
rect 9606 4097 9640 4131
rect 9864 4131 9916 4140
rect 9588 4088 9640 4097
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 10784 4131 10836 4140
rect 10784 4097 10793 4131
rect 10793 4097 10827 4131
rect 10827 4097 10836 4131
rect 10784 4088 10836 4097
rect 11796 4131 11848 4140
rect 11796 4097 11805 4131
rect 11805 4097 11839 4131
rect 11839 4097 11848 4131
rect 11796 4088 11848 4097
rect 8760 4020 8812 4072
rect 10508 4020 10560 4072
rect 11520 4063 11572 4072
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 11704 4020 11756 4072
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 12164 4131 12216 4140
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 12624 4088 12676 4140
rect 8852 3952 8904 4004
rect 11060 3952 11112 4004
rect 13176 4131 13228 4140
rect 13176 4097 13185 4131
rect 13185 4097 13219 4131
rect 13219 4097 13228 4131
rect 13176 4088 13228 4097
rect 15108 4131 15160 4140
rect 15108 4097 15117 4131
rect 15117 4097 15151 4131
rect 15151 4097 15160 4131
rect 15108 4088 15160 4097
rect 15292 4088 15344 4140
rect 15568 4088 15620 4140
rect 16120 4088 16172 4140
rect 16488 4088 16540 4140
rect 13728 4020 13780 4072
rect 16396 4020 16448 4072
rect 18420 4088 18472 4140
rect 19340 4156 19392 4208
rect 22744 4224 22796 4276
rect 30656 4224 30708 4276
rect 31760 4224 31812 4276
rect 32588 4224 32640 4276
rect 34336 4224 34388 4276
rect 23480 4156 23532 4208
rect 28816 4156 28868 4208
rect 31392 4156 31444 4208
rect 35808 4156 35860 4208
rect 39764 4224 39816 4276
rect 44640 4224 44692 4276
rect 49608 4224 49660 4276
rect 52460 4224 52512 4276
rect 52644 4224 52696 4276
rect 49056 4199 49108 4208
rect 21180 4088 21232 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 17960 4063 18012 4072
rect 17960 4029 17969 4063
rect 17969 4029 18003 4063
rect 18003 4029 18012 4063
rect 17960 4020 18012 4029
rect 18328 4020 18380 4072
rect 19064 4063 19116 4072
rect 19064 4029 19073 4063
rect 19073 4029 19107 4063
rect 19107 4029 19116 4063
rect 19064 4020 19116 4029
rect 20720 4020 20772 4072
rect 22192 4131 22244 4140
rect 22192 4097 22201 4131
rect 22201 4097 22235 4131
rect 22235 4097 22244 4131
rect 22192 4088 22244 4097
rect 23848 4088 23900 4140
rect 24124 4131 24176 4140
rect 24124 4097 24133 4131
rect 24133 4097 24167 4131
rect 24167 4097 24176 4131
rect 24124 4088 24176 4097
rect 26332 4088 26384 4140
rect 30932 4088 30984 4140
rect 32588 4131 32640 4140
rect 32588 4097 32597 4131
rect 32597 4097 32631 4131
rect 32631 4097 32640 4131
rect 32588 4088 32640 4097
rect 33416 4131 33468 4140
rect 33416 4097 33425 4131
rect 33425 4097 33459 4131
rect 33459 4097 33468 4131
rect 33416 4088 33468 4097
rect 37556 4088 37608 4140
rect 39120 4131 39172 4140
rect 39120 4097 39129 4131
rect 39129 4097 39163 4131
rect 39163 4097 39172 4131
rect 39120 4088 39172 4097
rect 41696 4131 41748 4140
rect 41696 4097 41705 4131
rect 41705 4097 41739 4131
rect 41739 4097 41748 4131
rect 41696 4088 41748 4097
rect 42984 4088 43036 4140
rect 49056 4165 49065 4199
rect 49065 4165 49099 4199
rect 49099 4165 49108 4199
rect 49056 4156 49108 4165
rect 53012 4199 53064 4208
rect 53012 4165 53021 4199
rect 53021 4165 53055 4199
rect 53055 4165 53064 4199
rect 53012 4156 53064 4165
rect 53656 4224 53708 4276
rect 54760 4224 54812 4276
rect 45744 4131 45796 4140
rect 3056 3884 3108 3936
rect 4160 3884 4212 3936
rect 8392 3884 8444 3936
rect 8944 3884 8996 3936
rect 9220 3884 9272 3936
rect 9588 3884 9640 3936
rect 10968 3884 11020 3936
rect 11428 3884 11480 3936
rect 12624 3884 12676 3936
rect 12992 3884 13044 3936
rect 13084 3927 13136 3936
rect 13084 3893 13093 3927
rect 13093 3893 13127 3927
rect 13127 3893 13136 3927
rect 13084 3884 13136 3893
rect 13360 3884 13412 3936
rect 15108 3884 15160 3936
rect 17868 3884 17920 3936
rect 17960 3884 18012 3936
rect 18236 3884 18288 3936
rect 22560 3952 22612 4004
rect 21088 3884 21140 3936
rect 21824 3884 21876 3936
rect 23204 3884 23256 3936
rect 24308 3884 24360 3936
rect 30380 4020 30432 4072
rect 25504 3995 25556 4004
rect 25504 3961 25513 3995
rect 25513 3961 25547 3995
rect 25547 3961 25556 3995
rect 25504 3952 25556 3961
rect 29736 3952 29788 4004
rect 35900 4020 35952 4072
rect 32772 3995 32824 4004
rect 32772 3961 32781 3995
rect 32781 3961 32815 3995
rect 32815 3961 32824 3995
rect 32772 3952 32824 3961
rect 35624 3952 35676 4004
rect 37464 3952 37516 4004
rect 40132 4020 40184 4072
rect 45744 4097 45753 4131
rect 45753 4097 45787 4131
rect 45787 4097 45796 4131
rect 45744 4088 45796 4097
rect 26424 3927 26476 3936
rect 26424 3893 26433 3927
rect 26433 3893 26467 3927
rect 26467 3893 26476 3927
rect 26424 3884 26476 3893
rect 27896 3884 27948 3936
rect 28632 3884 28684 3936
rect 31392 3927 31444 3936
rect 31392 3893 31401 3927
rect 31401 3893 31435 3927
rect 31435 3893 31444 3927
rect 31392 3884 31444 3893
rect 35164 3927 35216 3936
rect 35164 3893 35173 3927
rect 35173 3893 35207 3927
rect 35207 3893 35216 3927
rect 35164 3884 35216 3893
rect 35992 3927 36044 3936
rect 35992 3893 36001 3927
rect 36001 3893 36035 3927
rect 36035 3893 36044 3927
rect 35992 3884 36044 3893
rect 36360 3884 36412 3936
rect 37740 3927 37792 3936
rect 37740 3893 37749 3927
rect 37749 3893 37783 3927
rect 37783 3893 37792 3927
rect 37740 3884 37792 3893
rect 39764 3884 39816 3936
rect 45192 4020 45244 4072
rect 49332 4131 49384 4140
rect 49332 4097 49341 4131
rect 49341 4097 49375 4131
rect 49375 4097 49384 4131
rect 49332 4088 49384 4097
rect 49700 4088 49752 4140
rect 49792 4131 49844 4140
rect 49792 4097 49801 4131
rect 49801 4097 49835 4131
rect 49835 4097 49844 4131
rect 49792 4088 49844 4097
rect 51356 4088 51408 4140
rect 52184 4088 52236 4140
rect 55312 4088 55364 4140
rect 56692 4131 56744 4140
rect 56692 4097 56701 4131
rect 56701 4097 56735 4131
rect 56735 4097 56744 4131
rect 56692 4088 56744 4097
rect 57244 4088 57296 4140
rect 47032 4020 47084 4072
rect 49608 4020 49660 4072
rect 53656 4020 53708 4072
rect 53748 4020 53800 4072
rect 44180 3952 44232 4004
rect 49884 3995 49936 4004
rect 49884 3961 49893 3995
rect 49893 3961 49927 3995
rect 49927 3961 49936 3995
rect 49884 3952 49936 3961
rect 49976 3952 50028 4004
rect 55220 3952 55272 4004
rect 43076 3927 43128 3936
rect 43076 3893 43085 3927
rect 43085 3893 43119 3927
rect 43119 3893 43128 3927
rect 43076 3884 43128 3893
rect 43628 3884 43680 3936
rect 45928 3927 45980 3936
rect 45928 3893 45937 3927
rect 45937 3893 45971 3927
rect 45971 3893 45980 3927
rect 45928 3884 45980 3893
rect 46664 3927 46716 3936
rect 46664 3893 46673 3927
rect 46673 3893 46707 3927
rect 46707 3893 46716 3927
rect 46664 3884 46716 3893
rect 47584 3927 47636 3936
rect 47584 3893 47593 3927
rect 47593 3893 47627 3927
rect 47627 3893 47636 3927
rect 47584 3884 47636 3893
rect 47768 3884 47820 3936
rect 54484 3927 54536 3936
rect 54484 3893 54493 3927
rect 54493 3893 54527 3927
rect 54527 3893 54536 3927
rect 54484 3884 54536 3893
rect 55312 3884 55364 3936
rect 55680 3884 55732 3936
rect 56324 3884 56376 3936
rect 8174 3782 8226 3834
rect 8238 3782 8290 3834
rect 8302 3782 8354 3834
rect 8366 3782 8418 3834
rect 8430 3782 8482 3834
rect 22622 3782 22674 3834
rect 22686 3782 22738 3834
rect 22750 3782 22802 3834
rect 22814 3782 22866 3834
rect 22878 3782 22930 3834
rect 37070 3782 37122 3834
rect 37134 3782 37186 3834
rect 37198 3782 37250 3834
rect 37262 3782 37314 3834
rect 37326 3782 37378 3834
rect 51518 3782 51570 3834
rect 51582 3782 51634 3834
rect 51646 3782 51698 3834
rect 51710 3782 51762 3834
rect 51774 3782 51826 3834
rect 3792 3723 3844 3732
rect 3792 3689 3801 3723
rect 3801 3689 3835 3723
rect 3835 3689 3844 3723
rect 3792 3680 3844 3689
rect 6368 3723 6420 3732
rect 6368 3689 6377 3723
rect 6377 3689 6411 3723
rect 6411 3689 6420 3723
rect 6368 3680 6420 3689
rect 8852 3680 8904 3732
rect 9772 3680 9824 3732
rect 10784 3680 10836 3732
rect 2412 3544 2464 3596
rect 7656 3612 7708 3664
rect 13084 3612 13136 3664
rect 2964 3476 3016 3528
rect 4160 3544 4212 3596
rect 4436 3587 4488 3596
rect 4436 3553 4445 3587
rect 4445 3553 4479 3587
rect 4479 3553 4488 3587
rect 4436 3544 4488 3553
rect 5448 3544 5500 3596
rect 7196 3544 7248 3596
rect 8576 3544 8628 3596
rect 8852 3544 8904 3596
rect 12164 3544 12216 3596
rect 12348 3587 12400 3596
rect 12348 3553 12357 3587
rect 12357 3553 12391 3587
rect 12391 3553 12400 3587
rect 12348 3544 12400 3553
rect 3148 3383 3200 3392
rect 3148 3349 3157 3383
rect 3157 3349 3191 3383
rect 3191 3349 3200 3383
rect 5540 3408 5592 3460
rect 6644 3476 6696 3528
rect 7104 3476 7156 3528
rect 7748 3519 7800 3528
rect 7748 3485 7757 3519
rect 7757 3485 7791 3519
rect 7791 3485 7800 3519
rect 7748 3476 7800 3485
rect 10232 3476 10284 3528
rect 10508 3476 10560 3528
rect 9680 3451 9732 3460
rect 9680 3417 9689 3451
rect 9689 3417 9723 3451
rect 9723 3417 9732 3451
rect 9680 3408 9732 3417
rect 10416 3451 10468 3460
rect 10416 3417 10425 3451
rect 10425 3417 10459 3451
rect 10459 3417 10468 3451
rect 10416 3408 10468 3417
rect 12992 3476 13044 3528
rect 14372 3680 14424 3732
rect 15384 3680 15436 3732
rect 13728 3612 13780 3664
rect 17592 3680 17644 3732
rect 17868 3680 17920 3732
rect 18236 3723 18288 3732
rect 18236 3689 18245 3723
rect 18245 3689 18279 3723
rect 18279 3689 18288 3723
rect 18236 3680 18288 3689
rect 19156 3680 19208 3732
rect 13912 3544 13964 3596
rect 15660 3544 15712 3596
rect 16120 3544 16172 3596
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 14556 3476 14608 3528
rect 13176 3451 13228 3460
rect 13176 3417 13185 3451
rect 13185 3417 13219 3451
rect 13219 3417 13228 3451
rect 13176 3408 13228 3417
rect 3148 3340 3200 3349
rect 4528 3340 4580 3392
rect 5448 3383 5500 3392
rect 5448 3349 5457 3383
rect 5457 3349 5491 3383
rect 5491 3349 5500 3383
rect 5448 3340 5500 3349
rect 6552 3383 6604 3392
rect 6552 3349 6561 3383
rect 6561 3349 6595 3383
rect 6595 3349 6604 3383
rect 6552 3340 6604 3349
rect 8300 3340 8352 3392
rect 10692 3383 10744 3392
rect 10692 3349 10701 3383
rect 10701 3349 10735 3383
rect 10735 3349 10744 3383
rect 10692 3340 10744 3349
rect 11612 3340 11664 3392
rect 12164 3383 12216 3392
rect 12164 3349 12173 3383
rect 12173 3349 12207 3383
rect 12207 3349 12216 3383
rect 12164 3340 12216 3349
rect 12256 3383 12308 3392
rect 12256 3349 12265 3383
rect 12265 3349 12299 3383
rect 12299 3349 12308 3383
rect 12256 3340 12308 3349
rect 12624 3340 12676 3392
rect 13544 3408 13596 3460
rect 15108 3476 15160 3528
rect 15568 3408 15620 3460
rect 19616 3612 19668 3664
rect 18052 3544 18104 3596
rect 18328 3587 18380 3596
rect 18328 3553 18337 3587
rect 18337 3553 18371 3587
rect 18371 3553 18380 3587
rect 18328 3544 18380 3553
rect 19708 3587 19760 3596
rect 18512 3519 18564 3528
rect 18512 3485 18521 3519
rect 18521 3485 18555 3519
rect 18555 3485 18564 3519
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 22008 3680 22060 3732
rect 25320 3723 25372 3732
rect 25320 3689 25329 3723
rect 25329 3689 25363 3723
rect 25363 3689 25372 3723
rect 25320 3680 25372 3689
rect 30932 3723 30984 3732
rect 24584 3612 24636 3664
rect 26424 3612 26476 3664
rect 21180 3587 21232 3596
rect 21180 3553 21189 3587
rect 21189 3553 21223 3587
rect 21223 3553 21232 3587
rect 21180 3544 21232 3553
rect 26148 3544 26200 3596
rect 26976 3544 27028 3596
rect 18512 3476 18564 3485
rect 21640 3519 21692 3528
rect 21640 3485 21649 3519
rect 21649 3485 21683 3519
rect 21683 3485 21692 3519
rect 21640 3476 21692 3485
rect 23112 3519 23164 3528
rect 23112 3485 23121 3519
rect 23121 3485 23155 3519
rect 23155 3485 23164 3519
rect 23112 3476 23164 3485
rect 23388 3476 23440 3528
rect 24676 3476 24728 3528
rect 26056 3519 26108 3528
rect 26056 3485 26065 3519
rect 26065 3485 26099 3519
rect 26099 3485 26108 3519
rect 26056 3476 26108 3485
rect 26700 3476 26752 3528
rect 29000 3476 29052 3528
rect 30932 3689 30941 3723
rect 30941 3689 30975 3723
rect 30975 3689 30984 3723
rect 30932 3680 30984 3689
rect 35440 3723 35492 3732
rect 35440 3689 35449 3723
rect 35449 3689 35483 3723
rect 35483 3689 35492 3723
rect 35440 3680 35492 3689
rect 39212 3680 39264 3732
rect 30380 3587 30432 3596
rect 30380 3553 30389 3587
rect 30389 3553 30423 3587
rect 30423 3553 30432 3587
rect 30380 3544 30432 3553
rect 35164 3612 35216 3664
rect 40132 3680 40184 3732
rect 40224 3680 40276 3732
rect 42248 3680 42300 3732
rect 45744 3723 45796 3732
rect 45744 3689 45753 3723
rect 45753 3689 45787 3723
rect 45787 3689 45796 3723
rect 45744 3680 45796 3689
rect 47032 3680 47084 3732
rect 48044 3680 48096 3732
rect 31208 3544 31260 3596
rect 35348 3544 35400 3596
rect 35992 3587 36044 3596
rect 35992 3553 36001 3587
rect 36001 3553 36035 3587
rect 36035 3553 36044 3587
rect 35992 3544 36044 3553
rect 36912 3544 36964 3596
rect 38660 3587 38712 3596
rect 38660 3553 38669 3587
rect 38669 3553 38703 3587
rect 38703 3553 38712 3587
rect 38660 3544 38712 3553
rect 31576 3476 31628 3528
rect 18144 3408 18196 3460
rect 18328 3408 18380 3460
rect 21088 3408 21140 3460
rect 24860 3451 24912 3460
rect 24860 3417 24869 3451
rect 24869 3417 24903 3451
rect 24903 3417 24912 3451
rect 24860 3408 24912 3417
rect 32588 3476 32640 3528
rect 33140 3476 33192 3528
rect 33600 3476 33652 3528
rect 33784 3408 33836 3460
rect 33968 3476 34020 3528
rect 36176 3476 36228 3528
rect 38752 3476 38804 3528
rect 41604 3544 41656 3596
rect 36452 3408 36504 3460
rect 38200 3408 38252 3460
rect 38844 3451 38896 3460
rect 38844 3417 38853 3451
rect 38853 3417 38887 3451
rect 38887 3417 38896 3451
rect 38844 3408 38896 3417
rect 17868 3340 17920 3392
rect 19800 3340 19852 3392
rect 19984 3383 20036 3392
rect 19984 3349 19993 3383
rect 19993 3349 20027 3383
rect 20027 3349 20036 3383
rect 19984 3340 20036 3349
rect 21732 3340 21784 3392
rect 23572 3340 23624 3392
rect 24308 3340 24360 3392
rect 25688 3340 25740 3392
rect 26240 3340 26292 3392
rect 29092 3340 29144 3392
rect 30472 3383 30524 3392
rect 30472 3349 30481 3383
rect 30481 3349 30515 3383
rect 30515 3349 30524 3383
rect 30472 3340 30524 3349
rect 33876 3340 33928 3392
rect 34060 3383 34112 3392
rect 34060 3349 34069 3383
rect 34069 3349 34103 3383
rect 34103 3349 34112 3383
rect 34060 3340 34112 3349
rect 36084 3340 36136 3392
rect 36268 3383 36320 3392
rect 36268 3349 36277 3383
rect 36277 3349 36311 3383
rect 36311 3349 36320 3383
rect 36268 3340 36320 3349
rect 39948 3476 40000 3528
rect 44272 3612 44324 3664
rect 50160 3655 50212 3664
rect 50160 3621 50169 3655
rect 50169 3621 50203 3655
rect 50203 3621 50212 3655
rect 50160 3612 50212 3621
rect 51172 3612 51224 3664
rect 55220 3680 55272 3732
rect 56048 3680 56100 3732
rect 44640 3544 44692 3596
rect 45192 3587 45244 3596
rect 45192 3553 45201 3587
rect 45201 3553 45235 3587
rect 45235 3553 45244 3587
rect 45192 3544 45244 3553
rect 45928 3544 45980 3596
rect 49332 3587 49384 3596
rect 49332 3553 49341 3587
rect 49341 3553 49375 3587
rect 49375 3553 49384 3587
rect 49332 3544 49384 3553
rect 52184 3544 52236 3596
rect 52552 3587 52604 3596
rect 52552 3553 52561 3587
rect 52561 3553 52595 3587
rect 52595 3553 52604 3587
rect 52552 3544 52604 3553
rect 52644 3544 52696 3596
rect 42432 3476 42484 3528
rect 42616 3476 42668 3528
rect 42892 3476 42944 3528
rect 45376 3476 45428 3528
rect 46572 3519 46624 3528
rect 46572 3485 46581 3519
rect 46581 3485 46615 3519
rect 46615 3485 46624 3519
rect 46572 3476 46624 3485
rect 46664 3476 46716 3528
rect 49424 3476 49476 3528
rect 50712 3476 50764 3528
rect 50896 3519 50948 3528
rect 50896 3485 50905 3519
rect 50905 3485 50939 3519
rect 50939 3485 50948 3519
rect 50896 3476 50948 3485
rect 51172 3519 51224 3528
rect 51172 3485 51181 3519
rect 51181 3485 51215 3519
rect 51215 3485 51224 3519
rect 51172 3476 51224 3485
rect 39488 3340 39540 3392
rect 40224 3340 40276 3392
rect 47032 3408 47084 3460
rect 49332 3408 49384 3460
rect 52828 3408 52880 3460
rect 41788 3383 41840 3392
rect 41788 3349 41797 3383
rect 41797 3349 41831 3383
rect 41831 3349 41840 3383
rect 41788 3340 41840 3349
rect 45468 3340 45520 3392
rect 46940 3383 46992 3392
rect 46940 3349 46949 3383
rect 46949 3349 46983 3383
rect 46983 3349 46992 3383
rect 46940 3340 46992 3349
rect 47124 3383 47176 3392
rect 47124 3349 47133 3383
rect 47133 3349 47167 3383
rect 47167 3349 47176 3383
rect 47124 3340 47176 3349
rect 47584 3383 47636 3392
rect 47584 3349 47593 3383
rect 47593 3349 47627 3383
rect 47627 3349 47636 3383
rect 47584 3340 47636 3349
rect 48872 3340 48924 3392
rect 55496 3612 55548 3664
rect 55404 3544 55456 3596
rect 55864 3587 55916 3596
rect 55864 3553 55873 3587
rect 55873 3553 55907 3587
rect 55907 3553 55916 3587
rect 55864 3544 55916 3553
rect 56232 3544 56284 3596
rect 57428 3476 57480 3528
rect 54024 3383 54076 3392
rect 54024 3349 54033 3383
rect 54033 3349 54067 3383
rect 54067 3349 54076 3383
rect 54024 3340 54076 3349
rect 55312 3340 55364 3392
rect 55680 3383 55732 3392
rect 55680 3349 55689 3383
rect 55689 3349 55723 3383
rect 55723 3349 55732 3383
rect 55680 3340 55732 3349
rect 55772 3383 55824 3392
rect 55772 3349 55781 3383
rect 55781 3349 55815 3383
rect 55815 3349 55824 3383
rect 55772 3340 55824 3349
rect 55956 3340 56008 3392
rect 15398 3238 15450 3290
rect 15462 3238 15514 3290
rect 15526 3238 15578 3290
rect 15590 3238 15642 3290
rect 15654 3238 15706 3290
rect 29846 3238 29898 3290
rect 29910 3238 29962 3290
rect 29974 3238 30026 3290
rect 30038 3238 30090 3290
rect 30102 3238 30154 3290
rect 44294 3238 44346 3290
rect 44358 3238 44410 3290
rect 44422 3238 44474 3290
rect 44486 3238 44538 3290
rect 44550 3238 44602 3290
rect 4436 3000 4488 3052
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 5080 2932 5132 2984
rect 4988 2864 5040 2916
rect 5540 3068 5592 3120
rect 6828 3179 6880 3188
rect 6828 3145 6837 3179
rect 6837 3145 6871 3179
rect 6871 3145 6880 3179
rect 6828 3136 6880 3145
rect 7288 3136 7340 3188
rect 10140 3136 10192 3188
rect 11612 3179 11664 3188
rect 11612 3145 11621 3179
rect 11621 3145 11655 3179
rect 11655 3145 11664 3179
rect 11612 3136 11664 3145
rect 5632 3043 5684 3052
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 7380 3068 7432 3120
rect 7748 3068 7800 3120
rect 11704 3068 11756 3120
rect 5632 3000 5684 3009
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 7196 3000 7248 3052
rect 8760 3043 8812 3052
rect 7564 2932 7616 2984
rect 8760 3009 8769 3043
rect 8769 3009 8803 3043
rect 8803 3009 8812 3043
rect 8760 3000 8812 3009
rect 13360 3136 13412 3188
rect 13544 3136 13596 3188
rect 13728 3136 13780 3188
rect 15660 3136 15712 3188
rect 15844 3136 15896 3188
rect 16396 3136 16448 3188
rect 15200 3068 15252 3120
rect 18052 3136 18104 3188
rect 18512 3136 18564 3188
rect 19800 3136 19852 3188
rect 24124 3136 24176 3188
rect 24676 3136 24728 3188
rect 31208 3179 31260 3188
rect 31208 3145 31217 3179
rect 31217 3145 31251 3179
rect 31251 3145 31260 3179
rect 31208 3136 31260 3145
rect 31576 3179 31628 3188
rect 31576 3145 31585 3179
rect 31585 3145 31619 3179
rect 31619 3145 31628 3179
rect 31576 3136 31628 3145
rect 32312 3136 32364 3188
rect 34796 3136 34848 3188
rect 35256 3136 35308 3188
rect 12532 3000 12584 3052
rect 12716 3000 12768 3052
rect 12900 3043 12952 3052
rect 12900 3009 12909 3043
rect 12909 3009 12943 3043
rect 12943 3009 12952 3043
rect 13268 3043 13320 3052
rect 12900 3000 12952 3009
rect 13268 3009 13277 3043
rect 13277 3009 13311 3043
rect 13311 3009 13320 3043
rect 13268 3000 13320 3009
rect 13360 3000 13412 3052
rect 13544 3000 13596 3052
rect 14004 3000 14056 3052
rect 15752 3000 15804 3052
rect 16304 3000 16356 3052
rect 18328 3000 18380 3052
rect 19248 3000 19300 3052
rect 8300 2932 8352 2984
rect 9404 2932 9456 2984
rect 10232 2932 10284 2984
rect 12348 2932 12400 2984
rect 12992 2932 13044 2984
rect 13636 2932 13688 2984
rect 13820 2932 13872 2984
rect 14556 2932 14608 2984
rect 15292 2932 15344 2984
rect 16396 2932 16448 2984
rect 20444 3000 20496 3052
rect 28632 3111 28684 3120
rect 28632 3077 28641 3111
rect 28641 3077 28675 3111
rect 28675 3077 28684 3111
rect 28632 3068 28684 3077
rect 31392 3068 31444 3120
rect 33876 3111 33928 3120
rect 33876 3077 33885 3111
rect 33885 3077 33919 3111
rect 33919 3077 33928 3111
rect 33876 3068 33928 3077
rect 24676 3000 24728 3052
rect 24860 3000 24912 3052
rect 26608 3000 26660 3052
rect 27344 3000 27396 3052
rect 29092 3000 29144 3052
rect 5540 2864 5592 2916
rect 2780 2796 2832 2848
rect 2964 2796 3016 2848
rect 4068 2796 4120 2848
rect 4344 2839 4396 2848
rect 4344 2805 4353 2839
rect 4353 2805 4387 2839
rect 4387 2805 4396 2839
rect 4344 2796 4396 2805
rect 4436 2796 4488 2848
rect 5264 2796 5316 2848
rect 5356 2796 5408 2848
rect 8944 2864 8996 2916
rect 9220 2864 9272 2916
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 6368 2796 6420 2848
rect 7472 2796 7524 2848
rect 8576 2839 8628 2848
rect 8576 2805 8585 2839
rect 8585 2805 8619 2839
rect 8619 2805 8628 2839
rect 8576 2796 8628 2805
rect 10784 2796 10836 2848
rect 13912 2864 13964 2916
rect 24492 2932 24544 2984
rect 30380 2932 30432 2984
rect 32772 3000 32824 3052
rect 33508 3000 33560 3052
rect 35164 3000 35216 3052
rect 31760 2932 31812 2984
rect 34520 2932 34572 2984
rect 34612 2932 34664 2984
rect 36820 2932 36872 2984
rect 38936 3136 38988 3188
rect 39856 3136 39908 3188
rect 41696 3136 41748 3188
rect 40592 3068 40644 3120
rect 41604 3068 41656 3120
rect 42524 3136 42576 3188
rect 45008 3136 45060 3188
rect 43076 3068 43128 3120
rect 43168 3068 43220 3120
rect 46112 3136 46164 3188
rect 49424 3136 49476 3188
rect 49608 3136 49660 3188
rect 52644 3136 52696 3188
rect 47032 3111 47084 3120
rect 40132 3000 40184 3052
rect 38108 2932 38160 2984
rect 40592 2932 40644 2984
rect 43904 3000 43956 3052
rect 12256 2796 12308 2848
rect 12624 2796 12676 2848
rect 13360 2796 13412 2848
rect 14372 2839 14424 2848
rect 14372 2805 14381 2839
rect 14381 2805 14415 2839
rect 14415 2805 14424 2839
rect 14372 2796 14424 2805
rect 15568 2839 15620 2848
rect 15568 2805 15577 2839
rect 15577 2805 15611 2839
rect 15611 2805 15620 2839
rect 15568 2796 15620 2805
rect 19340 2864 19392 2916
rect 20996 2864 21048 2916
rect 23756 2864 23808 2916
rect 23848 2864 23900 2916
rect 26884 2864 26936 2916
rect 31484 2864 31536 2916
rect 24032 2796 24084 2848
rect 25964 2796 26016 2848
rect 26516 2796 26568 2848
rect 29552 2796 29604 2848
rect 30196 2796 30248 2848
rect 34244 2796 34296 2848
rect 36452 2907 36504 2916
rect 36452 2873 36461 2907
rect 36461 2873 36495 2907
rect 36495 2873 36504 2907
rect 36452 2864 36504 2873
rect 36544 2864 36596 2916
rect 38660 2864 38712 2916
rect 35348 2839 35400 2848
rect 35348 2805 35357 2839
rect 35357 2805 35391 2839
rect 35391 2805 35400 2839
rect 35348 2796 35400 2805
rect 36728 2796 36780 2848
rect 41236 2864 41288 2916
rect 43076 2907 43128 2916
rect 43076 2873 43085 2907
rect 43085 2873 43119 2907
rect 43119 2873 43128 2907
rect 43076 2864 43128 2873
rect 42432 2839 42484 2848
rect 42432 2805 42441 2839
rect 42441 2805 42475 2839
rect 42475 2805 42484 2839
rect 42432 2796 42484 2805
rect 42800 2796 42852 2848
rect 44272 2864 44324 2916
rect 43260 2796 43312 2848
rect 45192 3000 45244 3052
rect 47032 3077 47041 3111
rect 47041 3077 47075 3111
rect 47075 3077 47084 3111
rect 47032 3068 47084 3077
rect 46572 3000 46624 3052
rect 49884 3068 49936 3120
rect 50068 3111 50120 3120
rect 50068 3077 50077 3111
rect 50077 3077 50111 3111
rect 50111 3077 50120 3111
rect 50068 3068 50120 3077
rect 50712 3068 50764 3120
rect 47216 3000 47268 3052
rect 50804 3000 50856 3052
rect 52460 3068 52512 3120
rect 51356 3000 51408 3052
rect 55864 3068 55916 3120
rect 56048 3111 56100 3120
rect 56048 3077 56057 3111
rect 56057 3077 56091 3111
rect 56091 3077 56100 3111
rect 56048 3068 56100 3077
rect 55956 3000 56008 3052
rect 56324 3000 56376 3052
rect 45560 2932 45612 2984
rect 45284 2864 45336 2916
rect 48596 2864 48648 2916
rect 55496 2932 55548 2984
rect 56232 2975 56284 2984
rect 56232 2941 56241 2975
rect 56241 2941 56275 2975
rect 56275 2941 56284 2975
rect 56232 2932 56284 2941
rect 47676 2796 47728 2848
rect 49884 2796 49936 2848
rect 50436 2796 50488 2848
rect 50988 2864 51040 2916
rect 52368 2864 52420 2916
rect 54208 2839 54260 2848
rect 54208 2805 54217 2839
rect 54217 2805 54251 2839
rect 54251 2805 54260 2839
rect 54208 2796 54260 2805
rect 55588 2796 55640 2848
rect 55772 2796 55824 2848
rect 56600 2796 56652 2848
rect 8174 2694 8226 2746
rect 8238 2694 8290 2746
rect 8302 2694 8354 2746
rect 8366 2694 8418 2746
rect 8430 2694 8482 2746
rect 22622 2694 22674 2746
rect 22686 2694 22738 2746
rect 22750 2694 22802 2746
rect 22814 2694 22866 2746
rect 22878 2694 22930 2746
rect 37070 2694 37122 2746
rect 37134 2694 37186 2746
rect 37198 2694 37250 2746
rect 37262 2694 37314 2746
rect 37326 2694 37378 2746
rect 51518 2694 51570 2746
rect 51582 2694 51634 2746
rect 51646 2694 51698 2746
rect 51710 2694 51762 2746
rect 51774 2694 51826 2746
rect 4620 2592 4672 2644
rect 5080 2592 5132 2644
rect 5540 2592 5592 2644
rect 7288 2592 7340 2644
rect 5448 2524 5500 2576
rect 7104 2524 7156 2576
rect 2872 2456 2924 2508
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 3884 2431 3936 2440
rect 3884 2397 3893 2431
rect 3893 2397 3927 2431
rect 3927 2397 3936 2431
rect 3884 2388 3936 2397
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 5264 2456 5316 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 5632 2499 5684 2508
rect 5632 2465 5666 2499
rect 5666 2465 5684 2499
rect 5632 2456 5684 2465
rect 10416 2592 10468 2644
rect 10508 2524 10560 2576
rect 8852 2456 8904 2508
rect 11612 2592 11664 2644
rect 13268 2592 13320 2644
rect 14004 2592 14056 2644
rect 16488 2592 16540 2644
rect 20720 2592 20772 2644
rect 24584 2592 24636 2644
rect 26700 2592 26752 2644
rect 33876 2592 33928 2644
rect 34520 2592 34572 2644
rect 34796 2592 34848 2644
rect 36820 2592 36872 2644
rect 38016 2592 38068 2644
rect 38844 2592 38896 2644
rect 40316 2592 40368 2644
rect 44272 2592 44324 2644
rect 49516 2635 49568 2644
rect 49516 2601 49525 2635
rect 49525 2601 49559 2635
rect 49559 2601 49568 2635
rect 49516 2592 49568 2601
rect 49608 2592 49660 2644
rect 4988 2388 5040 2440
rect 4344 2252 4396 2304
rect 5356 2252 5408 2304
rect 5724 2320 5776 2372
rect 7380 2388 7432 2440
rect 9220 2431 9272 2440
rect 9220 2397 9229 2431
rect 9229 2397 9263 2431
rect 9263 2397 9272 2431
rect 9220 2388 9272 2397
rect 12624 2456 12676 2508
rect 14096 2524 14148 2576
rect 19064 2524 19116 2576
rect 22652 2524 22704 2576
rect 25136 2524 25188 2576
rect 26608 2524 26660 2576
rect 30380 2524 30432 2576
rect 32036 2524 32088 2576
rect 33692 2524 33744 2576
rect 37832 2524 37884 2576
rect 15568 2456 15620 2508
rect 18420 2456 18472 2508
rect 12256 2431 12308 2440
rect 7104 2320 7156 2372
rect 12256 2397 12265 2431
rect 12265 2397 12299 2431
rect 12299 2397 12308 2431
rect 12256 2388 12308 2397
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 12900 2388 12952 2440
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 7748 2252 7800 2304
rect 8760 2252 8812 2304
rect 9220 2252 9272 2304
rect 14004 2320 14056 2372
rect 11612 2252 11664 2304
rect 13176 2252 13228 2304
rect 18328 2388 18380 2440
rect 22928 2456 22980 2508
rect 22284 2388 22336 2440
rect 22468 2388 22520 2440
rect 22100 2320 22152 2372
rect 18788 2252 18840 2304
rect 23296 2388 23348 2440
rect 24216 2456 24268 2508
rect 24676 2499 24728 2508
rect 24676 2465 24685 2499
rect 24685 2465 24719 2499
rect 24719 2465 24728 2499
rect 24676 2456 24728 2465
rect 24768 2456 24820 2508
rect 26976 2499 27028 2508
rect 23664 2388 23716 2440
rect 26976 2465 26985 2499
rect 26985 2465 27019 2499
rect 27019 2465 27028 2499
rect 26976 2456 27028 2465
rect 29276 2456 29328 2508
rect 30656 2456 30708 2508
rect 24860 2320 24912 2372
rect 24492 2252 24544 2304
rect 26332 2320 26384 2372
rect 27528 2320 27580 2372
rect 30932 2388 30984 2440
rect 31208 2388 31260 2440
rect 36268 2456 36320 2508
rect 32956 2388 33008 2440
rect 37372 2456 37424 2508
rect 40868 2456 40920 2508
rect 45192 2524 45244 2576
rect 45836 2524 45888 2576
rect 50436 2524 50488 2576
rect 44548 2456 44600 2508
rect 44640 2456 44692 2508
rect 49700 2456 49752 2508
rect 57428 2592 57480 2644
rect 55864 2524 55916 2576
rect 56692 2456 56744 2508
rect 38016 2388 38068 2440
rect 25596 2295 25648 2304
rect 25596 2261 25605 2295
rect 25605 2261 25639 2295
rect 25639 2261 25648 2295
rect 25596 2252 25648 2261
rect 25780 2295 25832 2304
rect 25780 2261 25789 2295
rect 25789 2261 25823 2295
rect 25823 2261 25832 2295
rect 25780 2252 25832 2261
rect 28356 2295 28408 2304
rect 28356 2261 28365 2295
rect 28365 2261 28399 2295
rect 28399 2261 28408 2295
rect 28356 2252 28408 2261
rect 35440 2320 35492 2372
rect 33876 2252 33928 2304
rect 37004 2252 37056 2304
rect 37096 2252 37148 2304
rect 39948 2388 40000 2440
rect 39764 2320 39816 2372
rect 40132 2252 40184 2304
rect 41972 2252 42024 2304
rect 46848 2388 46900 2440
rect 51448 2431 51500 2440
rect 45284 2320 45336 2372
rect 51448 2397 51457 2431
rect 51457 2397 51491 2431
rect 51491 2397 51500 2431
rect 51448 2388 51500 2397
rect 52736 2431 52788 2440
rect 52736 2397 52745 2431
rect 52745 2397 52779 2431
rect 52779 2397 52788 2431
rect 52736 2388 52788 2397
rect 54760 2388 54812 2440
rect 56232 2431 56284 2440
rect 56232 2397 56241 2431
rect 56241 2397 56275 2431
rect 56275 2397 56284 2431
rect 56232 2388 56284 2397
rect 44824 2252 44876 2304
rect 45468 2252 45520 2304
rect 47584 2252 47636 2304
rect 50804 2252 50856 2304
rect 51172 2252 51224 2304
rect 15398 2150 15450 2202
rect 15462 2150 15514 2202
rect 15526 2150 15578 2202
rect 15590 2150 15642 2202
rect 15654 2150 15706 2202
rect 29846 2150 29898 2202
rect 29910 2150 29962 2202
rect 29974 2150 30026 2202
rect 30038 2150 30090 2202
rect 30102 2150 30154 2202
rect 44294 2150 44346 2202
rect 44358 2150 44410 2202
rect 44422 2150 44474 2202
rect 44486 2150 44538 2202
rect 44550 2150 44602 2202
rect 3884 2048 3936 2100
rect 8944 2048 8996 2100
rect 10508 2048 10560 2100
rect 4712 1980 4764 2032
rect 11152 1980 11204 2032
rect 12256 2048 12308 2100
rect 18236 2048 18288 2100
rect 18420 2048 18472 2100
rect 21548 2048 21600 2100
rect 37004 2048 37056 2100
rect 40132 2048 40184 2100
rect 41420 2048 41472 2100
rect 45192 2048 45244 2100
rect 46388 2048 46440 2100
rect 51448 2048 51500 2100
rect 13820 1980 13872 2032
rect 18328 1980 18380 2032
rect 20168 1980 20220 2032
rect 23296 1980 23348 2032
rect 45376 1980 45428 2032
rect 46940 1980 46992 2032
rect 52736 1980 52788 2032
rect 4528 1912 4580 1964
rect 25596 1912 25648 1964
rect 30472 1912 30524 1964
rect 41604 1912 41656 1964
rect 7748 1844 7800 1896
rect 12440 1844 12492 1896
rect 12624 1844 12676 1896
rect 18604 1844 18656 1896
rect 23112 1844 23164 1896
rect 41788 1844 41840 1896
rect 49424 1912 49476 1964
rect 56232 1912 56284 1964
rect 54208 1844 54260 1896
rect 3056 1776 3108 1828
rect 8208 1776 8260 1828
rect 10692 1776 10744 1828
rect 24768 1776 24820 1828
rect 6552 1708 6604 1760
rect 18144 1708 18196 1760
rect 22468 1708 22520 1760
rect 40040 1708 40092 1760
rect 43076 1708 43128 1760
rect 44732 1708 44784 1760
rect 46848 1708 46900 1760
rect 47124 1776 47176 1828
rect 55772 1776 55824 1828
rect 54024 1708 54076 1760
rect 12440 1640 12492 1692
rect 21640 1640 21692 1692
rect 23664 1640 23716 1692
rect 44824 1640 44876 1692
rect 7196 1436 7248 1488
rect 7932 1436 7984 1488
rect 7012 1368 7064 1420
rect 7748 1368 7800 1420
rect 9220 1368 9272 1420
rect 25412 1368 25464 1420
rect 27528 1368 27580 1420
rect 35900 1368 35952 1420
rect 37096 1368 37148 1420
rect 38384 1368 38436 1420
rect 39948 1368 40000 1420
rect 48320 1368 48372 1420
rect 49608 1368 49660 1420
rect 8024 1300 8076 1352
<< metal2 >>
rect 3974 9200 4030 10000
rect 4434 9200 4490 10000
rect 4894 9330 4950 10000
rect 4894 9302 5028 9330
rect 4894 9200 4950 9302
rect 4448 7410 4476 9200
rect 5000 7410 5028 9302
rect 5354 9200 5410 10000
rect 5814 9200 5870 10000
rect 6274 9330 6330 10000
rect 6274 9302 6408 9330
rect 6274 9200 6330 9302
rect 5828 7410 5856 9200
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 5816 7404 5868 7410
rect 5816 7346 5868 7352
rect 6380 6866 6408 9302
rect 6734 9200 6790 10000
rect 7194 9330 7250 10000
rect 7654 9330 7710 10000
rect 7116 9302 7250 9330
rect 7116 7410 7144 9302
rect 7194 9200 7250 9302
rect 7576 9302 7710 9330
rect 7576 7410 7604 9302
rect 7654 9200 7710 9302
rect 8114 9200 8170 10000
rect 8574 9330 8630 10000
rect 8404 9302 8630 9330
rect 8404 7410 8432 9302
rect 8574 9200 8630 9302
rect 9034 9330 9090 10000
rect 9034 9302 9168 9330
rect 9034 9200 9090 9302
rect 9140 7410 9168 9302
rect 9494 9200 9550 10000
rect 9954 9200 10010 10000
rect 10414 9200 10470 10000
rect 10874 9200 10930 10000
rect 11334 9330 11390 10000
rect 11794 9330 11850 10000
rect 11334 9302 11468 9330
rect 11334 9200 11390 9302
rect 9968 7410 9996 9200
rect 10428 7410 10456 9200
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 8174 7100 8482 7109
rect 8174 7098 8180 7100
rect 8236 7098 8260 7100
rect 8316 7098 8340 7100
rect 8396 7098 8420 7100
rect 8476 7098 8482 7100
rect 8236 7046 8238 7098
rect 8418 7046 8420 7098
rect 8174 7044 8180 7046
rect 8236 7044 8260 7046
rect 8316 7044 8340 7046
rect 8396 7044 8420 7046
rect 8476 7044 8482 7046
rect 8174 7035 8482 7044
rect 11440 6866 11468 9302
rect 11794 9302 11928 9330
rect 11794 9200 11850 9302
rect 11900 7410 11928 9302
rect 12254 9200 12310 10000
rect 12714 9330 12770 10000
rect 12636 9302 12770 9330
rect 12636 7410 12664 9302
rect 12714 9200 12770 9302
rect 13174 9330 13230 10000
rect 13174 9302 13308 9330
rect 13174 9200 13230 9302
rect 13280 7410 13308 9302
rect 13634 9200 13690 10000
rect 14094 9200 14150 10000
rect 14554 9330 14610 10000
rect 14554 9302 14688 9330
rect 14554 9200 14610 9302
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 14108 6866 14136 9200
rect 14660 7410 14688 9302
rect 15014 9200 15070 10000
rect 15474 9330 15530 10000
rect 15304 9302 15530 9330
rect 15304 7410 15332 9302
rect 15474 9200 15530 9302
rect 15934 9200 15990 10000
rect 16394 9200 16450 10000
rect 16854 9330 16910 10000
rect 17314 9330 17370 10000
rect 16854 9302 16988 9330
rect 16854 9200 16910 9302
rect 15398 7644 15706 7653
rect 15398 7642 15404 7644
rect 15460 7642 15484 7644
rect 15540 7642 15564 7644
rect 15620 7642 15644 7644
rect 15700 7642 15706 7644
rect 15460 7590 15462 7642
rect 15642 7590 15644 7642
rect 15398 7588 15404 7590
rect 15460 7588 15484 7590
rect 15540 7588 15564 7590
rect 15620 7588 15644 7590
rect 15700 7588 15706 7590
rect 15398 7579 15706 7588
rect 15948 7410 15976 9200
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15936 7404 15988 7410
rect 15936 7346 15988 7352
rect 16960 6866 16988 9302
rect 17236 9302 17370 9330
rect 17236 7410 17264 9302
rect 17314 9200 17370 9302
rect 17774 9200 17830 10000
rect 18234 9330 18290 10000
rect 18064 9302 18290 9330
rect 18064 7410 18092 9302
rect 18234 9200 18290 9302
rect 18694 9200 18750 10000
rect 19154 9200 19210 10000
rect 19614 9330 19670 10000
rect 19536 9302 19670 9330
rect 18708 7410 18736 9200
rect 19536 7410 19564 9302
rect 19614 9200 19670 9302
rect 20074 9330 20130 10000
rect 20074 9302 20208 9330
rect 20074 9200 20130 9302
rect 20180 7410 20208 9302
rect 20534 9200 20590 10000
rect 20994 9200 21050 10000
rect 21454 9330 21510 10000
rect 21284 9302 21510 9330
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 18052 7404 18104 7410
rect 18052 7346 18104 7352
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 21008 6866 21036 9200
rect 21284 7410 21312 9302
rect 21454 9200 21510 9302
rect 21914 9200 21970 10000
rect 22374 9200 22430 10000
rect 22834 9330 22890 10000
rect 22834 9302 22968 9330
rect 22834 9200 22890 9302
rect 22388 7410 22416 9200
rect 22940 7410 22968 9302
rect 23294 9200 23350 10000
rect 23754 9330 23810 10000
rect 23676 9302 23810 9330
rect 23676 7410 23704 9302
rect 23754 9200 23810 9302
rect 24214 9330 24270 10000
rect 24214 9302 24440 9330
rect 24214 9200 24270 9302
rect 21272 7404 21324 7410
rect 21272 7346 21324 7352
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22928 7404 22980 7410
rect 22928 7346 22980 7352
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 22622 7100 22930 7109
rect 22622 7098 22628 7100
rect 22684 7098 22708 7100
rect 22764 7098 22788 7100
rect 22844 7098 22868 7100
rect 22924 7098 22930 7100
rect 22684 7046 22686 7098
rect 22866 7046 22868 7098
rect 22622 7044 22628 7046
rect 22684 7044 22708 7046
rect 22764 7044 22788 7046
rect 22844 7044 22868 7046
rect 22924 7044 22930 7046
rect 22622 7035 22930 7044
rect 24412 6866 24440 9302
rect 24674 9200 24730 10000
rect 25134 9200 25190 10000
rect 25594 9200 25650 10000
rect 26054 9200 26110 10000
rect 26514 9330 26570 10000
rect 26436 9302 26570 9330
rect 25148 7410 25176 9200
rect 25608 7410 25636 9200
rect 26436 7410 26464 9302
rect 26514 9200 26570 9302
rect 26974 9200 27030 10000
rect 27434 9200 27490 10000
rect 27894 9330 27950 10000
rect 27724 9302 27950 9330
rect 25136 7404 25188 7410
rect 25136 7346 25188 7352
rect 25596 7404 25648 7410
rect 25596 7346 25648 7352
rect 26424 7404 26476 7410
rect 26424 7346 26476 7352
rect 26988 6866 27016 9200
rect 27724 7410 27752 9302
rect 27894 9200 27950 9302
rect 28354 9200 28410 10000
rect 28814 9200 28870 10000
rect 29274 9330 29330 10000
rect 29012 9302 29330 9330
rect 28368 7410 28396 9200
rect 29012 7410 29040 9302
rect 29274 9200 29330 9302
rect 29734 9200 29790 10000
rect 30194 9200 30250 10000
rect 30654 9330 30710 10000
rect 30576 9302 30710 9330
rect 29748 7410 29776 9200
rect 29846 7644 30154 7653
rect 29846 7642 29852 7644
rect 29908 7642 29932 7644
rect 29988 7642 30012 7644
rect 30068 7642 30092 7644
rect 30148 7642 30154 7644
rect 29908 7590 29910 7642
rect 30090 7590 30092 7642
rect 29846 7588 29852 7590
rect 29908 7588 29932 7590
rect 29988 7588 30012 7590
rect 30068 7588 30092 7590
rect 30148 7588 30154 7590
rect 29846 7579 30154 7588
rect 30576 7410 30604 9302
rect 30654 9200 30710 9302
rect 31114 9330 31170 10000
rect 31114 9302 31248 9330
rect 31114 9200 31170 9302
rect 31220 7410 31248 9302
rect 31574 9200 31630 10000
rect 32034 9330 32090 10000
rect 32494 9330 32550 10000
rect 32034 9302 32168 9330
rect 32034 9200 32090 9302
rect 32140 7410 32168 9302
rect 32494 9302 32812 9330
rect 32494 9200 32550 9302
rect 32784 7410 32812 9302
rect 32954 9200 33010 10000
rect 33414 9200 33470 10000
rect 33874 9200 33930 10000
rect 34334 9200 34390 10000
rect 34794 9200 34850 10000
rect 35254 9200 35310 10000
rect 35714 9200 35770 10000
rect 36174 9330 36230 10000
rect 36174 9302 36308 9330
rect 36174 9200 36230 9302
rect 33428 7410 33456 9200
rect 33888 7410 33916 9200
rect 34808 7410 34836 9200
rect 27712 7404 27764 7410
rect 27712 7346 27764 7352
rect 28356 7404 28408 7410
rect 28356 7346 28408 7352
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 29736 7404 29788 7410
rect 29736 7346 29788 7352
rect 30564 7404 30616 7410
rect 30564 7346 30616 7352
rect 31208 7404 31260 7410
rect 31208 7346 31260 7352
rect 32128 7404 32180 7410
rect 32128 7346 32180 7352
rect 32772 7404 32824 7410
rect 32772 7346 32824 7352
rect 33416 7404 33468 7410
rect 33416 7346 33468 7352
rect 33876 7404 33928 7410
rect 33876 7346 33928 7352
rect 34796 7404 34848 7410
rect 34796 7346 34848 7352
rect 35268 7342 35296 9200
rect 35256 7336 35308 7342
rect 35256 7278 35308 7284
rect 36280 6866 36308 9302
rect 36634 9200 36690 10000
rect 37094 9200 37150 10000
rect 37554 9200 37610 10000
rect 38014 9200 38070 10000
rect 38474 9200 38530 10000
rect 38934 9200 38990 10000
rect 39394 9200 39450 10000
rect 39854 9200 39910 10000
rect 40314 9330 40370 10000
rect 40774 9330 40830 10000
rect 40314 9302 40540 9330
rect 40314 9200 40370 9302
rect 36648 7410 36676 9200
rect 37568 7410 37596 9200
rect 38028 7410 38056 9200
rect 38948 7410 38976 9200
rect 36636 7404 36688 7410
rect 36636 7346 36688 7352
rect 37556 7404 37608 7410
rect 37556 7346 37608 7352
rect 38016 7404 38068 7410
rect 38016 7346 38068 7352
rect 38936 7404 38988 7410
rect 38936 7346 38988 7352
rect 37070 7100 37378 7109
rect 37070 7098 37076 7100
rect 37132 7098 37156 7100
rect 37212 7098 37236 7100
rect 37292 7098 37316 7100
rect 37372 7098 37378 7100
rect 37132 7046 37134 7098
rect 37314 7046 37316 7098
rect 37070 7044 37076 7046
rect 37132 7044 37156 7046
rect 37212 7044 37236 7046
rect 37292 7044 37316 7046
rect 37372 7044 37378 7046
rect 37070 7035 37378 7044
rect 39408 6866 39436 9200
rect 40512 7410 40540 9302
rect 40774 9302 41184 9330
rect 40774 9200 40830 9302
rect 41156 7410 41184 9302
rect 41234 9200 41290 10000
rect 41694 9200 41750 10000
rect 42154 9330 42210 10000
rect 42154 9302 42472 9330
rect 42154 9200 42210 9302
rect 41708 7410 41736 9200
rect 40500 7404 40552 7410
rect 40500 7346 40552 7352
rect 41144 7404 41196 7410
rect 41144 7346 41196 7352
rect 41696 7404 41748 7410
rect 41696 7346 41748 7352
rect 42444 7274 42472 9302
rect 42614 9200 42670 10000
rect 43074 9200 43130 10000
rect 43534 9330 43590 10000
rect 43534 9302 43668 9330
rect 43534 9200 43590 9302
rect 43088 7410 43116 9200
rect 43076 7404 43128 7410
rect 43076 7346 43128 7352
rect 42432 7268 42484 7274
rect 42432 7210 42484 7216
rect 43640 6866 43668 9302
rect 43994 9200 44050 10000
rect 44454 9200 44510 10000
rect 44914 9330 44970 10000
rect 44914 9302 45232 9330
rect 44914 9200 44970 9302
rect 44468 7970 44496 9200
rect 44468 7942 44680 7970
rect 44294 7644 44602 7653
rect 44294 7642 44300 7644
rect 44356 7642 44380 7644
rect 44436 7642 44460 7644
rect 44516 7642 44540 7644
rect 44596 7642 44602 7644
rect 44356 7590 44358 7642
rect 44538 7590 44540 7642
rect 44294 7588 44300 7590
rect 44356 7588 44380 7590
rect 44436 7588 44460 7590
rect 44516 7588 44540 7590
rect 44596 7588 44602 7590
rect 44294 7579 44602 7588
rect 44652 7410 44680 7942
rect 45204 7410 45232 9302
rect 45374 9200 45430 10000
rect 45834 9200 45890 10000
rect 46294 9200 46350 10000
rect 46754 9200 46810 10000
rect 47214 9330 47270 10000
rect 47214 9302 47624 9330
rect 47214 9200 47270 9302
rect 45848 7410 45876 9200
rect 44640 7404 44692 7410
rect 44640 7346 44692 7352
rect 45192 7404 45244 7410
rect 45192 7346 45244 7352
rect 45836 7404 45888 7410
rect 45836 7346 45888 7352
rect 46308 6866 46336 9200
rect 47596 7410 47624 9302
rect 47674 9200 47730 10000
rect 48134 9200 48190 10000
rect 48594 9330 48650 10000
rect 48594 9302 48912 9330
rect 48594 9200 48650 9302
rect 47688 7410 47716 9200
rect 48884 7410 48912 9302
rect 49054 9200 49110 10000
rect 49514 9200 49570 10000
rect 49974 9330 50030 10000
rect 49974 9302 50200 9330
rect 49974 9200 50030 9302
rect 47584 7404 47636 7410
rect 47584 7346 47636 7352
rect 47676 7404 47728 7410
rect 47676 7346 47728 7352
rect 48872 7404 48924 7410
rect 48872 7346 48924 7352
rect 49068 6866 49096 9200
rect 50172 7410 50200 9302
rect 50434 9200 50490 10000
rect 50894 9200 50950 10000
rect 51354 9330 51410 10000
rect 51814 9330 51870 10000
rect 51354 9302 51488 9330
rect 51354 9200 51410 9302
rect 50448 7410 50476 9200
rect 51460 7410 51488 9302
rect 51814 9302 52224 9330
rect 51814 9200 51870 9302
rect 52196 7410 52224 9302
rect 52274 9200 52330 10000
rect 52734 9330 52790 10000
rect 53194 9330 53250 10000
rect 52734 9302 53144 9330
rect 52734 9200 52790 9302
rect 53116 7410 53144 9302
rect 53194 9302 53512 9330
rect 53194 9200 53250 9302
rect 53484 7410 53512 9302
rect 53654 9200 53710 10000
rect 54114 9330 54170 10000
rect 54574 9330 54630 10000
rect 54114 9302 54248 9330
rect 54114 9200 54170 9302
rect 50160 7404 50212 7410
rect 50160 7346 50212 7352
rect 50436 7404 50488 7410
rect 50436 7346 50488 7352
rect 51448 7404 51500 7410
rect 51448 7346 51500 7352
rect 52184 7404 52236 7410
rect 52184 7346 52236 7352
rect 53104 7404 53156 7410
rect 53104 7346 53156 7352
rect 53472 7404 53524 7410
rect 53472 7346 53524 7352
rect 51518 7100 51826 7109
rect 51518 7098 51524 7100
rect 51580 7098 51604 7100
rect 51660 7098 51684 7100
rect 51740 7098 51764 7100
rect 51820 7098 51826 7100
rect 51580 7046 51582 7098
rect 51762 7046 51764 7098
rect 51518 7044 51524 7046
rect 51580 7044 51604 7046
rect 51660 7044 51684 7046
rect 51740 7044 51764 7046
rect 51820 7044 51826 7046
rect 51518 7035 51826 7044
rect 54220 6866 54248 9302
rect 54574 9302 54984 9330
rect 54574 9200 54630 9302
rect 54956 7426 54984 9302
rect 55034 9200 55090 10000
rect 55494 9200 55550 10000
rect 55954 9330 56010 10000
rect 55954 9302 56272 9330
rect 55954 9200 56010 9302
rect 54956 7410 55260 7426
rect 55508 7410 55536 9200
rect 56244 7410 56272 9302
rect 54956 7404 55272 7410
rect 54956 7398 55220 7404
rect 55220 7346 55272 7352
rect 55496 7404 55548 7410
rect 55496 7346 55548 7352
rect 56232 7404 56284 7410
rect 56232 7346 56284 7352
rect 6368 6860 6420 6866
rect 6368 6802 6420 6808
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 26976 6860 27028 6866
rect 26976 6802 27028 6808
rect 36268 6860 36320 6866
rect 36268 6802 36320 6808
rect 39396 6860 39448 6866
rect 39396 6802 39448 6808
rect 43628 6860 43680 6866
rect 43628 6802 43680 6808
rect 46296 6860 46348 6866
rect 46296 6802 46348 6808
rect 49056 6860 49108 6866
rect 49056 6802 49108 6808
rect 54208 6860 54260 6866
rect 54208 6802 54260 6808
rect 27344 6724 27396 6730
rect 27344 6666 27396 6672
rect 47032 6724 47084 6730
rect 47032 6666 47084 6672
rect 48136 6724 48188 6730
rect 48136 6666 48188 6672
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 8668 6248 8720 6254
rect 8668 6190 8720 6196
rect 8174 6012 8482 6021
rect 8174 6010 8180 6012
rect 8236 6010 8260 6012
rect 8316 6010 8340 6012
rect 8396 6010 8420 6012
rect 8476 6010 8482 6012
rect 8236 5958 8238 6010
rect 8418 5958 8420 6010
rect 8174 5956 8180 5958
rect 8236 5956 8260 5958
rect 8316 5956 8340 5958
rect 8396 5956 8420 5958
rect 8476 5956 8482 5958
rect 8174 5947 8482 5956
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 4344 5840 4396 5846
rect 4344 5782 4396 5788
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3424 5024 3476 5030
rect 3424 4966 3476 4972
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3252 4214 3280 4558
rect 3148 4208 3200 4214
rect 3148 4150 3200 4156
rect 3240 4208 3292 4214
rect 3240 4150 3292 4156
rect 3056 3936 3108 3942
rect 3056 3878 3108 3884
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2424 2446 2452 3538
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2976 2854 3004 3470
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2792 2496 2820 2790
rect 2872 2508 2924 2514
rect 2792 2468 2872 2496
rect 2872 2450 2924 2456
rect 3068 2446 3096 3878
rect 3160 3398 3188 4150
rect 3436 4146 3464 4966
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3804 4282 3832 4558
rect 4080 4554 4108 5102
rect 4172 4622 4200 5578
rect 4356 5370 4384 5782
rect 5460 5522 5488 5850
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7748 5568 7800 5574
rect 5460 5494 5580 5522
rect 7748 5510 7800 5516
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 4264 5222 4476 5250
rect 4264 4826 4292 5222
rect 4448 5166 4476 5222
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4632 4826 4660 5170
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4724 4622 4752 4966
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3804 3738 3832 4082
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3148 3392 3200 3398
rect 3146 3360 3148 3369
rect 3200 3360 3202 3369
rect 3146 3295 3202 3304
rect 4080 2854 4108 4490
rect 4172 4146 4200 4558
rect 5184 4486 5212 5170
rect 5368 5137 5396 5170
rect 5354 5128 5410 5137
rect 5354 5063 5410 5072
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4264 4146 4292 4422
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4172 3602 4200 3878
rect 4434 3632 4490 3641
rect 4160 3596 4212 3602
rect 5460 3602 5488 5306
rect 5552 5234 5580 5494
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5448 3596 5500 3602
rect 4434 3567 4436 3576
rect 4160 3538 4212 3544
rect 4488 3567 4490 3576
rect 4436 3538 4488 3544
rect 5276 3556 5448 3584
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4448 2854 4476 2994
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 4344 2848 4396 2854
rect 4344 2790 4396 2796
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 4080 2553 4108 2790
rect 4066 2544 4122 2553
rect 4066 2479 4122 2488
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3068 1834 3096 2382
rect 3896 2106 3924 2382
rect 4356 2310 4384 2790
rect 4344 2304 4396 2310
rect 4344 2246 4396 2252
rect 3884 2100 3936 2106
rect 3884 2042 3936 2048
rect 4540 1970 4568 3334
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4632 2650 4660 2994
rect 5080 2984 5132 2990
rect 5080 2926 5132 2932
rect 4988 2916 5040 2922
rect 4988 2858 5040 2864
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 5000 2446 5028 2858
rect 5092 2650 5120 2926
rect 5276 2854 5304 3556
rect 5500 3556 5672 3584
rect 5448 3538 5500 3544
rect 5446 3496 5502 3505
rect 5446 3431 5502 3440
rect 5540 3460 5592 3466
rect 5460 3398 5488 3431
rect 5540 3402 5592 3408
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5552 3126 5580 3402
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5552 2922 5580 3062
rect 5644 3058 5672 3556
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5276 2514 5304 2790
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 4724 2038 4752 2382
rect 5368 2310 5396 2790
rect 5552 2774 5580 2858
rect 5828 2854 5856 4558
rect 6288 4554 6316 5238
rect 6564 4622 6592 5238
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6276 4548 6328 4554
rect 6276 4490 6328 4496
rect 6288 4457 6316 4490
rect 6274 4448 6330 4457
rect 6274 4383 6330 4392
rect 6826 4312 6882 4321
rect 6826 4247 6882 4256
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6380 2854 6408 3674
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 5552 2746 5672 2774
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5448 2576 5500 2582
rect 5448 2518 5500 2524
rect 5460 2394 5488 2518
rect 5552 2514 5580 2586
rect 5644 2514 5672 2746
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5460 2378 5764 2394
rect 5460 2372 5776 2378
rect 5460 2366 5724 2372
rect 5724 2314 5776 2320
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 4712 2032 4764 2038
rect 4712 1974 4764 1980
rect 4528 1964 4580 1970
rect 4528 1906 4580 1912
rect 3056 1828 3108 1834
rect 3056 1770 3108 1776
rect 6564 1766 6592 3334
rect 6656 3058 6684 3470
rect 6840 3194 6868 4247
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6552 1760 6604 1766
rect 6552 1702 6604 1708
rect 7024 1426 7052 5170
rect 7196 5092 7248 5098
rect 7196 5034 7248 5040
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 7116 4622 7144 4966
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 7208 3602 7236 5034
rect 7760 4622 7788 5510
rect 7852 5234 7880 5714
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7300 4146 7328 4422
rect 7668 4185 7696 4422
rect 7654 4176 7710 4185
rect 7288 4140 7340 4146
rect 7654 4111 7710 4120
rect 7288 4082 7340 4088
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7116 2774 7144 3470
rect 7208 3058 7236 3538
rect 7300 3194 7328 4082
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 7196 3052 7248 3058
rect 7248 3012 7328 3040
rect 7196 2994 7248 3000
rect 7116 2746 7236 2774
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7116 2378 7144 2518
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7208 1494 7236 2746
rect 7300 2650 7328 3012
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7392 2446 7420 3062
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7286 2000 7342 2009
rect 7286 1935 7342 1944
rect 7196 1488 7248 1494
rect 7196 1430 7248 1436
rect 7012 1420 7064 1426
rect 7012 1362 7064 1368
rect 7300 800 7328 1935
rect 7392 800 7420 2382
rect 7484 800 7512 2790
rect 7576 800 7604 2926
rect 7668 800 7696 3606
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7760 3126 7788 3470
rect 7748 3120 7800 3126
rect 7748 3062 7800 3068
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 7760 1902 7788 2246
rect 7748 1896 7800 1902
rect 7748 1838 7800 1844
rect 7748 1420 7800 1426
rect 7748 1362 7800 1368
rect 7760 800 7788 1362
rect 7852 800 7880 5170
rect 8036 2632 8064 5646
rect 8680 5234 8708 6190
rect 9876 6186 9904 6598
rect 15398 6556 15706 6565
rect 15398 6554 15404 6556
rect 15460 6554 15484 6556
rect 15540 6554 15564 6556
rect 15620 6554 15644 6556
rect 15700 6554 15706 6556
rect 15460 6502 15462 6554
rect 15642 6502 15644 6554
rect 15398 6500 15404 6502
rect 15460 6500 15484 6502
rect 15540 6500 15564 6502
rect 15620 6500 15644 6502
rect 15700 6500 15706 6502
rect 15398 6491 15706 6500
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 8772 5234 8800 6054
rect 9324 5710 9352 6054
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 8174 4924 8482 4933
rect 8174 4922 8180 4924
rect 8236 4922 8260 4924
rect 8316 4922 8340 4924
rect 8396 4922 8420 4924
rect 8476 4922 8482 4924
rect 8236 4870 8238 4922
rect 8418 4870 8420 4922
rect 8174 4868 8180 4870
rect 8236 4868 8260 4870
rect 8316 4868 8340 4870
rect 8396 4868 8420 4870
rect 8476 4868 8482 4870
rect 8174 4859 8482 4868
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8312 4593 8340 4626
rect 8298 4584 8354 4593
rect 8298 4519 8354 4528
rect 8392 3936 8444 3942
rect 8444 3896 8616 3924
rect 8392 3878 8444 3884
rect 8174 3836 8482 3845
rect 8174 3834 8180 3836
rect 8236 3834 8260 3836
rect 8316 3834 8340 3836
rect 8396 3834 8420 3836
rect 8476 3834 8482 3836
rect 8236 3782 8238 3834
rect 8418 3782 8420 3834
rect 8174 3780 8180 3782
rect 8236 3780 8260 3782
rect 8316 3780 8340 3782
rect 8396 3780 8420 3782
rect 8476 3780 8482 3782
rect 8174 3771 8482 3780
rect 8588 3602 8616 3896
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8312 2990 8340 3334
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8174 2748 8482 2757
rect 8174 2746 8180 2748
rect 8236 2746 8260 2748
rect 8316 2746 8340 2748
rect 8396 2746 8420 2748
rect 8476 2746 8482 2748
rect 8236 2694 8238 2746
rect 8418 2694 8420 2746
rect 8174 2692 8180 2694
rect 8236 2692 8260 2694
rect 8316 2692 8340 2694
rect 8396 2692 8420 2694
rect 8476 2692 8482 2694
rect 8174 2683 8482 2692
rect 8036 2604 8156 2632
rect 7932 1488 7984 1494
rect 7932 1430 7984 1436
rect 7944 800 7972 1430
rect 8024 1352 8076 1358
rect 8024 1294 8076 1300
rect 8036 800 8064 1294
rect 8128 800 8156 2604
rect 8208 1828 8260 1834
rect 8208 1770 8260 1776
rect 8220 800 8248 1770
rect 8588 1578 8616 2790
rect 8404 1550 8616 1578
rect 8404 800 8432 1550
rect 8680 1442 8708 5170
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8772 3233 8800 4014
rect 8852 4004 8904 4010
rect 8852 3946 8904 3952
rect 8864 3738 8892 3946
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8852 3732 8904 3738
rect 8852 3674 8904 3680
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8758 3224 8814 3233
rect 8758 3159 8814 3168
rect 8758 3088 8814 3097
rect 8758 3023 8760 3032
rect 8812 3023 8814 3032
rect 8760 2994 8812 3000
rect 8864 2514 8892 3538
rect 8956 2922 8984 3878
rect 8944 2916 8996 2922
rect 8944 2858 8996 2864
rect 8852 2508 8904 2514
rect 8852 2450 8904 2456
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 8588 1414 8708 1442
rect 8588 800 8616 1414
rect 8772 800 8800 2246
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 8956 800 8984 2042
rect 9140 800 9168 4082
rect 9232 3942 9260 5170
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 9232 2446 9260 2858
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9232 1426 9260 2246
rect 9220 1420 9272 1426
rect 9220 1362 9272 1368
rect 9324 800 9352 5646
rect 9508 5234 9536 6054
rect 9876 5642 9904 6122
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 10520 5914 10548 6054
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 9864 5636 9916 5642
rect 9864 5578 9916 5584
rect 9876 5370 9904 5578
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9404 4684 9456 4690
rect 9404 4626 9456 4632
rect 9416 3754 9444 4626
rect 9508 4026 9536 5170
rect 9678 4720 9734 4729
rect 9876 4690 9904 5306
rect 9678 4655 9734 4664
rect 9864 4684 9916 4690
rect 9692 4554 9720 4655
rect 9864 4626 9916 4632
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9600 4146 9628 4422
rect 9876 4146 9904 4626
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9968 4282 9996 4558
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9508 3998 9904 4026
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9416 3726 9536 3754
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9416 1737 9444 2926
rect 9402 1728 9458 1737
rect 9402 1663 9458 1672
rect 9508 800 9536 3726
rect 9600 800 9628 3878
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9692 3369 9720 3402
rect 9678 3360 9734 3369
rect 9678 3295 9734 3304
rect 9784 800 9812 3674
rect 9876 800 9904 3998
rect 10060 800 10088 5646
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10244 4622 10272 4966
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10152 800 10180 3130
rect 10244 2990 10272 3470
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10336 800 10364 4694
rect 10520 4078 10548 5850
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 10600 5024 10652 5030
rect 10600 4966 10652 4972
rect 10508 4072 10560 4078
rect 10508 4014 10560 4020
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10428 2650 10456 3402
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10520 2582 10548 3470
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10520 2106 10548 2518
rect 10508 2100 10560 2106
rect 10508 2042 10560 2048
rect 10612 800 10640 4966
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10796 3738 10824 4082
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10692 3392 10744 3398
rect 10692 3334 10744 3340
rect 10704 1834 10732 3334
rect 10784 2848 10836 2854
rect 10782 2816 10784 2825
rect 10836 2816 10838 2825
rect 10782 2751 10838 2760
rect 10692 1828 10744 1834
rect 10692 1770 10744 1776
rect 10888 800 10916 5646
rect 11796 5228 11848 5234
rect 11796 5170 11848 5176
rect 11058 5128 11114 5137
rect 11058 5063 11114 5072
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10980 3942 11008 4966
rect 11072 4010 11100 5063
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11532 4078 11560 4490
rect 11716 4078 11744 4762
rect 11808 4758 11836 5170
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11808 4146 11836 4694
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11992 4146 12020 4422
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 11152 2032 11204 2038
rect 11152 1974 11204 1980
rect 11164 800 11192 1974
rect 11440 800 11468 3878
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11624 3194 11652 3334
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11704 3120 11756 3126
rect 11704 3062 11756 3068
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11624 2310 11652 2586
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11716 800 11744 3062
rect 12084 2774 12112 5646
rect 12716 5296 12768 5302
rect 12360 5222 12572 5250
rect 12716 5238 12768 5244
rect 12360 5166 12388 5222
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12176 3913 12204 4082
rect 12162 3904 12218 3913
rect 12162 3839 12218 3848
rect 12176 3602 12204 3839
rect 12346 3632 12402 3641
rect 12164 3596 12216 3602
rect 12346 3567 12348 3576
rect 12164 3538 12216 3544
rect 12400 3567 12402 3576
rect 12348 3538 12400 3544
rect 12164 3392 12216 3398
rect 12164 3334 12216 3340
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 11992 2746 12112 2774
rect 11992 800 12020 2746
rect 12176 1873 12204 3334
rect 12268 2854 12296 3334
rect 12348 2984 12400 2990
rect 12348 2926 12400 2932
rect 12256 2848 12308 2854
rect 12256 2790 12308 2796
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12268 2106 12296 2382
rect 12256 2100 12308 2106
rect 12256 2042 12308 2048
rect 12162 1864 12218 1873
rect 12162 1799 12218 1808
rect 12360 1442 12388 2926
rect 12452 2774 12480 5034
rect 12544 3058 12572 5222
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12636 4729 12664 5102
rect 12622 4720 12678 4729
rect 12622 4655 12678 4664
rect 12728 4622 12756 5238
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12636 4146 12664 4490
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12624 3936 12676 3942
rect 12624 3878 12676 3884
rect 12636 3398 12664 3878
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12728 3176 12756 4422
rect 12636 3148 12756 3176
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12636 2854 12664 3148
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 12452 2746 12572 2774
rect 12440 1896 12492 1902
rect 12440 1838 12492 1844
rect 12452 1698 12480 1838
rect 12440 1692 12492 1698
rect 12440 1634 12492 1640
rect 12268 1414 12388 1442
rect 12268 800 12296 1414
rect 12544 800 12572 2746
rect 12624 2508 12676 2514
rect 12624 2450 12676 2456
rect 12636 1902 12664 2450
rect 12728 2446 12756 2994
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12624 1896 12676 1902
rect 12624 1838 12676 1844
rect 12820 800 12848 5646
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 12912 3058 12940 5510
rect 13452 5296 13504 5302
rect 13450 5264 13452 5273
rect 13504 5264 13506 5273
rect 13450 5199 13506 5208
rect 13084 4820 13136 4826
rect 13084 4762 13136 4768
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 13004 4457 13032 4694
rect 12990 4448 13046 4457
rect 12990 4383 13046 4392
rect 13004 3942 13032 4383
rect 13096 4026 13124 4762
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13188 4146 13216 4626
rect 14384 4622 14412 5510
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 14002 4176 14058 4185
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 13096 3998 13216 4026
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13096 3777 13124 3878
rect 13082 3768 13138 3777
rect 13082 3703 13138 3712
rect 13084 3664 13136 3670
rect 13084 3606 13136 3612
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 12912 2446 12940 2994
rect 13004 2990 13032 3470
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 13096 800 13124 3606
rect 13188 3466 13216 3998
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13372 3505 13400 3878
rect 13358 3496 13414 3505
rect 13176 3460 13228 3466
rect 13556 3466 13584 4150
rect 14002 4111 14058 4120
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13740 3670 13768 4014
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13910 3632 13966 3641
rect 13358 3431 13414 3440
rect 13544 3460 13596 3466
rect 13176 3402 13228 3408
rect 13544 3402 13596 3408
rect 13188 2310 13216 3402
rect 13266 3224 13322 3233
rect 13556 3194 13584 3402
rect 13740 3194 13768 3606
rect 13910 3567 13912 3576
rect 13964 3567 13966 3576
rect 13912 3538 13964 3544
rect 13266 3159 13322 3168
rect 13360 3188 13412 3194
rect 13280 3058 13308 3159
rect 13360 3130 13412 3136
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13372 3058 13400 3130
rect 14016 3058 14044 4111
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 13360 3052 13412 3058
rect 13360 2994 13412 3000
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 13280 2650 13308 2994
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 13372 2446 13400 2790
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13556 1170 13584 2994
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13372 1142 13584 1170
rect 13372 800 13400 1142
rect 13648 800 13676 2926
rect 13832 2038 13860 2926
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13820 2032 13872 2038
rect 13820 1974 13872 1980
rect 13924 800 13952 2858
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14016 2378 14044 2586
rect 14108 2582 14136 3470
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 14004 2372 14056 2378
rect 14004 2314 14056 2320
rect 14200 800 14228 4558
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14384 2854 14412 3674
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14476 800 14504 4966
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 14568 2990 14596 3470
rect 14556 2984 14608 2990
rect 14556 2926 14608 2932
rect 14752 800 14780 5646
rect 15398 5468 15706 5477
rect 15398 5466 15404 5468
rect 15460 5466 15484 5468
rect 15540 5466 15564 5468
rect 15620 5466 15644 5468
rect 15700 5466 15706 5468
rect 15460 5414 15462 5466
rect 15642 5414 15644 5466
rect 15398 5412 15404 5414
rect 15460 5412 15484 5414
rect 15540 5412 15564 5414
rect 15620 5412 15644 5414
rect 15700 5412 15706 5414
rect 15398 5403 15706 5412
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15028 800 15056 4966
rect 15384 4616 15436 4622
rect 15304 4576 15384 4604
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15120 3942 15148 4082
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 15120 3534 15148 3878
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15212 3126 15240 4422
rect 15304 4282 15332 4576
rect 15384 4558 15436 4564
rect 15398 4380 15706 4389
rect 15398 4378 15404 4380
rect 15460 4378 15484 4380
rect 15540 4378 15564 4380
rect 15620 4378 15644 4380
rect 15700 4378 15706 4380
rect 15460 4326 15462 4378
rect 15642 4326 15644 4378
rect 15398 4324 15404 4326
rect 15460 4324 15484 4326
rect 15540 4324 15564 4326
rect 15620 4324 15644 4326
rect 15700 4324 15706 4326
rect 15398 4315 15706 4324
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15200 3120 15252 3126
rect 15200 3062 15252 3068
rect 15304 2990 15332 4082
rect 15396 3738 15424 4218
rect 15658 4176 15714 4185
rect 15568 4140 15620 4146
rect 15658 4111 15714 4120
rect 15568 4082 15620 4088
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15580 3466 15608 4082
rect 15672 3602 15700 4111
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15398 3292 15706 3301
rect 15398 3290 15404 3292
rect 15460 3290 15484 3292
rect 15540 3290 15564 3292
rect 15620 3290 15644 3292
rect 15700 3290 15706 3292
rect 15460 3238 15462 3290
rect 15642 3238 15644 3290
rect 15398 3236 15404 3238
rect 15460 3236 15484 3238
rect 15540 3236 15564 3238
rect 15620 3236 15644 3238
rect 15700 3236 15706 3238
rect 15398 3227 15706 3236
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15568 2848 15620 2854
rect 15290 2816 15346 2825
rect 15568 2790 15620 2796
rect 15290 2751 15346 2760
rect 15304 800 15332 2751
rect 15580 2514 15608 2790
rect 15672 2774 15700 3130
rect 15764 3058 15792 4966
rect 15844 4548 15896 4554
rect 15844 4490 15896 4496
rect 15856 4162 15884 4490
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15948 4282 15976 4422
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15856 4134 15976 4162
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15672 2746 15792 2774
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15398 2204 15706 2213
rect 15398 2202 15404 2204
rect 15460 2202 15484 2204
rect 15540 2202 15564 2204
rect 15620 2202 15644 2204
rect 15700 2202 15706 2204
rect 15460 2150 15462 2202
rect 15642 2150 15644 2202
rect 15398 2148 15404 2150
rect 15460 2148 15484 2150
rect 15540 2148 15564 2150
rect 15620 2148 15644 2150
rect 15700 2148 15706 2150
rect 15398 2139 15706 2148
rect 15764 1442 15792 2746
rect 15580 1414 15792 1442
rect 15580 800 15608 1414
rect 15856 800 15884 3130
rect 15948 800 15976 4134
rect 16040 2774 16068 5034
rect 16120 4752 16172 4758
rect 16120 4694 16172 4700
rect 16132 4554 16160 4694
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16132 3602 16160 4082
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 16040 2746 16160 2774
rect 16132 800 16160 2746
rect 16224 800 16252 5646
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16316 3058 16344 5510
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16500 4146 16528 5102
rect 16776 5030 16804 5170
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16408 3194 16436 4014
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16396 2984 16448 2990
rect 16396 2926 16448 2932
rect 16408 800 16436 2926
rect 16488 2644 16540 2650
rect 16488 2586 16540 2592
rect 16500 800 16528 2586
rect 16684 800 16712 4626
rect 16776 800 16804 4966
rect 16960 800 16988 5646
rect 20732 5574 20760 6054
rect 20824 5914 20852 6190
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 25136 6112 25188 6118
rect 25136 6054 25188 6060
rect 26976 6112 27028 6118
rect 26976 6054 27028 6060
rect 22622 6012 22930 6021
rect 22622 6010 22628 6012
rect 22684 6010 22708 6012
rect 22764 6010 22788 6012
rect 22844 6010 22868 6012
rect 22924 6010 22930 6012
rect 22684 5958 22686 6010
rect 22866 5958 22868 6010
rect 22622 5956 22628 5958
rect 22684 5956 22708 5958
rect 22764 5956 22788 5958
rect 22844 5956 22868 5958
rect 22924 5956 22930 5958
rect 22622 5947 22930 5956
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 20720 5568 20772 5574
rect 20720 5510 20772 5516
rect 19248 5364 19300 5370
rect 19248 5306 19300 5312
rect 18328 5296 18380 5302
rect 18328 5238 18380 5244
rect 17960 5228 18012 5234
rect 17960 5170 18012 5176
rect 17592 5092 17644 5098
rect 17592 5034 17644 5040
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17144 800 17172 4966
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 17420 800 17448 4626
rect 17604 4622 17632 5034
rect 17592 4616 17644 4622
rect 17590 4584 17592 4593
rect 17644 4584 17646 4593
rect 17972 4554 18000 5170
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18052 4752 18104 4758
rect 18156 4729 18184 4762
rect 18052 4694 18104 4700
rect 18142 4720 18198 4729
rect 18064 4604 18092 4694
rect 18340 4690 18368 5238
rect 19156 5092 19208 5098
rect 19156 5034 19208 5040
rect 18972 5024 19024 5030
rect 18972 4966 19024 4972
rect 18984 4826 19012 4966
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 18142 4655 18198 4664
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18420 4616 18472 4622
rect 18064 4576 18184 4604
rect 17590 4519 17646 4528
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17972 4282 18000 4490
rect 17960 4276 18012 4282
rect 17960 4218 18012 4224
rect 17972 4078 18000 4218
rect 17960 4072 18012 4078
rect 17866 4040 17922 4049
rect 17960 4014 18012 4020
rect 17866 3975 17922 3984
rect 17880 3942 17908 3975
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17592 3732 17644 3738
rect 17868 3732 17920 3738
rect 17644 3692 17724 3720
rect 17592 3674 17644 3680
rect 17696 800 17724 3692
rect 17868 3674 17920 3680
rect 17880 3398 17908 3674
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17972 800 18000 3878
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18064 3194 18092 3538
rect 18156 3466 18184 4576
rect 18420 4558 18472 4564
rect 18432 4146 18460 4558
rect 19062 4176 19118 4185
rect 18420 4140 18472 4146
rect 18472 4100 18552 4128
rect 19062 4111 19118 4120
rect 18420 4082 18472 4088
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3738 18276 3878
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18340 3602 18368 4014
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 18524 3534 18552 4100
rect 19076 4078 19104 4111
rect 19064 4072 19116 4078
rect 19064 4014 19116 4020
rect 19168 3738 19196 5034
rect 19260 4690 19288 5306
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19260 4282 19288 4626
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18144 3460 18196 3466
rect 18144 3402 18196 3408
rect 18328 3460 18380 3466
rect 18328 3402 18380 3408
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 18156 1766 18184 3402
rect 18340 3058 18368 3402
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 18328 2440 18380 2446
rect 18328 2382 18380 2388
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 18144 1760 18196 1766
rect 18144 1702 18196 1708
rect 18248 800 18276 2042
rect 18340 2038 18368 2382
rect 18432 2106 18460 2450
rect 18420 2100 18472 2106
rect 18420 2042 18472 2048
rect 18328 2032 18380 2038
rect 18328 1974 18380 1980
rect 18524 800 18552 3130
rect 19260 3058 19288 4218
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 19352 3913 19380 4150
rect 19338 3904 19394 3913
rect 19338 3839 19394 3848
rect 19616 3664 19668 3670
rect 19616 3606 19668 3612
rect 19248 3052 19300 3058
rect 19248 2994 19300 3000
rect 18602 2952 18658 2961
rect 18602 2887 18658 2896
rect 19340 2916 19392 2922
rect 18616 1902 18644 2887
rect 19340 2858 19392 2864
rect 19064 2576 19116 2582
rect 19064 2518 19116 2524
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 18604 1896 18656 1902
rect 18604 1838 18656 1844
rect 18800 800 18828 2246
rect 19076 800 19104 2518
rect 19352 800 19380 2858
rect 19628 800 19656 3606
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 19720 3505 19748 3538
rect 19706 3496 19762 3505
rect 19706 3431 19762 3440
rect 19800 3392 19852 3398
rect 19800 3334 19852 3340
rect 19812 3194 19840 3334
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 19812 3097 19840 3130
rect 19798 3088 19854 3097
rect 19798 3023 19854 3032
rect 19904 800 19932 4966
rect 19996 3398 20024 5510
rect 20732 5370 20760 5510
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20824 5302 20852 5850
rect 22744 5636 22796 5642
rect 22744 5578 22796 5584
rect 21640 5568 21692 5574
rect 21640 5510 21692 5516
rect 22468 5568 22520 5574
rect 22468 5510 22520 5516
rect 20812 5296 20864 5302
rect 20812 5238 20864 5244
rect 21180 5296 21232 5302
rect 21180 5238 21232 5244
rect 21192 4146 21220 5238
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 20720 4072 20772 4078
rect 20718 4040 20720 4049
rect 20772 4040 20774 4049
rect 20718 3975 20774 3984
rect 21088 3936 21140 3942
rect 21088 3878 21140 3884
rect 21100 3466 21128 3878
rect 21192 3602 21220 4082
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19996 3097 20024 3334
rect 19982 3088 20038 3097
rect 19982 3023 20038 3032
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20168 2032 20220 2038
rect 20168 1974 20220 1980
rect 20180 800 20208 1974
rect 20456 800 20484 2994
rect 20996 2916 21048 2922
rect 20996 2858 21048 2864
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20732 800 20760 2586
rect 21008 800 21036 2858
rect 21284 800 21312 4558
rect 21652 3534 21680 5510
rect 22192 5160 22244 5166
rect 22192 5102 22244 5108
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22112 4758 22140 4966
rect 22100 4752 22152 4758
rect 22100 4694 22152 4700
rect 22204 4146 22232 5102
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21548 2100 21600 2106
rect 21548 2042 21600 2048
rect 21560 800 21588 2042
rect 21652 1698 21680 3470
rect 21732 3392 21784 3398
rect 21732 3334 21784 3340
rect 21744 3233 21772 3334
rect 21730 3224 21786 3233
rect 21730 3159 21786 3168
rect 21744 2961 21772 3159
rect 21730 2952 21786 2961
rect 21730 2887 21786 2896
rect 21640 1692 21692 1698
rect 21640 1634 21692 1640
rect 21836 800 21864 3878
rect 22020 3738 22048 4082
rect 22008 3732 22060 3738
rect 22008 3674 22060 3680
rect 22480 2446 22508 5510
rect 22756 5302 22784 5578
rect 23020 5568 23072 5574
rect 23020 5510 23072 5516
rect 22744 5296 22796 5302
rect 22744 5238 22796 5244
rect 23032 5030 23060 5510
rect 23020 5024 23072 5030
rect 23018 4992 23020 5001
rect 23072 4992 23074 5001
rect 22622 4924 22930 4933
rect 23018 4927 23074 4936
rect 22622 4922 22628 4924
rect 22684 4922 22708 4924
rect 22764 4922 22788 4924
rect 22844 4922 22868 4924
rect 22924 4922 22930 4924
rect 22684 4870 22686 4922
rect 22866 4870 22868 4922
rect 23032 4901 23060 4927
rect 22622 4868 22628 4870
rect 22684 4868 22708 4870
rect 22764 4868 22788 4870
rect 22844 4868 22868 4870
rect 22924 4868 22930 4870
rect 22622 4859 22930 4868
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22572 4010 22600 4558
rect 22756 4282 22784 4558
rect 22744 4276 22796 4282
rect 22744 4218 22796 4224
rect 22560 4004 22612 4010
rect 22560 3946 22612 3952
rect 23204 3936 23256 3942
rect 23204 3878 23256 3884
rect 22622 3836 22930 3845
rect 22622 3834 22628 3836
rect 22684 3834 22708 3836
rect 22764 3834 22788 3836
rect 22844 3834 22868 3836
rect 22924 3834 22930 3836
rect 22684 3782 22686 3834
rect 22866 3782 22868 3834
rect 22622 3780 22628 3782
rect 22684 3780 22708 3782
rect 22764 3780 22788 3782
rect 22844 3780 22868 3782
rect 22924 3780 22930 3782
rect 22622 3771 22930 3780
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 22622 2748 22930 2757
rect 22622 2746 22628 2748
rect 22684 2746 22708 2748
rect 22764 2746 22788 2748
rect 22844 2746 22868 2748
rect 22924 2746 22930 2748
rect 22684 2694 22686 2746
rect 22866 2694 22868 2746
rect 22622 2692 22628 2694
rect 22684 2692 22708 2694
rect 22764 2692 22788 2694
rect 22844 2692 22868 2694
rect 22924 2692 22930 2694
rect 22622 2683 22930 2692
rect 22652 2576 22704 2582
rect 22652 2518 22704 2524
rect 22284 2440 22336 2446
rect 22468 2440 22520 2446
rect 22336 2400 22416 2428
rect 22284 2382 22336 2388
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 22112 800 22140 2314
rect 22388 800 22416 2400
rect 22468 2382 22520 2388
rect 22480 1766 22508 2382
rect 22468 1760 22520 1766
rect 22468 1702 22520 1708
rect 22664 800 22692 2518
rect 22928 2508 22980 2514
rect 22928 2450 22980 2456
rect 22940 800 22968 2450
rect 23124 1902 23152 3470
rect 23112 1896 23164 1902
rect 23112 1838 23164 1844
rect 23216 800 23244 3878
rect 23308 2446 23336 6054
rect 25148 5574 25176 6054
rect 26792 5704 26844 5710
rect 26792 5646 26844 5652
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 24768 5568 24820 5574
rect 24768 5510 24820 5516
rect 25136 5568 25188 5574
rect 25136 5510 25188 5516
rect 25228 5568 25280 5574
rect 25228 5510 25280 5516
rect 26700 5568 26752 5574
rect 26700 5510 26752 5516
rect 23388 5296 23440 5302
rect 23388 5238 23440 5244
rect 23400 4758 23428 5238
rect 23388 4752 23440 4758
rect 23388 4694 23440 4700
rect 23492 4298 23520 5510
rect 24124 5364 24176 5370
rect 24124 5306 24176 5312
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 23400 4270 23520 4298
rect 23400 3534 23428 4270
rect 23480 4208 23532 4214
rect 23480 4150 23532 4156
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23308 2038 23336 2382
rect 23296 2032 23348 2038
rect 23492 2009 23520 4150
rect 23860 4146 23888 4966
rect 24136 4146 24164 5306
rect 24780 5166 24808 5510
rect 25148 5370 25176 5510
rect 25136 5364 25188 5370
rect 25136 5306 25188 5312
rect 24768 5160 24820 5166
rect 24768 5102 24820 5108
rect 25044 5160 25096 5166
rect 25044 5102 25096 5108
rect 24584 5092 24636 5098
rect 24584 5034 24636 5040
rect 24596 4622 24624 5034
rect 24216 4616 24268 4622
rect 24216 4558 24268 4564
rect 24584 4616 24636 4622
rect 24584 4558 24636 4564
rect 23848 4140 23900 4146
rect 23848 4082 23900 4088
rect 24124 4140 24176 4146
rect 24124 4082 24176 4088
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23296 1974 23348 1980
rect 23478 2000 23534 2009
rect 23478 1935 23534 1944
rect 23584 898 23612 3334
rect 23860 2922 23888 4082
rect 24136 3194 24164 4082
rect 24228 3924 24256 4558
rect 24780 4162 24808 5102
rect 24952 5024 25004 5030
rect 24952 4966 25004 4972
rect 24964 4185 24992 4966
rect 25056 4758 25084 5102
rect 25044 4752 25096 4758
rect 25044 4694 25096 4700
rect 25148 4690 25176 5306
rect 25240 5302 25268 5510
rect 25780 5364 25832 5370
rect 25780 5306 25832 5312
rect 25228 5296 25280 5302
rect 25228 5238 25280 5244
rect 25320 5228 25372 5234
rect 25320 5170 25372 5176
rect 25136 4684 25188 4690
rect 25136 4626 25188 4632
rect 24950 4176 25006 4185
rect 24780 4134 24900 4162
rect 24872 4049 24900 4134
rect 24950 4111 25006 4120
rect 24858 4040 24914 4049
rect 24858 3975 24914 3984
rect 24308 3936 24360 3942
rect 24228 3896 24308 3924
rect 24124 3188 24176 3194
rect 24124 3130 24176 3136
rect 23756 2916 23808 2922
rect 23756 2858 23808 2864
rect 23848 2916 23900 2922
rect 23848 2858 23900 2864
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 23676 1698 23704 2382
rect 23664 1692 23716 1698
rect 23664 1634 23716 1640
rect 23492 870 23612 898
rect 23492 800 23520 870
rect 23768 800 23796 2858
rect 24032 2848 24084 2854
rect 24032 2790 24084 2796
rect 24044 800 24072 2790
rect 24228 2514 24256 3896
rect 24308 3878 24360 3884
rect 25332 3738 25360 5170
rect 25792 4622 25820 5306
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 26148 4480 26200 4486
rect 26148 4422 26200 4428
rect 25502 4040 25558 4049
rect 25502 3975 25504 3984
rect 25556 3975 25558 3984
rect 25778 4040 25834 4049
rect 25778 3975 25834 3984
rect 25504 3946 25556 3952
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 24584 3664 24636 3670
rect 24584 3606 24636 3612
rect 24308 3392 24360 3398
rect 24308 3334 24360 3340
rect 24216 2508 24268 2514
rect 24216 2450 24268 2456
rect 24320 800 24348 3334
rect 24596 3074 24624 3606
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 24688 3194 24716 3470
rect 24860 3460 24912 3466
rect 24860 3402 24912 3408
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24596 3058 24716 3074
rect 24872 3058 24900 3402
rect 25688 3392 25740 3398
rect 25688 3334 25740 3340
rect 24596 3052 24728 3058
rect 24596 3046 24676 3052
rect 24676 2994 24728 3000
rect 24860 3052 24912 3058
rect 24860 2994 24912 3000
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 24504 2310 24532 2926
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 24492 2304 24544 2310
rect 24492 2246 24544 2252
rect 24596 800 24624 2586
rect 24688 2514 24716 2994
rect 25136 2576 25188 2582
rect 25136 2518 25188 2524
rect 24676 2508 24728 2514
rect 24676 2450 24728 2456
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 24780 1834 24808 2450
rect 24860 2372 24912 2378
rect 24860 2314 24912 2320
rect 24768 1828 24820 1834
rect 24768 1770 24820 1776
rect 24872 800 24900 2314
rect 25148 800 25176 2518
rect 25596 2304 25648 2310
rect 25596 2246 25648 2252
rect 25608 1970 25636 2246
rect 25596 1964 25648 1970
rect 25596 1906 25648 1912
rect 25412 1420 25464 1426
rect 25412 1362 25464 1368
rect 25424 800 25452 1362
rect 25700 800 25728 3334
rect 25792 2310 25820 3975
rect 26160 3602 26188 4422
rect 26332 4140 26384 4146
rect 26332 4082 26384 4088
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 26056 3528 26108 3534
rect 26054 3496 26056 3505
rect 26108 3496 26110 3505
rect 26054 3431 26110 3440
rect 26240 3392 26292 3398
rect 26240 3334 26292 3340
rect 25964 2848 26016 2854
rect 25964 2790 26016 2796
rect 25780 2304 25832 2310
rect 25780 2246 25832 2252
rect 25976 800 26004 2790
rect 26252 800 26280 3334
rect 26344 2378 26372 4082
rect 26424 3936 26476 3942
rect 26424 3878 26476 3884
rect 26436 3670 26464 3878
rect 26424 3664 26476 3670
rect 26424 3606 26476 3612
rect 26712 3534 26740 5510
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 26608 3052 26660 3058
rect 26608 2994 26660 3000
rect 26516 2848 26568 2854
rect 26516 2790 26568 2796
rect 26332 2372 26384 2378
rect 26332 2314 26384 2320
rect 26528 800 26556 2790
rect 26620 2582 26648 2994
rect 26712 2961 26740 3470
rect 26698 2952 26754 2961
rect 26698 2887 26754 2896
rect 26712 2650 26740 2887
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 26608 2576 26660 2582
rect 26608 2518 26660 2524
rect 26804 800 26832 5646
rect 26884 5568 26936 5574
rect 26884 5510 26936 5516
rect 26896 4690 26924 5510
rect 26988 5234 27016 6054
rect 26976 5228 27028 5234
rect 26976 5170 27028 5176
rect 26884 4684 26936 4690
rect 26884 4626 26936 4632
rect 26988 3602 27016 5170
rect 27160 5024 27212 5030
rect 27160 4966 27212 4972
rect 26976 3596 27028 3602
rect 26976 3538 27028 3544
rect 26884 2916 26936 2922
rect 26884 2858 26936 2864
rect 26896 2553 26924 2858
rect 26882 2544 26938 2553
rect 26988 2514 27016 3538
rect 27172 2530 27200 4966
rect 27250 3088 27306 3097
rect 27356 3058 27384 6666
rect 33508 6656 33560 6662
rect 33508 6598 33560 6604
rect 29846 6556 30154 6565
rect 29846 6554 29852 6556
rect 29908 6554 29932 6556
rect 29988 6554 30012 6556
rect 30068 6554 30092 6556
rect 30148 6554 30154 6556
rect 29908 6502 29910 6554
rect 30090 6502 30092 6554
rect 29846 6500 29852 6502
rect 29908 6500 29932 6502
rect 29988 6500 30012 6502
rect 30068 6500 30092 6502
rect 30148 6500 30154 6502
rect 29846 6491 30154 6500
rect 30288 6248 30340 6254
rect 30288 6190 30340 6196
rect 28264 6112 28316 6118
rect 28264 6054 28316 6060
rect 27712 5840 27764 5846
rect 27712 5782 27764 5788
rect 27620 5772 27672 5778
rect 27620 5714 27672 5720
rect 27250 3023 27306 3032
rect 27344 3052 27396 3058
rect 26882 2479 26938 2488
rect 26976 2508 27028 2514
rect 26976 2450 27028 2456
rect 27080 2502 27200 2530
rect 27080 800 27108 2502
rect 27264 2417 27292 3023
rect 27344 2994 27396 3000
rect 27632 2774 27660 5714
rect 27356 2746 27660 2774
rect 27250 2408 27306 2417
rect 27250 2343 27306 2352
rect 27356 800 27384 2746
rect 27724 2666 27752 5782
rect 28172 5296 28224 5302
rect 28172 5238 28224 5244
rect 27896 3936 27948 3942
rect 27896 3878 27948 3884
rect 27632 2638 27752 2666
rect 27528 2372 27580 2378
rect 27528 2314 27580 2320
rect 27540 1426 27568 2314
rect 27528 1420 27580 1426
rect 27528 1362 27580 1368
rect 27632 800 27660 2638
rect 27908 800 27936 3878
rect 28184 800 28212 5238
rect 28276 4729 28304 6054
rect 29736 5704 29788 5710
rect 29736 5646 29788 5652
rect 28816 5568 28868 5574
rect 28816 5510 28868 5516
rect 29460 5568 29512 5574
rect 29460 5510 29512 5516
rect 28448 5024 28500 5030
rect 28448 4966 28500 4972
rect 28262 4720 28318 4729
rect 28262 4655 28318 4664
rect 28276 4622 28304 4655
rect 28264 4616 28316 4622
rect 28264 4558 28316 4564
rect 28276 3233 28304 4558
rect 28262 3224 28318 3233
rect 28262 3159 28318 3168
rect 28356 2304 28408 2310
rect 28356 2246 28408 2252
rect 28368 1737 28396 2246
rect 28354 1728 28410 1737
rect 28354 1663 28410 1672
rect 28460 800 28488 4966
rect 28724 4616 28776 4622
rect 28724 4558 28776 4564
rect 28632 3936 28684 3942
rect 28632 3878 28684 3884
rect 28644 3126 28672 3878
rect 28632 3120 28684 3126
rect 28632 3062 28684 3068
rect 28736 800 28764 4558
rect 28828 4214 28856 5510
rect 29472 5166 29500 5510
rect 29552 5364 29604 5370
rect 29552 5306 29604 5312
rect 29460 5160 29512 5166
rect 29460 5102 29512 5108
rect 29472 4758 29500 5102
rect 29460 4752 29512 4758
rect 29460 4694 29512 4700
rect 29564 4690 29592 5306
rect 29748 5098 29776 5646
rect 29846 5468 30154 5477
rect 29846 5466 29852 5468
rect 29908 5466 29932 5468
rect 29988 5466 30012 5468
rect 30068 5466 30092 5468
rect 30148 5466 30154 5468
rect 29908 5414 29910 5466
rect 30090 5414 30092 5466
rect 29846 5412 29852 5414
rect 29908 5412 29932 5414
rect 29988 5412 30012 5414
rect 30068 5412 30092 5414
rect 30148 5412 30154 5414
rect 29846 5403 30154 5412
rect 30300 5166 30328 6190
rect 33520 6186 33548 6598
rect 44294 6556 44602 6565
rect 44294 6554 44300 6556
rect 44356 6554 44380 6556
rect 44436 6554 44460 6556
rect 44516 6554 44540 6556
rect 44596 6554 44602 6556
rect 44356 6502 44358 6554
rect 44538 6502 44540 6554
rect 44294 6500 44300 6502
rect 44356 6500 44380 6502
rect 44436 6500 44460 6502
rect 44516 6500 44540 6502
rect 44596 6500 44602 6502
rect 44294 6491 44602 6500
rect 38384 6248 38436 6254
rect 38384 6190 38436 6196
rect 42984 6248 43036 6254
rect 42984 6190 43036 6196
rect 33508 6180 33560 6186
rect 33508 6122 33560 6128
rect 30472 6112 30524 6118
rect 30472 6054 30524 6060
rect 31760 6112 31812 6118
rect 31760 6054 31812 6060
rect 33232 6112 33284 6118
rect 33232 6054 33284 6060
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30392 5273 30420 5510
rect 30378 5264 30434 5273
rect 30378 5199 30434 5208
rect 30288 5160 30340 5166
rect 30288 5102 30340 5108
rect 29736 5092 29788 5098
rect 29736 5034 29788 5040
rect 30286 4992 30342 5001
rect 30484 4978 30512 6054
rect 31024 5840 31076 5846
rect 31022 5808 31024 5817
rect 31076 5808 31078 5817
rect 31022 5743 31078 5752
rect 31668 5772 31720 5778
rect 31036 5370 31064 5743
rect 31668 5714 31720 5720
rect 31024 5364 31076 5370
rect 31024 5306 31076 5312
rect 31680 5234 31708 5714
rect 31668 5228 31720 5234
rect 31668 5170 31720 5176
rect 31680 5030 31708 5170
rect 30342 4950 30512 4978
rect 31668 5024 31720 5030
rect 31668 4966 31720 4972
rect 30286 4927 30342 4936
rect 30300 4826 30328 4927
rect 30288 4820 30340 4826
rect 30288 4762 30340 4768
rect 29552 4684 29604 4690
rect 29552 4626 29604 4632
rect 30300 4457 30328 4762
rect 30656 4616 30708 4622
rect 30656 4558 30708 4564
rect 31392 4616 31444 4622
rect 31392 4558 31444 4564
rect 30286 4448 30342 4457
rect 29846 4380 30154 4389
rect 30286 4383 30342 4392
rect 29846 4378 29852 4380
rect 29908 4378 29932 4380
rect 29988 4378 30012 4380
rect 30068 4378 30092 4380
rect 30148 4378 30154 4380
rect 29908 4326 29910 4378
rect 30090 4326 30092 4378
rect 29846 4324 29852 4326
rect 29908 4324 29932 4326
rect 29988 4324 30012 4326
rect 30068 4324 30092 4326
rect 30148 4324 30154 4326
rect 29846 4315 30154 4324
rect 30668 4282 30696 4558
rect 30656 4276 30708 4282
rect 30656 4218 30708 4224
rect 31404 4214 31432 4558
rect 31772 4282 31800 6054
rect 31852 5908 31904 5914
rect 31852 5850 31904 5856
rect 33048 5908 33100 5914
rect 33048 5850 33100 5856
rect 31864 5642 31892 5850
rect 33060 5778 33088 5850
rect 33048 5772 33100 5778
rect 33048 5714 33100 5720
rect 32864 5704 32916 5710
rect 32126 5672 32182 5681
rect 31852 5636 31904 5642
rect 32864 5646 32916 5652
rect 32126 5607 32128 5616
rect 31852 5578 31904 5584
rect 32180 5607 32182 5616
rect 32128 5578 32180 5584
rect 32036 5568 32088 5574
rect 32088 5516 32168 5522
rect 32036 5510 32168 5516
rect 32048 5494 32168 5510
rect 32140 5234 32168 5494
rect 32128 5228 32180 5234
rect 32128 5170 32180 5176
rect 32140 4758 32168 5170
rect 32876 5166 32904 5646
rect 33244 5234 33272 6054
rect 33416 5568 33468 5574
rect 33416 5510 33468 5516
rect 33428 5302 33456 5510
rect 33416 5296 33468 5302
rect 33416 5238 33468 5244
rect 33232 5228 33284 5234
rect 33232 5170 33284 5176
rect 32864 5160 32916 5166
rect 32864 5102 32916 5108
rect 32128 4752 32180 4758
rect 32128 4694 32180 4700
rect 32586 4584 32642 4593
rect 32586 4519 32642 4528
rect 32600 4486 32628 4519
rect 32588 4480 32640 4486
rect 32588 4422 32640 4428
rect 32600 4282 32628 4422
rect 31760 4276 31812 4282
rect 31760 4218 31812 4224
rect 32588 4276 32640 4282
rect 32588 4218 32640 4224
rect 28816 4208 28868 4214
rect 28816 4150 28868 4156
rect 31392 4208 31444 4214
rect 31392 4150 31444 4156
rect 30932 4140 30984 4146
rect 30932 4082 30984 4088
rect 30380 4072 30432 4078
rect 30380 4014 30432 4020
rect 29736 4004 29788 4010
rect 29736 3946 29788 3952
rect 29000 3528 29052 3534
rect 29000 3470 29052 3476
rect 29012 800 29040 3470
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 29104 3058 29132 3334
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 29552 2848 29604 2854
rect 29552 2790 29604 2796
rect 29276 2508 29328 2514
rect 29276 2450 29328 2456
rect 29288 800 29316 2450
rect 29564 800 29592 2790
rect 29748 1986 29776 3946
rect 30392 3602 30420 4014
rect 30944 3738 30972 4082
rect 31404 3942 31432 4150
rect 32600 4146 32628 4218
rect 32588 4140 32640 4146
rect 32588 4082 32640 4088
rect 33416 4140 33468 4146
rect 33520 4128 33548 6122
rect 34612 6112 34664 6118
rect 34612 6054 34664 6060
rect 35072 6112 35124 6118
rect 35072 6054 35124 6060
rect 35716 6112 35768 6118
rect 35716 6054 35768 6060
rect 35808 6112 35860 6118
rect 35808 6054 35860 6060
rect 36268 6112 36320 6118
rect 36268 6054 36320 6060
rect 34624 5846 34652 6054
rect 34704 5908 34756 5914
rect 34704 5850 34756 5856
rect 34612 5840 34664 5846
rect 34716 5817 34744 5850
rect 34612 5782 34664 5788
rect 34702 5808 34758 5817
rect 34702 5743 34758 5752
rect 34888 5772 34940 5778
rect 34888 5714 34940 5720
rect 34152 5704 34204 5710
rect 34152 5646 34204 5652
rect 33966 5536 34022 5545
rect 33966 5471 34022 5480
rect 33876 5228 33928 5234
rect 33876 5170 33928 5176
rect 33888 5137 33916 5170
rect 33980 5166 34008 5471
rect 34164 5234 34192 5646
rect 34152 5228 34204 5234
rect 34152 5170 34204 5176
rect 34900 5166 34928 5714
rect 33968 5160 34020 5166
rect 33874 5128 33930 5137
rect 33968 5102 34020 5108
rect 34888 5160 34940 5166
rect 34888 5102 34940 5108
rect 33874 5063 33930 5072
rect 33888 4622 33916 5063
rect 34336 5024 34388 5030
rect 34336 4966 34388 4972
rect 33876 4616 33928 4622
rect 33876 4558 33928 4564
rect 34348 4282 34376 4966
rect 35084 4622 35112 6054
rect 35728 5914 35756 6054
rect 35532 5908 35584 5914
rect 35716 5908 35768 5914
rect 35532 5850 35584 5856
rect 35636 5868 35716 5896
rect 35544 5710 35572 5850
rect 35532 5704 35584 5710
rect 35532 5646 35584 5652
rect 35348 5636 35400 5642
rect 35348 5578 35400 5584
rect 35360 5234 35388 5578
rect 35348 5228 35400 5234
rect 35348 5170 35400 5176
rect 35440 5024 35492 5030
rect 35440 4966 35492 4972
rect 35452 4690 35480 4966
rect 35636 4826 35664 5868
rect 35716 5850 35768 5856
rect 35820 5778 35848 6054
rect 35808 5772 35860 5778
rect 35808 5714 35860 5720
rect 36280 5710 36308 6054
rect 37070 6012 37378 6021
rect 37070 6010 37076 6012
rect 37132 6010 37156 6012
rect 37212 6010 37236 6012
rect 37292 6010 37316 6012
rect 37372 6010 37378 6012
rect 37132 5958 37134 6010
rect 37314 5958 37316 6010
rect 37070 5956 37076 5958
rect 37132 5956 37156 5958
rect 37212 5956 37236 5958
rect 37292 5956 37316 5958
rect 37372 5956 37378 5958
rect 37070 5947 37378 5956
rect 36268 5704 36320 5710
rect 36268 5646 36320 5652
rect 36452 5704 36504 5710
rect 36452 5646 36504 5652
rect 36464 5545 36492 5646
rect 36450 5536 36506 5545
rect 36450 5471 36506 5480
rect 36728 5228 36780 5234
rect 36728 5170 36780 5176
rect 35808 5160 35860 5166
rect 36740 5137 36768 5170
rect 35808 5102 35860 5108
rect 36726 5128 36782 5137
rect 35820 4826 35848 5102
rect 36726 5063 36782 5072
rect 37556 5024 37608 5030
rect 37556 4966 37608 4972
rect 38200 5024 38252 5030
rect 38200 4966 38252 4972
rect 37070 4924 37378 4933
rect 37070 4922 37076 4924
rect 37132 4922 37156 4924
rect 37212 4922 37236 4924
rect 37292 4922 37316 4924
rect 37372 4922 37378 4924
rect 37132 4870 37134 4922
rect 37314 4870 37316 4922
rect 37070 4868 37076 4870
rect 37132 4868 37156 4870
rect 37212 4868 37236 4870
rect 37292 4868 37316 4870
rect 37372 4868 37378 4870
rect 37070 4859 37378 4868
rect 35624 4820 35676 4826
rect 35624 4762 35676 4768
rect 35808 4820 35860 4826
rect 35808 4762 35860 4768
rect 35440 4684 35492 4690
rect 35440 4626 35492 4632
rect 37568 4622 37596 4966
rect 37646 4720 37702 4729
rect 37646 4655 37702 4664
rect 37660 4622 37688 4655
rect 35072 4616 35124 4622
rect 37556 4616 37608 4622
rect 35072 4558 35124 4564
rect 35438 4584 35494 4593
rect 34428 4548 34480 4554
rect 35728 4554 36032 4570
rect 37556 4558 37608 4564
rect 37648 4616 37700 4622
rect 37648 4558 37700 4564
rect 35438 4519 35494 4528
rect 35716 4548 36032 4554
rect 34428 4490 34480 4496
rect 34336 4276 34388 4282
rect 34336 4218 34388 4224
rect 33468 4100 33548 4128
rect 33416 4082 33468 4088
rect 32772 4004 32824 4010
rect 32772 3946 32824 3952
rect 31392 3936 31444 3942
rect 32784 3913 32812 3946
rect 31392 3878 31444 3884
rect 32770 3904 32826 3913
rect 30932 3732 30984 3738
rect 30932 3674 30984 3680
rect 30380 3596 30432 3602
rect 30380 3538 30432 3544
rect 31208 3596 31260 3602
rect 31208 3538 31260 3544
rect 29846 3292 30154 3301
rect 29846 3290 29852 3292
rect 29908 3290 29932 3292
rect 29988 3290 30012 3292
rect 30068 3290 30092 3292
rect 30148 3290 30154 3292
rect 29908 3238 29910 3290
rect 30090 3238 30092 3290
rect 29846 3236 29852 3238
rect 29908 3236 29932 3238
rect 29988 3236 30012 3238
rect 30068 3236 30092 3238
rect 30148 3236 30154 3238
rect 29846 3227 30154 3236
rect 30392 2990 30420 3538
rect 30484 3398 30512 3429
rect 30472 3392 30524 3398
rect 30470 3360 30472 3369
rect 30524 3360 30526 3369
rect 30470 3295 30526 3304
rect 30380 2984 30432 2990
rect 30380 2926 30432 2932
rect 30196 2848 30248 2854
rect 30196 2790 30248 2796
rect 29846 2204 30154 2213
rect 29846 2202 29852 2204
rect 29908 2202 29932 2204
rect 29988 2202 30012 2204
rect 30068 2202 30092 2204
rect 30148 2202 30154 2204
rect 29908 2150 29910 2202
rect 30090 2150 30092 2202
rect 29846 2148 29852 2150
rect 29908 2148 29932 2150
rect 29988 2148 30012 2150
rect 30068 2148 30092 2150
rect 30148 2148 30154 2150
rect 29846 2139 30154 2148
rect 29748 1958 29868 1986
rect 29840 800 29868 1958
rect 30208 1442 30236 2790
rect 30380 2576 30432 2582
rect 30380 2518 30432 2524
rect 30116 1414 30236 1442
rect 30116 800 30144 1414
rect 30392 800 30420 2518
rect 30484 1970 30512 3295
rect 31220 3194 31248 3538
rect 31208 3188 31260 3194
rect 31208 3130 31260 3136
rect 31404 3126 31432 3878
rect 32770 3839 32826 3848
rect 31576 3528 31628 3534
rect 31576 3470 31628 3476
rect 32588 3528 32640 3534
rect 32588 3470 32640 3476
rect 31588 3194 31616 3470
rect 31576 3188 31628 3194
rect 31576 3130 31628 3136
rect 32312 3188 32364 3194
rect 32312 3130 32364 3136
rect 31392 3120 31444 3126
rect 31392 3062 31444 3068
rect 31760 2984 31812 2990
rect 31760 2926 31812 2932
rect 31484 2916 31536 2922
rect 31484 2858 31536 2864
rect 30656 2508 30708 2514
rect 30656 2450 30708 2456
rect 30472 1964 30524 1970
rect 30472 1906 30524 1912
rect 30668 800 30696 2450
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 31208 2440 31260 2446
rect 31208 2382 31260 2388
rect 30944 800 30972 2382
rect 31220 800 31248 2382
rect 31496 800 31524 2858
rect 31772 800 31800 2926
rect 32036 2576 32088 2582
rect 32036 2518 32088 2524
rect 32048 800 32076 2518
rect 32324 800 32352 3130
rect 32600 800 32628 3470
rect 32784 3058 32812 3839
rect 33140 3528 33192 3534
rect 33140 3470 33192 3476
rect 32772 3052 32824 3058
rect 32772 2994 32824 3000
rect 32956 2440 33008 2446
rect 32956 2382 33008 2388
rect 32968 1306 32996 2382
rect 32876 1278 32996 1306
rect 32876 800 32904 1278
rect 33152 800 33180 3470
rect 33520 3058 33548 4100
rect 34440 3641 34468 4490
rect 35164 3936 35216 3942
rect 35164 3878 35216 3884
rect 35176 3670 35204 3878
rect 35452 3738 35480 4519
rect 35768 4542 36032 4548
rect 35716 4490 35768 4496
rect 35808 4480 35860 4486
rect 35808 4422 35860 4428
rect 35820 4214 35848 4422
rect 35808 4208 35860 4214
rect 35808 4150 35860 4156
rect 35900 4072 35952 4078
rect 35900 4014 35952 4020
rect 35624 4004 35676 4010
rect 35624 3946 35676 3952
rect 35440 3732 35492 3738
rect 35440 3674 35492 3680
rect 35164 3664 35216 3670
rect 34426 3632 34482 3641
rect 35164 3606 35216 3612
rect 34426 3567 34482 3576
rect 35348 3596 35400 3602
rect 35348 3538 35400 3544
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 33968 3528 34020 3534
rect 33968 3470 34020 3476
rect 33508 3052 33560 3058
rect 33508 2994 33560 3000
rect 33612 2774 33640 3470
rect 33784 3460 33836 3466
rect 33784 3402 33836 3408
rect 33520 2746 33640 2774
rect 33796 2774 33824 3402
rect 33876 3392 33928 3398
rect 33876 3334 33928 3340
rect 33888 3126 33916 3334
rect 33876 3120 33928 3126
rect 33876 3062 33928 3068
rect 33796 2746 33916 2774
rect 33520 1578 33548 2746
rect 33888 2650 33916 2746
rect 33876 2644 33928 2650
rect 33876 2586 33928 2592
rect 33692 2576 33744 2582
rect 33692 2518 33744 2524
rect 33428 1550 33548 1578
rect 33428 800 33456 1550
rect 33704 800 33732 2518
rect 33888 2310 33916 2586
rect 33876 2304 33928 2310
rect 33876 2246 33928 2252
rect 33980 800 34008 3470
rect 34060 3392 34112 3398
rect 34058 3360 34060 3369
rect 34112 3360 34114 3369
rect 34058 3295 34114 3304
rect 34796 3188 34848 3194
rect 34796 3130 34848 3136
rect 35256 3188 35308 3194
rect 35256 3130 35308 3136
rect 34520 2984 34572 2990
rect 34520 2926 34572 2932
rect 34612 2984 34664 2990
rect 34612 2926 34664 2932
rect 34244 2848 34296 2854
rect 34244 2790 34296 2796
rect 34256 800 34284 2790
rect 34532 2650 34560 2926
rect 34520 2644 34572 2650
rect 34520 2586 34572 2592
rect 34624 1442 34652 2926
rect 34808 2650 34836 3130
rect 35164 3052 35216 3058
rect 34900 3012 35164 3040
rect 34796 2644 34848 2650
rect 34796 2586 34848 2592
rect 34900 1442 34928 3012
rect 35164 2994 35216 3000
rect 35268 2774 35296 3130
rect 35360 2854 35388 3538
rect 35348 2848 35400 2854
rect 35348 2790 35400 2796
rect 35176 2746 35296 2774
rect 35176 1578 35204 2746
rect 35440 2372 35492 2378
rect 35440 2314 35492 2320
rect 34532 1414 34652 1442
rect 34808 1414 34928 1442
rect 35084 1550 35204 1578
rect 34532 800 34560 1414
rect 34808 800 34836 1414
rect 35084 800 35112 1550
rect 35452 1170 35480 2314
rect 35360 1142 35480 1170
rect 35360 800 35388 1142
rect 35636 800 35664 3946
rect 35912 3913 35940 4014
rect 36004 3942 36032 4542
rect 37462 4448 37518 4457
rect 37462 4383 37518 4392
rect 37476 4010 37504 4383
rect 37556 4140 37608 4146
rect 37556 4082 37608 4088
rect 37464 4004 37516 4010
rect 37464 3946 37516 3952
rect 35992 3936 36044 3942
rect 35898 3904 35954 3913
rect 35992 3878 36044 3884
rect 36360 3936 36412 3942
rect 36360 3878 36412 3884
rect 35898 3839 35954 3848
rect 35990 3632 36046 3641
rect 35990 3567 35992 3576
rect 36044 3567 36046 3576
rect 35992 3538 36044 3544
rect 36176 3528 36228 3534
rect 36082 3496 36138 3505
rect 36176 3470 36228 3476
rect 36082 3431 36138 3440
rect 36096 3398 36124 3431
rect 36084 3392 36136 3398
rect 36084 3334 36136 3340
rect 35900 1420 35952 1426
rect 35900 1362 35952 1368
rect 35912 800 35940 1362
rect 36188 800 36216 3470
rect 36268 3392 36320 3398
rect 36268 3334 36320 3340
rect 36280 2514 36308 3334
rect 36372 3097 36400 3878
rect 37070 3836 37378 3845
rect 37070 3834 37076 3836
rect 37132 3834 37156 3836
rect 37212 3834 37236 3836
rect 37292 3834 37316 3836
rect 37372 3834 37378 3836
rect 37132 3782 37134 3834
rect 37314 3782 37316 3834
rect 37070 3780 37076 3782
rect 37132 3780 37156 3782
rect 37212 3780 37236 3782
rect 37292 3780 37316 3782
rect 37372 3780 37378 3782
rect 37070 3771 37378 3780
rect 36912 3596 36964 3602
rect 36912 3538 36964 3544
rect 36452 3460 36504 3466
rect 36452 3402 36504 3408
rect 36358 3088 36414 3097
rect 36358 3023 36414 3032
rect 36464 2922 36492 3402
rect 36820 2984 36872 2990
rect 36820 2926 36872 2932
rect 36452 2916 36504 2922
rect 36452 2858 36504 2864
rect 36544 2916 36596 2922
rect 36544 2858 36596 2864
rect 36268 2508 36320 2514
rect 36268 2450 36320 2456
rect 36556 1442 36584 2858
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 36464 1414 36584 1442
rect 36464 800 36492 1414
rect 36740 800 36768 2790
rect 36832 2650 36860 2926
rect 36820 2644 36872 2650
rect 36820 2586 36872 2592
rect 36924 1850 36952 3538
rect 37070 2748 37378 2757
rect 37070 2746 37076 2748
rect 37132 2746 37156 2748
rect 37212 2746 37236 2748
rect 37292 2746 37316 2748
rect 37372 2746 37378 2748
rect 37132 2694 37134 2746
rect 37314 2694 37316 2746
rect 37070 2692 37076 2694
rect 37132 2692 37156 2694
rect 37212 2692 37236 2694
rect 37292 2692 37316 2694
rect 37372 2692 37378 2694
rect 37070 2683 37378 2692
rect 37372 2508 37424 2514
rect 37292 2468 37372 2496
rect 37004 2304 37056 2310
rect 37004 2246 37056 2252
rect 37096 2304 37148 2310
rect 37096 2246 37148 2252
rect 37016 2106 37044 2246
rect 37004 2100 37056 2106
rect 37004 2042 37056 2048
rect 36924 1822 37044 1850
rect 37016 800 37044 1822
rect 37108 1426 37136 2246
rect 37096 1420 37148 1426
rect 37096 1362 37148 1368
rect 37292 800 37320 2468
rect 37372 2450 37424 2456
rect 37568 800 37596 4082
rect 37740 3936 37792 3942
rect 37740 3878 37792 3884
rect 37752 3641 37780 3878
rect 37738 3632 37794 3641
rect 37738 3567 37794 3576
rect 38212 3466 38240 4966
rect 38396 4622 38424 6190
rect 40040 6180 40092 6186
rect 40040 6122 40092 6128
rect 39764 6112 39816 6118
rect 39764 6054 39816 6060
rect 38660 5228 38712 5234
rect 38660 5170 38712 5176
rect 38752 5228 38804 5234
rect 38752 5170 38804 5176
rect 39488 5228 39540 5234
rect 39488 5170 39540 5176
rect 38672 4758 38700 5170
rect 38764 4826 38792 5170
rect 39212 5024 39264 5030
rect 39212 4966 39264 4972
rect 38752 4820 38804 4826
rect 38752 4762 38804 4768
rect 38660 4752 38712 4758
rect 38660 4694 38712 4700
rect 38764 4690 38792 4762
rect 39224 4758 39252 4966
rect 39500 4826 39528 5170
rect 39776 5030 39804 6054
rect 40052 5642 40080 6122
rect 42996 5914 43024 6190
rect 45560 6112 45612 6118
rect 45560 6054 45612 6060
rect 46940 6112 46992 6118
rect 46940 6054 46992 6060
rect 41696 5908 41748 5914
rect 41696 5850 41748 5856
rect 42984 5908 43036 5914
rect 42984 5850 43036 5856
rect 40132 5772 40184 5778
rect 40132 5714 40184 5720
rect 39856 5636 39908 5642
rect 39856 5578 39908 5584
rect 40040 5636 40092 5642
rect 40040 5578 40092 5584
rect 39868 5545 39896 5578
rect 39854 5536 39910 5545
rect 39854 5471 39910 5480
rect 40144 5234 40172 5714
rect 40500 5636 40552 5642
rect 40500 5578 40552 5584
rect 40512 5234 40540 5578
rect 40682 5536 40738 5545
rect 40682 5471 40738 5480
rect 40132 5228 40184 5234
rect 40132 5170 40184 5176
rect 40500 5228 40552 5234
rect 40500 5170 40552 5176
rect 39764 5024 39816 5030
rect 40144 5001 40172 5170
rect 40696 5166 40724 5471
rect 41708 5370 41736 5850
rect 42800 5704 42852 5710
rect 42800 5646 42852 5652
rect 41696 5364 41748 5370
rect 41696 5306 41748 5312
rect 42616 5364 42668 5370
rect 42616 5306 42668 5312
rect 41052 5228 41104 5234
rect 41052 5170 41104 5176
rect 41236 5228 41288 5234
rect 41236 5170 41288 5176
rect 40684 5160 40736 5166
rect 40222 5128 40278 5137
rect 40684 5102 40736 5108
rect 40222 5063 40224 5072
rect 40276 5063 40278 5072
rect 40224 5034 40276 5040
rect 39764 4966 39816 4972
rect 40130 4992 40186 5001
rect 39488 4820 39540 4826
rect 39488 4762 39540 4768
rect 39120 4752 39172 4758
rect 38934 4720 38990 4729
rect 38752 4684 38804 4690
rect 39120 4694 39172 4700
rect 39212 4752 39264 4758
rect 39212 4694 39264 4700
rect 38934 4655 38990 4664
rect 38752 4626 38804 4632
rect 38384 4616 38436 4622
rect 38384 4558 38436 4564
rect 38948 4486 38976 4655
rect 38936 4480 38988 4486
rect 38934 4448 38936 4457
rect 38988 4448 38990 4457
rect 38934 4383 38990 4392
rect 39132 4146 39160 4694
rect 39776 4282 39804 4966
rect 40130 4927 40186 4936
rect 41064 4690 41092 5170
rect 41248 4826 41276 5170
rect 41236 4820 41288 4826
rect 41236 4762 41288 4768
rect 41052 4684 41104 4690
rect 41052 4626 41104 4632
rect 41708 4672 41736 5306
rect 42432 5296 42484 5302
rect 42628 5273 42656 5306
rect 42614 5264 42670 5273
rect 42432 5238 42484 5244
rect 42444 5030 42472 5238
rect 42536 5222 42614 5250
rect 42432 5024 42484 5030
rect 42432 4966 42484 4972
rect 42432 4820 42484 4826
rect 42536 4808 42564 5222
rect 42614 5199 42670 5208
rect 42812 5166 42840 5646
rect 42800 5160 42852 5166
rect 42800 5102 42852 5108
rect 42484 4780 42564 4808
rect 42432 4762 42484 4768
rect 42892 4752 42944 4758
rect 42892 4694 42944 4700
rect 41788 4684 41840 4690
rect 41708 4644 41788 4672
rect 40592 4480 40644 4486
rect 40592 4422 40644 4428
rect 39764 4276 39816 4282
rect 39764 4218 39816 4224
rect 39120 4140 39172 4146
rect 39120 4082 39172 4088
rect 40132 4072 40184 4078
rect 40132 4014 40184 4020
rect 39764 3936 39816 3942
rect 39764 3878 39816 3884
rect 38658 3768 38714 3777
rect 38658 3703 38714 3712
rect 38842 3768 38898 3777
rect 38842 3703 38898 3712
rect 39212 3732 39264 3738
rect 38672 3602 38700 3703
rect 38660 3596 38712 3602
rect 38660 3538 38712 3544
rect 38752 3528 38804 3534
rect 38752 3470 38804 3476
rect 38200 3460 38252 3466
rect 38200 3402 38252 3408
rect 38108 2984 38160 2990
rect 38108 2926 38160 2932
rect 38016 2644 38068 2650
rect 38016 2586 38068 2592
rect 37832 2576 37884 2582
rect 37832 2518 37884 2524
rect 37844 800 37872 2518
rect 38028 2446 38056 2586
rect 38016 2440 38068 2446
rect 38016 2382 38068 2388
rect 38120 800 38148 2926
rect 38660 2916 38712 2922
rect 38660 2858 38712 2864
rect 38384 1420 38436 1426
rect 38384 1362 38436 1368
rect 38396 800 38424 1362
rect 38672 800 38700 2858
rect 38764 1873 38792 3470
rect 38856 3466 38884 3703
rect 39212 3674 39264 3680
rect 38844 3460 38896 3466
rect 38844 3402 38896 3408
rect 38856 2650 38884 3402
rect 38936 3188 38988 3194
rect 38936 3130 38988 3136
rect 38844 2644 38896 2650
rect 38844 2586 38896 2592
rect 38750 1864 38806 1873
rect 38750 1799 38806 1808
rect 38948 800 38976 3130
rect 39224 800 39252 3674
rect 39776 3505 39804 3878
rect 40144 3738 40172 4014
rect 40604 3913 40632 4422
rect 41708 4146 41736 4644
rect 41788 4626 41840 4632
rect 41696 4140 41748 4146
rect 41696 4082 41748 4088
rect 40590 3904 40646 3913
rect 40590 3839 40646 3848
rect 40132 3732 40184 3738
rect 40132 3674 40184 3680
rect 40224 3732 40276 3738
rect 40224 3674 40276 3680
rect 39948 3528 40000 3534
rect 39762 3496 39818 3505
rect 39762 3431 39818 3440
rect 39868 3488 39948 3516
rect 39488 3392 39540 3398
rect 39488 3334 39540 3340
rect 39500 800 39528 3334
rect 39868 3194 39896 3488
rect 39948 3470 40000 3476
rect 40236 3398 40264 3674
rect 40224 3392 40276 3398
rect 40224 3334 40276 3340
rect 39856 3188 39908 3194
rect 39856 3130 39908 3136
rect 40604 3126 40632 3839
rect 42248 3732 42300 3738
rect 42248 3674 42300 3680
rect 41604 3596 41656 3602
rect 41604 3538 41656 3544
rect 41616 3126 41644 3538
rect 41788 3392 41840 3398
rect 41788 3334 41840 3340
rect 41696 3188 41748 3194
rect 41696 3130 41748 3136
rect 40592 3120 40644 3126
rect 40592 3062 40644 3068
rect 41604 3120 41656 3126
rect 41604 3062 41656 3068
rect 40132 3052 40184 3058
rect 40132 2994 40184 3000
rect 39948 2440 40000 2446
rect 39948 2382 40000 2388
rect 39764 2372 39816 2378
rect 39764 2314 39816 2320
rect 39776 800 39804 2314
rect 39960 1426 39988 2382
rect 40144 2310 40172 2994
rect 40592 2984 40644 2990
rect 40592 2926 40644 2932
rect 40316 2644 40368 2650
rect 40316 2586 40368 2592
rect 40132 2304 40184 2310
rect 40132 2246 40184 2252
rect 40144 2106 40172 2246
rect 40132 2100 40184 2106
rect 40132 2042 40184 2048
rect 40040 1760 40092 1766
rect 40040 1702 40092 1708
rect 39948 1420 40000 1426
rect 39948 1362 40000 1368
rect 40052 800 40080 1702
rect 40328 800 40356 2586
rect 40604 800 40632 2926
rect 41236 2916 41288 2922
rect 41156 2876 41236 2904
rect 40868 2508 40920 2514
rect 40868 2450 40920 2456
rect 40880 800 40908 2450
rect 41156 800 41184 2876
rect 41236 2858 41288 2864
rect 41420 2100 41472 2106
rect 41420 2042 41472 2048
rect 41432 800 41460 2042
rect 41616 1970 41644 3062
rect 41604 1964 41656 1970
rect 41604 1906 41656 1912
rect 41708 800 41736 3130
rect 41800 1902 41828 3334
rect 41972 2304 42024 2310
rect 41972 2246 42024 2252
rect 41788 1896 41840 1902
rect 41788 1838 41840 1844
rect 41984 800 42012 2246
rect 42260 800 42288 3674
rect 42904 3618 42932 4694
rect 42996 4146 43024 5850
rect 45572 5710 45600 6054
rect 45560 5704 45612 5710
rect 43442 5672 43498 5681
rect 45560 5646 45612 5652
rect 43442 5607 43498 5616
rect 43076 5568 43128 5574
rect 43076 5510 43128 5516
rect 42984 4140 43036 4146
rect 42984 4082 43036 4088
rect 43088 4026 43116 5510
rect 43456 5234 43484 5607
rect 45192 5568 45244 5574
rect 45192 5510 45244 5516
rect 44294 5468 44602 5477
rect 44294 5466 44300 5468
rect 44356 5466 44380 5468
rect 44436 5466 44460 5468
rect 44516 5466 44540 5468
rect 44596 5466 44602 5468
rect 44356 5414 44358 5466
rect 44538 5414 44540 5466
rect 44294 5412 44300 5414
rect 44356 5412 44380 5414
rect 44436 5412 44460 5414
rect 44516 5412 44540 5414
rect 44596 5412 44602 5414
rect 44294 5403 44602 5412
rect 44362 5264 44418 5273
rect 43444 5228 43496 5234
rect 44730 5264 44786 5273
rect 44362 5199 44418 5208
rect 44548 5228 44600 5234
rect 43444 5170 43496 5176
rect 43444 5024 43496 5030
rect 43444 4966 43496 4972
rect 43456 4826 43484 4966
rect 44376 4826 44404 5199
rect 45204 5234 45232 5510
rect 44730 5199 44732 5208
rect 44548 5170 44600 5176
rect 44784 5199 44786 5208
rect 45192 5228 45244 5234
rect 44732 5170 44784 5176
rect 45192 5170 45244 5176
rect 44560 5098 44588 5170
rect 44548 5092 44600 5098
rect 44548 5034 44600 5040
rect 44640 5024 44692 5030
rect 44744 5001 44772 5170
rect 45204 5080 45232 5170
rect 45376 5092 45428 5098
rect 45204 5052 45376 5080
rect 45376 5034 45428 5040
rect 44640 4966 44692 4972
rect 44730 4992 44786 5001
rect 43444 4820 43496 4826
rect 43444 4762 43496 4768
rect 44364 4820 44416 4826
rect 44364 4762 44416 4768
rect 44376 4622 44404 4762
rect 44652 4622 44680 4966
rect 44730 4927 44786 4936
rect 43352 4616 43404 4622
rect 43352 4558 43404 4564
rect 44364 4616 44416 4622
rect 44364 4558 44416 4564
rect 44640 4616 44692 4622
rect 44640 4558 44692 4564
rect 45192 4616 45244 4622
rect 45192 4558 45244 4564
rect 42812 3590 42932 3618
rect 42996 3998 43116 4026
rect 42432 3528 42484 3534
rect 42432 3470 42484 3476
rect 42616 3528 42668 3534
rect 42812 3516 42840 3590
rect 42668 3488 42840 3516
rect 42892 3528 42944 3534
rect 42616 3470 42668 3476
rect 42996 3516 43024 3998
rect 43076 3936 43128 3942
rect 43074 3904 43076 3913
rect 43128 3904 43130 3913
rect 43074 3839 43130 3848
rect 42944 3488 43024 3516
rect 42892 3470 42944 3476
rect 42444 2854 42472 3470
rect 42524 3188 42576 3194
rect 42524 3130 42576 3136
rect 42432 2848 42484 2854
rect 42432 2790 42484 2796
rect 42536 800 42564 3130
rect 42904 3097 42932 3470
rect 43088 3182 43300 3210
rect 43088 3126 43116 3182
rect 43076 3120 43128 3126
rect 42890 3088 42946 3097
rect 43076 3062 43128 3068
rect 43168 3120 43220 3126
rect 43168 3062 43220 3068
rect 42890 3023 42946 3032
rect 43076 2916 43128 2922
rect 43076 2858 43128 2864
rect 42800 2848 42852 2854
rect 42800 2790 42852 2796
rect 42812 800 42840 2790
rect 43088 1766 43116 2858
rect 43076 1760 43128 1766
rect 43076 1702 43128 1708
rect 43180 1578 43208 3062
rect 43272 2854 43300 3182
rect 43260 2848 43312 2854
rect 43260 2790 43312 2796
rect 43088 1550 43208 1578
rect 43088 800 43116 1550
rect 43364 800 43392 4558
rect 44294 4380 44602 4389
rect 44294 4378 44300 4380
rect 44356 4378 44380 4380
rect 44436 4378 44460 4380
rect 44516 4378 44540 4380
rect 44596 4378 44602 4380
rect 44356 4326 44358 4378
rect 44538 4326 44540 4378
rect 44294 4324 44300 4326
rect 44356 4324 44380 4326
rect 44436 4324 44460 4326
rect 44516 4324 44540 4326
rect 44596 4324 44602 4326
rect 44294 4315 44602 4324
rect 44652 4282 44680 4558
rect 44640 4276 44692 4282
rect 44640 4218 44692 4224
rect 45204 4078 45232 4558
rect 45572 4486 45600 5646
rect 46952 5574 46980 6054
rect 46020 5568 46072 5574
rect 46020 5510 46072 5516
rect 46940 5568 46992 5574
rect 46940 5510 46992 5516
rect 46032 4690 46060 5510
rect 46388 5228 46440 5234
rect 46388 5170 46440 5176
rect 46296 5024 46348 5030
rect 46296 4966 46348 4972
rect 46308 4690 46336 4966
rect 46400 4690 46428 5170
rect 46756 5024 46808 5030
rect 46756 4966 46808 4972
rect 46020 4684 46072 4690
rect 46020 4626 46072 4632
rect 46296 4684 46348 4690
rect 46296 4626 46348 4632
rect 46388 4684 46440 4690
rect 46388 4626 46440 4632
rect 45560 4480 45612 4486
rect 45560 4422 45612 4428
rect 45744 4140 45796 4146
rect 45744 4082 45796 4088
rect 45192 4072 45244 4078
rect 44086 4040 44142 4049
rect 44270 4040 44326 4049
rect 44086 3975 44142 3984
rect 44180 4004 44232 4010
rect 43628 3936 43680 3942
rect 43628 3878 43680 3884
rect 43640 800 43668 3878
rect 44100 3505 44128 3975
rect 45192 4014 45244 4020
rect 44270 3975 44326 3984
rect 44180 3946 44232 3952
rect 44086 3496 44142 3505
rect 44086 3431 44142 3440
rect 43904 3052 43956 3058
rect 43904 2994 43956 3000
rect 43916 800 43944 2994
rect 44192 800 44220 3946
rect 44284 3670 44312 3975
rect 45756 3738 45784 4082
rect 45928 3936 45980 3942
rect 45928 3878 45980 3884
rect 46664 3936 46716 3942
rect 46664 3878 46716 3884
rect 45744 3732 45796 3738
rect 45744 3674 45796 3680
rect 44272 3664 44324 3670
rect 44272 3606 44324 3612
rect 44638 3632 44694 3641
rect 45940 3602 45968 3878
rect 44638 3567 44640 3576
rect 44692 3567 44694 3576
rect 45192 3596 45244 3602
rect 44640 3538 44692 3544
rect 45192 3538 45244 3544
rect 45928 3596 45980 3602
rect 45928 3538 45980 3544
rect 44294 3292 44602 3301
rect 44294 3290 44300 3292
rect 44356 3290 44380 3292
rect 44436 3290 44460 3292
rect 44516 3290 44540 3292
rect 44596 3290 44602 3292
rect 44356 3238 44358 3290
rect 44538 3238 44540 3290
rect 44294 3236 44300 3238
rect 44356 3236 44380 3238
rect 44436 3236 44460 3238
rect 44516 3236 44540 3238
rect 44596 3236 44602 3238
rect 44294 3227 44602 3236
rect 44272 2916 44324 2922
rect 44272 2858 44324 2864
rect 44284 2650 44312 2858
rect 44652 2666 44680 3538
rect 45204 3505 45232 3538
rect 46676 3534 46704 3878
rect 45376 3528 45428 3534
rect 45190 3496 45246 3505
rect 45376 3470 45428 3476
rect 46572 3528 46624 3534
rect 46572 3470 46624 3476
rect 46664 3528 46716 3534
rect 46664 3470 46716 3476
rect 45190 3431 45246 3440
rect 45008 3188 45060 3194
rect 45008 3130 45060 3136
rect 45020 3040 45048 3130
rect 45192 3052 45244 3058
rect 45020 3012 45192 3040
rect 45192 2994 45244 3000
rect 45284 2916 45336 2922
rect 45284 2858 45336 2864
rect 45296 2666 45324 2858
rect 44272 2644 44324 2650
rect 44272 2586 44324 2592
rect 44560 2638 44680 2666
rect 45020 2638 45324 2666
rect 44560 2514 44588 2638
rect 44548 2508 44600 2514
rect 44548 2450 44600 2456
rect 44640 2508 44692 2514
rect 44640 2450 44692 2456
rect 44294 2204 44602 2213
rect 44294 2202 44300 2204
rect 44356 2202 44380 2204
rect 44436 2202 44460 2204
rect 44516 2202 44540 2204
rect 44596 2202 44602 2204
rect 44356 2150 44358 2202
rect 44538 2150 44540 2202
rect 44294 2148 44300 2150
rect 44356 2148 44380 2150
rect 44436 2148 44460 2150
rect 44516 2148 44540 2150
rect 44596 2148 44602 2150
rect 44294 2139 44602 2148
rect 44652 1306 44680 2450
rect 44824 2304 44876 2310
rect 44824 2246 44876 2252
rect 44732 1760 44784 1766
rect 44732 1702 44784 1708
rect 44468 1278 44680 1306
rect 44468 800 44496 1278
rect 44744 800 44772 1702
rect 44836 1698 44864 2246
rect 44824 1692 44876 1698
rect 44824 1634 44876 1640
rect 45020 800 45048 2638
rect 45192 2576 45244 2582
rect 45192 2518 45244 2524
rect 45204 2106 45232 2518
rect 45284 2372 45336 2378
rect 45284 2314 45336 2320
rect 45192 2100 45244 2106
rect 45192 2042 45244 2048
rect 45296 800 45324 2314
rect 45388 2038 45416 3470
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 45480 2310 45508 3334
rect 46112 3188 46164 3194
rect 46112 3130 46164 3136
rect 45560 2984 45612 2990
rect 45560 2926 45612 2932
rect 45468 2304 45520 2310
rect 45468 2246 45520 2252
rect 45376 2032 45428 2038
rect 45376 1974 45428 1980
rect 45572 800 45600 2926
rect 45836 2576 45888 2582
rect 45836 2518 45888 2524
rect 45848 800 45876 2518
rect 46124 800 46152 3130
rect 46584 3058 46612 3470
rect 46572 3052 46624 3058
rect 46572 2994 46624 3000
rect 46584 2961 46612 2994
rect 46570 2952 46626 2961
rect 46570 2887 46626 2896
rect 46768 2530 46796 4966
rect 46952 3398 46980 5510
rect 47044 4078 47072 6666
rect 48148 5846 48176 6666
rect 52184 6656 52236 6662
rect 52184 6598 52236 6604
rect 50896 6180 50948 6186
rect 50896 6122 50948 6128
rect 49792 5908 49844 5914
rect 49792 5850 49844 5856
rect 48136 5840 48188 5846
rect 48136 5782 48188 5788
rect 49700 5636 49752 5642
rect 49700 5578 49752 5584
rect 48320 5296 48372 5302
rect 47122 5264 47178 5273
rect 48320 5238 48372 5244
rect 47122 5199 47178 5208
rect 47136 5098 47164 5199
rect 47124 5092 47176 5098
rect 47124 5034 47176 5040
rect 48332 4826 48360 5238
rect 49332 5160 49384 5166
rect 49160 5120 49332 5148
rect 48320 4820 48372 4826
rect 48320 4762 48372 4768
rect 48596 4752 48648 4758
rect 48594 4720 48596 4729
rect 48648 4720 48650 4729
rect 48594 4655 48650 4664
rect 49056 4208 49108 4214
rect 49056 4150 49108 4156
rect 47032 4072 47084 4078
rect 49068 4049 49096 4150
rect 47032 4014 47084 4020
rect 49054 4040 49110 4049
rect 47044 3738 47072 4014
rect 49054 3975 49110 3984
rect 47584 3936 47636 3942
rect 47584 3878 47636 3884
rect 47768 3936 47820 3942
rect 47768 3878 47820 3884
rect 47596 3777 47624 3878
rect 47582 3768 47638 3777
rect 47032 3732 47084 3738
rect 47582 3703 47638 3712
rect 47032 3674 47084 3680
rect 47030 3632 47086 3641
rect 47030 3567 47086 3576
rect 47044 3466 47072 3567
rect 47032 3460 47084 3466
rect 47032 3402 47084 3408
rect 46940 3392 46992 3398
rect 46938 3360 46940 3369
rect 46992 3360 46994 3369
rect 46938 3295 46994 3304
rect 47044 3126 47072 3402
rect 47124 3392 47176 3398
rect 47124 3334 47176 3340
rect 47584 3392 47636 3398
rect 47584 3334 47636 3340
rect 47032 3120 47084 3126
rect 47032 3062 47084 3068
rect 46676 2502 46796 2530
rect 46388 2100 46440 2106
rect 46388 2042 46440 2048
rect 46400 800 46428 2042
rect 46676 800 46704 2502
rect 46848 2440 46900 2446
rect 47136 2417 47164 3334
rect 47216 3052 47268 3058
rect 47216 2994 47268 3000
rect 46848 2382 46900 2388
rect 47122 2408 47178 2417
rect 46860 1766 46888 2382
rect 47122 2343 47178 2352
rect 46940 2032 46992 2038
rect 46940 1974 46992 1980
rect 46848 1760 46900 1766
rect 46848 1702 46900 1708
rect 46952 800 46980 1974
rect 47136 1834 47164 2343
rect 47124 1828 47176 1834
rect 47124 1770 47176 1776
rect 47228 800 47256 2994
rect 47596 2310 47624 3334
rect 47676 2848 47728 2854
rect 47676 2790 47728 2796
rect 47584 2304 47636 2310
rect 47584 2246 47636 2252
rect 47688 1442 47716 2790
rect 47504 1414 47716 1442
rect 47504 800 47532 1414
rect 47780 800 47808 3878
rect 48044 3732 48096 3738
rect 48044 3674 48096 3680
rect 48056 800 48084 3674
rect 48872 3392 48924 3398
rect 48872 3334 48924 3340
rect 48596 2916 48648 2922
rect 48596 2858 48648 2864
rect 48320 1420 48372 1426
rect 48320 1362 48372 1368
rect 48332 800 48360 1362
rect 48608 800 48636 2858
rect 48884 800 48912 3334
rect 49160 800 49188 5120
rect 49332 5102 49384 5108
rect 49608 5024 49660 5030
rect 49608 4966 49660 4972
rect 49620 4758 49648 4966
rect 49608 4752 49660 4758
rect 49608 4694 49660 4700
rect 49608 4616 49660 4622
rect 49608 4558 49660 4564
rect 49620 4282 49648 4558
rect 49608 4276 49660 4282
rect 49608 4218 49660 4224
rect 49712 4146 49740 5578
rect 49804 5574 49832 5850
rect 50252 5704 50304 5710
rect 50252 5646 50304 5652
rect 50528 5704 50580 5710
rect 50528 5646 50580 5652
rect 49792 5568 49844 5574
rect 49792 5510 49844 5516
rect 49804 4146 49832 5510
rect 50160 5092 50212 5098
rect 50160 5034 50212 5040
rect 50172 4622 50200 5034
rect 50160 4616 50212 4622
rect 50160 4558 50212 4564
rect 49884 4548 49936 4554
rect 49884 4490 49936 4496
rect 49332 4140 49384 4146
rect 49332 4082 49384 4088
rect 49700 4140 49752 4146
rect 49700 4082 49752 4088
rect 49792 4140 49844 4146
rect 49792 4082 49844 4088
rect 49344 3602 49372 4082
rect 49608 4072 49660 4078
rect 49608 4014 49660 4020
rect 49332 3596 49384 3602
rect 49332 3538 49384 3544
rect 49344 3466 49372 3538
rect 49424 3528 49476 3534
rect 49424 3470 49476 3476
rect 49332 3460 49384 3466
rect 49332 3402 49384 3408
rect 49344 2774 49372 3402
rect 49436 3194 49464 3470
rect 49620 3194 49648 4014
rect 49896 4010 49924 4490
rect 49884 4004 49936 4010
rect 49884 3946 49936 3952
rect 49976 4004 50028 4010
rect 49976 3946 50028 3952
rect 49424 3188 49476 3194
rect 49424 3130 49476 3136
rect 49608 3188 49660 3194
rect 49608 3130 49660 3136
rect 49884 3120 49936 3126
rect 49884 3062 49936 3068
rect 49896 2854 49924 3062
rect 49884 2848 49936 2854
rect 49884 2790 49936 2796
rect 49344 2746 49556 2774
rect 49528 2650 49556 2746
rect 49516 2644 49568 2650
rect 49516 2586 49568 2592
rect 49608 2644 49660 2650
rect 49608 2586 49660 2592
rect 49424 1964 49476 1970
rect 49424 1906 49476 1912
rect 49436 800 49464 1906
rect 49620 1426 49648 2586
rect 49700 2508 49752 2514
rect 49700 2450 49752 2456
rect 49608 1420 49660 1426
rect 49608 1362 49660 1368
rect 49712 800 49740 2450
rect 49988 800 50016 3946
rect 50160 3664 50212 3670
rect 50160 3606 50212 3612
rect 50066 3360 50122 3369
rect 50066 3295 50122 3304
rect 50080 3126 50108 3295
rect 50068 3120 50120 3126
rect 50068 3062 50120 3068
rect 50172 2553 50200 3606
rect 50158 2544 50214 2553
rect 50158 2479 50214 2488
rect 50264 800 50292 5646
rect 50436 2848 50488 2854
rect 50436 2790 50488 2796
rect 50448 2582 50476 2790
rect 50436 2576 50488 2582
rect 50436 2518 50488 2524
rect 50540 800 50568 5646
rect 50908 5234 50936 6122
rect 51356 6112 51408 6118
rect 51356 6054 51408 6060
rect 52000 6112 52052 6118
rect 52000 6054 52052 6060
rect 51172 5296 51224 5302
rect 51172 5238 51224 5244
rect 50896 5228 50948 5234
rect 50896 5170 50948 5176
rect 51184 4826 51212 5238
rect 51264 5160 51316 5166
rect 51264 5102 51316 5108
rect 51172 4820 51224 4826
rect 51172 4762 51224 4768
rect 50896 4480 50948 4486
rect 50896 4422 50948 4428
rect 50908 3534 50936 4422
rect 51276 3913 51304 5102
rect 51368 4146 51396 6054
rect 51518 6012 51826 6021
rect 51518 6010 51524 6012
rect 51580 6010 51604 6012
rect 51660 6010 51684 6012
rect 51740 6010 51764 6012
rect 51820 6010 51826 6012
rect 51580 5958 51582 6010
rect 51762 5958 51764 6010
rect 51518 5956 51524 5958
rect 51580 5956 51604 5958
rect 51660 5956 51684 5958
rect 51740 5956 51764 5958
rect 51820 5956 51826 5958
rect 51518 5947 51826 5956
rect 51448 5704 51500 5710
rect 51448 5646 51500 5652
rect 51908 5704 51960 5710
rect 51908 5646 51960 5652
rect 51356 4140 51408 4146
rect 51356 4082 51408 4088
rect 51262 3904 51318 3913
rect 51262 3839 51318 3848
rect 51172 3664 51224 3670
rect 51092 3624 51172 3652
rect 50712 3528 50764 3534
rect 50712 3470 50764 3476
rect 50896 3528 50948 3534
rect 50896 3470 50948 3476
rect 50724 3126 50752 3470
rect 50712 3120 50764 3126
rect 50712 3062 50764 3068
rect 50804 3052 50856 3058
rect 50856 3012 51028 3040
rect 50804 2994 50856 3000
rect 51000 2922 51028 3012
rect 50988 2916 51040 2922
rect 50988 2858 51040 2864
rect 50804 2304 50856 2310
rect 50804 2246 50856 2252
rect 50816 800 50844 2246
rect 51092 800 51120 3624
rect 51172 3606 51224 3612
rect 51172 3528 51224 3534
rect 51368 3516 51396 4082
rect 51224 3488 51396 3516
rect 51172 3470 51224 3476
rect 51184 3097 51212 3470
rect 51170 3088 51226 3097
rect 51170 3023 51226 3032
rect 51356 3052 51408 3058
rect 51184 2310 51212 3023
rect 51356 2994 51408 3000
rect 51172 2304 51224 2310
rect 51172 2246 51224 2252
rect 51368 800 51396 2994
rect 51460 2564 51488 5646
rect 51518 4924 51826 4933
rect 51518 4922 51524 4924
rect 51580 4922 51604 4924
rect 51660 4922 51684 4924
rect 51740 4922 51764 4924
rect 51820 4922 51826 4924
rect 51580 4870 51582 4922
rect 51762 4870 51764 4922
rect 51518 4868 51524 4870
rect 51580 4868 51604 4870
rect 51660 4868 51684 4870
rect 51740 4868 51764 4870
rect 51820 4868 51826 4870
rect 51518 4859 51826 4868
rect 51518 3836 51826 3845
rect 51518 3834 51524 3836
rect 51580 3834 51604 3836
rect 51660 3834 51684 3836
rect 51740 3834 51764 3836
rect 51820 3834 51826 3836
rect 51580 3782 51582 3834
rect 51762 3782 51764 3834
rect 51518 3780 51524 3782
rect 51580 3780 51604 3782
rect 51660 3780 51684 3782
rect 51740 3780 51764 3782
rect 51820 3780 51826 3782
rect 51518 3771 51826 3780
rect 51518 2748 51826 2757
rect 51518 2746 51524 2748
rect 51580 2746 51604 2748
rect 51660 2746 51684 2748
rect 51740 2746 51764 2748
rect 51820 2746 51826 2748
rect 51580 2694 51582 2746
rect 51762 2694 51764 2746
rect 51518 2692 51524 2694
rect 51580 2692 51604 2694
rect 51660 2692 51684 2694
rect 51740 2692 51764 2694
rect 51820 2692 51826 2694
rect 51518 2683 51826 2692
rect 51460 2536 51672 2564
rect 51448 2440 51500 2446
rect 51448 2382 51500 2388
rect 51460 2106 51488 2382
rect 51448 2100 51500 2106
rect 51448 2042 51500 2048
rect 51644 800 51672 2536
rect 51920 800 51948 5646
rect 52012 5234 52040 6054
rect 52196 5914 52224 6598
rect 52184 5908 52236 5914
rect 52184 5850 52236 5856
rect 52000 5228 52052 5234
rect 52000 5170 52052 5176
rect 52090 4584 52146 4593
rect 52090 4519 52146 4528
rect 52104 4486 52132 4519
rect 52092 4480 52144 4486
rect 52092 4422 52144 4428
rect 52196 4146 52224 5850
rect 52276 5772 52328 5778
rect 52276 5714 52328 5720
rect 52184 4140 52236 4146
rect 52184 4082 52236 4088
rect 52196 3602 52224 4082
rect 52184 3596 52236 3602
rect 52184 3538 52236 3544
rect 52288 2904 52316 5714
rect 54760 5636 54812 5642
rect 54760 5578 54812 5584
rect 54024 5364 54076 5370
rect 54024 5306 54076 5312
rect 52552 5092 52604 5098
rect 52552 5034 52604 5040
rect 52736 5092 52788 5098
rect 52736 5034 52788 5040
rect 52460 4820 52512 4826
rect 52460 4762 52512 4768
rect 52472 4282 52500 4762
rect 52460 4276 52512 4282
rect 52460 4218 52512 4224
rect 52564 3602 52592 5034
rect 52644 5024 52696 5030
rect 52644 4966 52696 4972
rect 52656 4282 52684 4966
rect 52644 4276 52696 4282
rect 52644 4218 52696 4224
rect 52552 3596 52604 3602
rect 52552 3538 52604 3544
rect 52644 3596 52696 3602
rect 52644 3538 52696 3544
rect 52656 3194 52684 3538
rect 52644 3188 52696 3194
rect 52644 3130 52696 3136
rect 52460 3120 52512 3126
rect 52460 3062 52512 3068
rect 52196 2876 52316 2904
rect 52368 2916 52420 2922
rect 52196 800 52224 2876
rect 52368 2858 52420 2864
rect 52380 800 52408 2858
rect 52472 800 52500 3062
rect 52748 2564 52776 5034
rect 52828 5024 52880 5030
rect 52828 4966 52880 4972
rect 53012 5024 53064 5030
rect 53012 4966 53064 4972
rect 52840 3466 52868 4966
rect 53024 4214 53052 4966
rect 53748 4684 53800 4690
rect 53748 4626 53800 4632
rect 53656 4276 53708 4282
rect 53656 4218 53708 4224
rect 53012 4208 53064 4214
rect 53012 4150 53064 4156
rect 53668 4078 53696 4218
rect 53760 4078 53788 4626
rect 54036 4622 54064 5306
rect 54024 4616 54076 4622
rect 54024 4558 54076 4564
rect 54772 4486 54800 5578
rect 55220 5568 55272 5574
rect 55220 5510 55272 5516
rect 54760 4480 54812 4486
rect 54760 4422 54812 4428
rect 54772 4282 54800 4422
rect 54760 4276 54812 4282
rect 54760 4218 54812 4224
rect 53656 4072 53708 4078
rect 53656 4014 53708 4020
rect 53748 4072 53800 4078
rect 53748 4014 53800 4020
rect 54484 3936 54536 3942
rect 54484 3878 54536 3884
rect 54496 3641 54524 3878
rect 54482 3632 54538 3641
rect 54482 3567 54538 3576
rect 52828 3460 52880 3466
rect 52828 3402 52880 3408
rect 54024 3392 54076 3398
rect 54024 3334 54076 3340
rect 52564 2536 52776 2564
rect 52564 800 52592 2536
rect 52736 2440 52788 2446
rect 52736 2382 52788 2388
rect 52748 2038 52776 2382
rect 52736 2032 52788 2038
rect 52736 1974 52788 1980
rect 54036 1766 54064 3334
rect 54208 2848 54260 2854
rect 54208 2790 54260 2796
rect 54220 1902 54248 2790
rect 54772 2446 54800 4218
rect 55232 4010 55260 5510
rect 55404 5296 55456 5302
rect 55404 5238 55456 5244
rect 55312 5024 55364 5030
rect 55312 4966 55364 4972
rect 55324 4146 55352 4966
rect 55312 4140 55364 4146
rect 55312 4082 55364 4088
rect 55220 4004 55272 4010
rect 55220 3946 55272 3952
rect 55232 3738 55260 3946
rect 55312 3936 55364 3942
rect 55312 3878 55364 3884
rect 55220 3732 55272 3738
rect 55220 3674 55272 3680
rect 55324 3398 55352 3878
rect 55416 3602 55444 5238
rect 55680 5228 55732 5234
rect 55680 5170 55732 5176
rect 55588 5160 55640 5166
rect 55494 5128 55550 5137
rect 55588 5102 55640 5108
rect 55494 5063 55550 5072
rect 55508 4622 55536 5063
rect 55496 4616 55548 4622
rect 55496 4558 55548 4564
rect 55496 3664 55548 3670
rect 55496 3606 55548 3612
rect 55404 3596 55456 3602
rect 55404 3538 55456 3544
rect 55312 3392 55364 3398
rect 55312 3334 55364 3340
rect 55508 2990 55536 3606
rect 55496 2984 55548 2990
rect 55496 2926 55548 2932
rect 55600 2854 55628 5102
rect 55692 4826 55720 5170
rect 55772 5024 55824 5030
rect 55772 4966 55824 4972
rect 55680 4820 55732 4826
rect 55680 4762 55732 4768
rect 55784 4026 55812 4966
rect 56600 4480 56652 4486
rect 56600 4422 56652 4428
rect 57244 4480 57296 4486
rect 57244 4422 57296 4428
rect 55784 3998 55904 4026
rect 55680 3936 55732 3942
rect 55680 3878 55732 3884
rect 55692 3398 55720 3878
rect 55876 3602 55904 3998
rect 56324 3936 56376 3942
rect 56324 3878 56376 3884
rect 56048 3732 56100 3738
rect 56048 3674 56100 3680
rect 55864 3596 55916 3602
rect 55864 3538 55916 3544
rect 55876 3505 55904 3538
rect 55862 3496 55918 3505
rect 55862 3431 55918 3440
rect 55680 3392 55732 3398
rect 55680 3334 55732 3340
rect 55772 3392 55824 3398
rect 55772 3334 55824 3340
rect 55956 3392 56008 3398
rect 55956 3334 56008 3340
rect 55784 2854 55812 3334
rect 55864 3120 55916 3126
rect 55864 3062 55916 3068
rect 55588 2848 55640 2854
rect 55588 2790 55640 2796
rect 55772 2848 55824 2854
rect 55772 2790 55824 2796
rect 54760 2440 54812 2446
rect 54760 2382 54812 2388
rect 54208 1896 54260 1902
rect 54208 1838 54260 1844
rect 55784 1834 55812 2790
rect 55876 2582 55904 3062
rect 55968 3058 55996 3334
rect 56060 3126 56088 3674
rect 56232 3596 56284 3602
rect 56232 3538 56284 3544
rect 56048 3120 56100 3126
rect 56048 3062 56100 3068
rect 55956 3052 56008 3058
rect 55956 2994 56008 3000
rect 56244 2990 56272 3538
rect 56336 3058 56364 3878
rect 56324 3052 56376 3058
rect 56324 2994 56376 3000
rect 56232 2984 56284 2990
rect 56232 2926 56284 2932
rect 56612 2854 56640 4422
rect 57256 4146 57284 4422
rect 56692 4140 56744 4146
rect 56692 4082 56744 4088
rect 57244 4140 57296 4146
rect 57244 4082 57296 4088
rect 56600 2848 56652 2854
rect 56600 2790 56652 2796
rect 55864 2576 55916 2582
rect 55864 2518 55916 2524
rect 56704 2514 56732 4082
rect 57428 3528 57480 3534
rect 57428 3470 57480 3476
rect 57440 2650 57468 3470
rect 57428 2644 57480 2650
rect 57428 2586 57480 2592
rect 56692 2508 56744 2514
rect 56692 2450 56744 2456
rect 56232 2440 56284 2446
rect 56232 2382 56284 2388
rect 56244 1970 56272 2382
rect 56232 1964 56284 1970
rect 56232 1906 56284 1912
rect 55772 1828 55824 1834
rect 55772 1770 55824 1776
rect 54024 1760 54076 1766
rect 54024 1702 54076 1708
rect 7286 0 7342 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7654 0 7710 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 7930 0 7986 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8206 0 8262 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8574 0 8630 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8850 0 8906 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9126 0 9182 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9494 0 9550 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9770 0 9826 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10046 0 10102 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10414 0 10470 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10690 0 10746 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 10966 0 11022 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11334 0 11390 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11610 0 11666 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11886 0 11942 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12254 0 12310 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12530 0 12586 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12806 0 12862 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13082 0 13138 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13450 0 13506 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13726 0 13782 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14002 0 14058 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14370 0 14426 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14646 0 14702 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 14922 0 14978 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15290 0 15346 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15566 0 15622 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15842 0 15898 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16210 0 16266 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16486 0 16542 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16762 0 16818 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17130 0 17186 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17406 0 17462 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17682 0 17738 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18050 0 18106 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18326 0 18382 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18602 0 18658 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 18970 0 19026 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19246 0 19302 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19522 0 19578 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19890 0 19946 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20166 0 20222 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20442 0 20498 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20810 0 20866 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21086 0 21142 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21362 0 21418 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21730 0 21786 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22006 0 22062 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22282 0 22338 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22650 0 22706 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 22926 0 22982 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23202 0 23258 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23570 0 23626 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23846 0 23902 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24122 0 24178 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24490 0 24546 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24766 0 24822 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25042 0 25098 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25410 0 25466 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25686 0 25742 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 25962 0 26018 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26238 0 26294 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26606 0 26662 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26882 0 26938 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27158 0 27214 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27526 0 27582 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27802 0 27858 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28078 0 28134 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28446 0 28502 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28722 0 28778 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 28998 0 29054 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29366 0 29422 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29642 0 29698 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 29918 0 29974 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30286 0 30342 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30562 0 30618 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30838 0 30894 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31206 0 31262 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31482 0 31538 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31758 0 31814 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32126 0 32182 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32402 0 32458 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32678 0 32734 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33046 0 33102 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33322 0 33378 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33598 0 33654 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 33966 0 34022 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34242 0 34298 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34518 0 34574 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34886 0 34942 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35162 0 35218 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35438 0 35494 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35806 0 35862 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36082 0 36138 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36358 0 36414 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36726 0 36782 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37002 0 37058 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37278 0 37334 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37646 0 37702 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 37922 0 37978 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38198 0 38254 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38566 0 38622 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38842 0 38898 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39118 0 39174 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39394 0 39450 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39762 0 39818 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40038 0 40094 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40314 0 40370 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40682 0 40738 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 40958 0 41014 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41234 0 41290 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41602 0 41658 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41878 0 41934 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42154 0 42210 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42522 0 42578 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42798 0 42854 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43074 0 43130 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43442 0 43498 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43718 0 43774 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 43994 0 44050 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44362 0 44418 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44638 0 44694 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 44914 0 44970 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45282 0 45338 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45558 0 45614 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45834 0 45890 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46202 0 46258 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46478 0 46534 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46754 0 46810 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47122 0 47178 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47398 0 47454 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47674 0 47730 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48042 0 48098 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48318 0 48374 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48594 0 48650 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 48962 0 49018 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49238 0 49294 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49514 0 49570 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49882 0 49938 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50158 0 50214 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50434 0 50490 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50802 0 50858 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51078 0 51134 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51354 0 51410 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51722 0 51778 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 51998 0 52054 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52274 0 52330 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52550 0 52606 800
<< via2 >>
rect 8180 7098 8236 7100
rect 8260 7098 8316 7100
rect 8340 7098 8396 7100
rect 8420 7098 8476 7100
rect 8180 7046 8226 7098
rect 8226 7046 8236 7098
rect 8260 7046 8290 7098
rect 8290 7046 8302 7098
rect 8302 7046 8316 7098
rect 8340 7046 8354 7098
rect 8354 7046 8366 7098
rect 8366 7046 8396 7098
rect 8420 7046 8430 7098
rect 8430 7046 8476 7098
rect 8180 7044 8236 7046
rect 8260 7044 8316 7046
rect 8340 7044 8396 7046
rect 8420 7044 8476 7046
rect 15404 7642 15460 7644
rect 15484 7642 15540 7644
rect 15564 7642 15620 7644
rect 15644 7642 15700 7644
rect 15404 7590 15450 7642
rect 15450 7590 15460 7642
rect 15484 7590 15514 7642
rect 15514 7590 15526 7642
rect 15526 7590 15540 7642
rect 15564 7590 15578 7642
rect 15578 7590 15590 7642
rect 15590 7590 15620 7642
rect 15644 7590 15654 7642
rect 15654 7590 15700 7642
rect 15404 7588 15460 7590
rect 15484 7588 15540 7590
rect 15564 7588 15620 7590
rect 15644 7588 15700 7590
rect 22628 7098 22684 7100
rect 22708 7098 22764 7100
rect 22788 7098 22844 7100
rect 22868 7098 22924 7100
rect 22628 7046 22674 7098
rect 22674 7046 22684 7098
rect 22708 7046 22738 7098
rect 22738 7046 22750 7098
rect 22750 7046 22764 7098
rect 22788 7046 22802 7098
rect 22802 7046 22814 7098
rect 22814 7046 22844 7098
rect 22868 7046 22878 7098
rect 22878 7046 22924 7098
rect 22628 7044 22684 7046
rect 22708 7044 22764 7046
rect 22788 7044 22844 7046
rect 22868 7044 22924 7046
rect 29852 7642 29908 7644
rect 29932 7642 29988 7644
rect 30012 7642 30068 7644
rect 30092 7642 30148 7644
rect 29852 7590 29898 7642
rect 29898 7590 29908 7642
rect 29932 7590 29962 7642
rect 29962 7590 29974 7642
rect 29974 7590 29988 7642
rect 30012 7590 30026 7642
rect 30026 7590 30038 7642
rect 30038 7590 30068 7642
rect 30092 7590 30102 7642
rect 30102 7590 30148 7642
rect 29852 7588 29908 7590
rect 29932 7588 29988 7590
rect 30012 7588 30068 7590
rect 30092 7588 30148 7590
rect 37076 7098 37132 7100
rect 37156 7098 37212 7100
rect 37236 7098 37292 7100
rect 37316 7098 37372 7100
rect 37076 7046 37122 7098
rect 37122 7046 37132 7098
rect 37156 7046 37186 7098
rect 37186 7046 37198 7098
rect 37198 7046 37212 7098
rect 37236 7046 37250 7098
rect 37250 7046 37262 7098
rect 37262 7046 37292 7098
rect 37316 7046 37326 7098
rect 37326 7046 37372 7098
rect 37076 7044 37132 7046
rect 37156 7044 37212 7046
rect 37236 7044 37292 7046
rect 37316 7044 37372 7046
rect 44300 7642 44356 7644
rect 44380 7642 44436 7644
rect 44460 7642 44516 7644
rect 44540 7642 44596 7644
rect 44300 7590 44346 7642
rect 44346 7590 44356 7642
rect 44380 7590 44410 7642
rect 44410 7590 44422 7642
rect 44422 7590 44436 7642
rect 44460 7590 44474 7642
rect 44474 7590 44486 7642
rect 44486 7590 44516 7642
rect 44540 7590 44550 7642
rect 44550 7590 44596 7642
rect 44300 7588 44356 7590
rect 44380 7588 44436 7590
rect 44460 7588 44516 7590
rect 44540 7588 44596 7590
rect 51524 7098 51580 7100
rect 51604 7098 51660 7100
rect 51684 7098 51740 7100
rect 51764 7098 51820 7100
rect 51524 7046 51570 7098
rect 51570 7046 51580 7098
rect 51604 7046 51634 7098
rect 51634 7046 51646 7098
rect 51646 7046 51660 7098
rect 51684 7046 51698 7098
rect 51698 7046 51710 7098
rect 51710 7046 51740 7098
rect 51764 7046 51774 7098
rect 51774 7046 51820 7098
rect 51524 7044 51580 7046
rect 51604 7044 51660 7046
rect 51684 7044 51740 7046
rect 51764 7044 51820 7046
rect 8180 6010 8236 6012
rect 8260 6010 8316 6012
rect 8340 6010 8396 6012
rect 8420 6010 8476 6012
rect 8180 5958 8226 6010
rect 8226 5958 8236 6010
rect 8260 5958 8290 6010
rect 8290 5958 8302 6010
rect 8302 5958 8316 6010
rect 8340 5958 8354 6010
rect 8354 5958 8366 6010
rect 8366 5958 8396 6010
rect 8420 5958 8430 6010
rect 8430 5958 8476 6010
rect 8180 5956 8236 5958
rect 8260 5956 8316 5958
rect 8340 5956 8396 5958
rect 8420 5956 8476 5958
rect 3146 3340 3148 3360
rect 3148 3340 3200 3360
rect 3200 3340 3202 3360
rect 3146 3304 3202 3340
rect 5354 5072 5410 5128
rect 4434 3596 4490 3632
rect 4434 3576 4436 3596
rect 4436 3576 4488 3596
rect 4488 3576 4490 3596
rect 4066 2488 4122 2544
rect 5446 3440 5502 3496
rect 6274 4392 6330 4448
rect 6826 4256 6882 4312
rect 7654 4120 7710 4176
rect 7286 1944 7342 2000
rect 15404 6554 15460 6556
rect 15484 6554 15540 6556
rect 15564 6554 15620 6556
rect 15644 6554 15700 6556
rect 15404 6502 15450 6554
rect 15450 6502 15460 6554
rect 15484 6502 15514 6554
rect 15514 6502 15526 6554
rect 15526 6502 15540 6554
rect 15564 6502 15578 6554
rect 15578 6502 15590 6554
rect 15590 6502 15620 6554
rect 15644 6502 15654 6554
rect 15654 6502 15700 6554
rect 15404 6500 15460 6502
rect 15484 6500 15540 6502
rect 15564 6500 15620 6502
rect 15644 6500 15700 6502
rect 8180 4922 8236 4924
rect 8260 4922 8316 4924
rect 8340 4922 8396 4924
rect 8420 4922 8476 4924
rect 8180 4870 8226 4922
rect 8226 4870 8236 4922
rect 8260 4870 8290 4922
rect 8290 4870 8302 4922
rect 8302 4870 8316 4922
rect 8340 4870 8354 4922
rect 8354 4870 8366 4922
rect 8366 4870 8396 4922
rect 8420 4870 8430 4922
rect 8430 4870 8476 4922
rect 8180 4868 8236 4870
rect 8260 4868 8316 4870
rect 8340 4868 8396 4870
rect 8420 4868 8476 4870
rect 8298 4528 8354 4584
rect 8180 3834 8236 3836
rect 8260 3834 8316 3836
rect 8340 3834 8396 3836
rect 8420 3834 8476 3836
rect 8180 3782 8226 3834
rect 8226 3782 8236 3834
rect 8260 3782 8290 3834
rect 8290 3782 8302 3834
rect 8302 3782 8316 3834
rect 8340 3782 8354 3834
rect 8354 3782 8366 3834
rect 8366 3782 8396 3834
rect 8420 3782 8430 3834
rect 8430 3782 8476 3834
rect 8180 3780 8236 3782
rect 8260 3780 8316 3782
rect 8340 3780 8396 3782
rect 8420 3780 8476 3782
rect 8180 2746 8236 2748
rect 8260 2746 8316 2748
rect 8340 2746 8396 2748
rect 8420 2746 8476 2748
rect 8180 2694 8226 2746
rect 8226 2694 8236 2746
rect 8260 2694 8290 2746
rect 8290 2694 8302 2746
rect 8302 2694 8316 2746
rect 8340 2694 8354 2746
rect 8354 2694 8366 2746
rect 8366 2694 8396 2746
rect 8420 2694 8430 2746
rect 8430 2694 8476 2746
rect 8180 2692 8236 2694
rect 8260 2692 8316 2694
rect 8340 2692 8396 2694
rect 8420 2692 8476 2694
rect 8758 3168 8814 3224
rect 8758 3052 8814 3088
rect 8758 3032 8760 3052
rect 8760 3032 8812 3052
rect 8812 3032 8814 3052
rect 9678 4664 9734 4720
rect 9402 1672 9458 1728
rect 9678 3304 9734 3360
rect 10782 2796 10784 2816
rect 10784 2796 10836 2816
rect 10836 2796 10838 2816
rect 10782 2760 10838 2796
rect 11058 5072 11114 5128
rect 12162 3848 12218 3904
rect 12346 3596 12402 3632
rect 12346 3576 12348 3596
rect 12348 3576 12400 3596
rect 12400 3576 12402 3596
rect 12162 1808 12218 1864
rect 12622 4664 12678 4720
rect 13450 5244 13452 5264
rect 13452 5244 13504 5264
rect 13504 5244 13506 5264
rect 13450 5208 13506 5244
rect 12990 4392 13046 4448
rect 13082 3712 13138 3768
rect 13358 3440 13414 3496
rect 14002 4120 14058 4176
rect 13266 3168 13322 3224
rect 13910 3596 13966 3632
rect 13910 3576 13912 3596
rect 13912 3576 13964 3596
rect 13964 3576 13966 3596
rect 15404 5466 15460 5468
rect 15484 5466 15540 5468
rect 15564 5466 15620 5468
rect 15644 5466 15700 5468
rect 15404 5414 15450 5466
rect 15450 5414 15460 5466
rect 15484 5414 15514 5466
rect 15514 5414 15526 5466
rect 15526 5414 15540 5466
rect 15564 5414 15578 5466
rect 15578 5414 15590 5466
rect 15590 5414 15620 5466
rect 15644 5414 15654 5466
rect 15654 5414 15700 5466
rect 15404 5412 15460 5414
rect 15484 5412 15540 5414
rect 15564 5412 15620 5414
rect 15644 5412 15700 5414
rect 15404 4378 15460 4380
rect 15484 4378 15540 4380
rect 15564 4378 15620 4380
rect 15644 4378 15700 4380
rect 15404 4326 15450 4378
rect 15450 4326 15460 4378
rect 15484 4326 15514 4378
rect 15514 4326 15526 4378
rect 15526 4326 15540 4378
rect 15564 4326 15578 4378
rect 15578 4326 15590 4378
rect 15590 4326 15620 4378
rect 15644 4326 15654 4378
rect 15654 4326 15700 4378
rect 15404 4324 15460 4326
rect 15484 4324 15540 4326
rect 15564 4324 15620 4326
rect 15644 4324 15700 4326
rect 15658 4120 15714 4176
rect 15404 3290 15460 3292
rect 15484 3290 15540 3292
rect 15564 3290 15620 3292
rect 15644 3290 15700 3292
rect 15404 3238 15450 3290
rect 15450 3238 15460 3290
rect 15484 3238 15514 3290
rect 15514 3238 15526 3290
rect 15526 3238 15540 3290
rect 15564 3238 15578 3290
rect 15578 3238 15590 3290
rect 15590 3238 15620 3290
rect 15644 3238 15654 3290
rect 15654 3238 15700 3290
rect 15404 3236 15460 3238
rect 15484 3236 15540 3238
rect 15564 3236 15620 3238
rect 15644 3236 15700 3238
rect 15290 2760 15346 2816
rect 15404 2202 15460 2204
rect 15484 2202 15540 2204
rect 15564 2202 15620 2204
rect 15644 2202 15700 2204
rect 15404 2150 15450 2202
rect 15450 2150 15460 2202
rect 15484 2150 15514 2202
rect 15514 2150 15526 2202
rect 15526 2150 15540 2202
rect 15564 2150 15578 2202
rect 15578 2150 15590 2202
rect 15590 2150 15620 2202
rect 15644 2150 15654 2202
rect 15654 2150 15700 2202
rect 15404 2148 15460 2150
rect 15484 2148 15540 2150
rect 15564 2148 15620 2150
rect 15644 2148 15700 2150
rect 22628 6010 22684 6012
rect 22708 6010 22764 6012
rect 22788 6010 22844 6012
rect 22868 6010 22924 6012
rect 22628 5958 22674 6010
rect 22674 5958 22684 6010
rect 22708 5958 22738 6010
rect 22738 5958 22750 6010
rect 22750 5958 22764 6010
rect 22788 5958 22802 6010
rect 22802 5958 22814 6010
rect 22814 5958 22844 6010
rect 22868 5958 22878 6010
rect 22878 5958 22924 6010
rect 22628 5956 22684 5958
rect 22708 5956 22764 5958
rect 22788 5956 22844 5958
rect 22868 5956 22924 5958
rect 17590 4564 17592 4584
rect 17592 4564 17644 4584
rect 17644 4564 17646 4584
rect 17590 4528 17646 4564
rect 18142 4664 18198 4720
rect 17866 3984 17922 4040
rect 19062 4120 19118 4176
rect 19338 3848 19394 3904
rect 18602 2896 18658 2952
rect 19706 3440 19762 3496
rect 19798 3032 19854 3088
rect 20718 4020 20720 4040
rect 20720 4020 20772 4040
rect 20772 4020 20774 4040
rect 20718 3984 20774 4020
rect 19982 3032 20038 3088
rect 21730 3168 21786 3224
rect 21730 2896 21786 2952
rect 23018 4972 23020 4992
rect 23020 4972 23072 4992
rect 23072 4972 23074 4992
rect 23018 4936 23074 4972
rect 22628 4922 22684 4924
rect 22708 4922 22764 4924
rect 22788 4922 22844 4924
rect 22868 4922 22924 4924
rect 22628 4870 22674 4922
rect 22674 4870 22684 4922
rect 22708 4870 22738 4922
rect 22738 4870 22750 4922
rect 22750 4870 22764 4922
rect 22788 4870 22802 4922
rect 22802 4870 22814 4922
rect 22814 4870 22844 4922
rect 22868 4870 22878 4922
rect 22878 4870 22924 4922
rect 22628 4868 22684 4870
rect 22708 4868 22764 4870
rect 22788 4868 22844 4870
rect 22868 4868 22924 4870
rect 22628 3834 22684 3836
rect 22708 3834 22764 3836
rect 22788 3834 22844 3836
rect 22868 3834 22924 3836
rect 22628 3782 22674 3834
rect 22674 3782 22684 3834
rect 22708 3782 22738 3834
rect 22738 3782 22750 3834
rect 22750 3782 22764 3834
rect 22788 3782 22802 3834
rect 22802 3782 22814 3834
rect 22814 3782 22844 3834
rect 22868 3782 22878 3834
rect 22878 3782 22924 3834
rect 22628 3780 22684 3782
rect 22708 3780 22764 3782
rect 22788 3780 22844 3782
rect 22868 3780 22924 3782
rect 22628 2746 22684 2748
rect 22708 2746 22764 2748
rect 22788 2746 22844 2748
rect 22868 2746 22924 2748
rect 22628 2694 22674 2746
rect 22674 2694 22684 2746
rect 22708 2694 22738 2746
rect 22738 2694 22750 2746
rect 22750 2694 22764 2746
rect 22788 2694 22802 2746
rect 22802 2694 22814 2746
rect 22814 2694 22844 2746
rect 22868 2694 22878 2746
rect 22878 2694 22924 2746
rect 22628 2692 22684 2694
rect 22708 2692 22764 2694
rect 22788 2692 22844 2694
rect 22868 2692 22924 2694
rect 23478 1944 23534 2000
rect 24950 4120 25006 4176
rect 24858 3984 24914 4040
rect 25502 4004 25558 4040
rect 25502 3984 25504 4004
rect 25504 3984 25556 4004
rect 25556 3984 25558 4004
rect 25778 3984 25834 4040
rect 26054 3476 26056 3496
rect 26056 3476 26108 3496
rect 26108 3476 26110 3496
rect 26054 3440 26110 3476
rect 26698 2896 26754 2952
rect 26882 2488 26938 2544
rect 27250 3032 27306 3088
rect 29852 6554 29908 6556
rect 29932 6554 29988 6556
rect 30012 6554 30068 6556
rect 30092 6554 30148 6556
rect 29852 6502 29898 6554
rect 29898 6502 29908 6554
rect 29932 6502 29962 6554
rect 29962 6502 29974 6554
rect 29974 6502 29988 6554
rect 30012 6502 30026 6554
rect 30026 6502 30038 6554
rect 30038 6502 30068 6554
rect 30092 6502 30102 6554
rect 30102 6502 30148 6554
rect 29852 6500 29908 6502
rect 29932 6500 29988 6502
rect 30012 6500 30068 6502
rect 30092 6500 30148 6502
rect 27250 2352 27306 2408
rect 28262 4664 28318 4720
rect 28262 3168 28318 3224
rect 28354 1672 28410 1728
rect 29852 5466 29908 5468
rect 29932 5466 29988 5468
rect 30012 5466 30068 5468
rect 30092 5466 30148 5468
rect 29852 5414 29898 5466
rect 29898 5414 29908 5466
rect 29932 5414 29962 5466
rect 29962 5414 29974 5466
rect 29974 5414 29988 5466
rect 30012 5414 30026 5466
rect 30026 5414 30038 5466
rect 30038 5414 30068 5466
rect 30092 5414 30102 5466
rect 30102 5414 30148 5466
rect 29852 5412 29908 5414
rect 29932 5412 29988 5414
rect 30012 5412 30068 5414
rect 30092 5412 30148 5414
rect 44300 6554 44356 6556
rect 44380 6554 44436 6556
rect 44460 6554 44516 6556
rect 44540 6554 44596 6556
rect 44300 6502 44346 6554
rect 44346 6502 44356 6554
rect 44380 6502 44410 6554
rect 44410 6502 44422 6554
rect 44422 6502 44436 6554
rect 44460 6502 44474 6554
rect 44474 6502 44486 6554
rect 44486 6502 44516 6554
rect 44540 6502 44550 6554
rect 44550 6502 44596 6554
rect 44300 6500 44356 6502
rect 44380 6500 44436 6502
rect 44460 6500 44516 6502
rect 44540 6500 44596 6502
rect 30378 5208 30434 5264
rect 30286 4936 30342 4992
rect 31022 5788 31024 5808
rect 31024 5788 31076 5808
rect 31076 5788 31078 5808
rect 31022 5752 31078 5788
rect 30286 4392 30342 4448
rect 29852 4378 29908 4380
rect 29932 4378 29988 4380
rect 30012 4378 30068 4380
rect 30092 4378 30148 4380
rect 29852 4326 29898 4378
rect 29898 4326 29908 4378
rect 29932 4326 29962 4378
rect 29962 4326 29974 4378
rect 29974 4326 29988 4378
rect 30012 4326 30026 4378
rect 30026 4326 30038 4378
rect 30038 4326 30068 4378
rect 30092 4326 30102 4378
rect 30102 4326 30148 4378
rect 29852 4324 29908 4326
rect 29932 4324 29988 4326
rect 30012 4324 30068 4326
rect 30092 4324 30148 4326
rect 32126 5636 32182 5672
rect 32126 5616 32128 5636
rect 32128 5616 32180 5636
rect 32180 5616 32182 5636
rect 32586 4528 32642 4584
rect 34702 5752 34758 5808
rect 33966 5480 34022 5536
rect 33874 5072 33930 5128
rect 37076 6010 37132 6012
rect 37156 6010 37212 6012
rect 37236 6010 37292 6012
rect 37316 6010 37372 6012
rect 37076 5958 37122 6010
rect 37122 5958 37132 6010
rect 37156 5958 37186 6010
rect 37186 5958 37198 6010
rect 37198 5958 37212 6010
rect 37236 5958 37250 6010
rect 37250 5958 37262 6010
rect 37262 5958 37292 6010
rect 37316 5958 37326 6010
rect 37326 5958 37372 6010
rect 37076 5956 37132 5958
rect 37156 5956 37212 5958
rect 37236 5956 37292 5958
rect 37316 5956 37372 5958
rect 36450 5480 36506 5536
rect 36726 5072 36782 5128
rect 37076 4922 37132 4924
rect 37156 4922 37212 4924
rect 37236 4922 37292 4924
rect 37316 4922 37372 4924
rect 37076 4870 37122 4922
rect 37122 4870 37132 4922
rect 37156 4870 37186 4922
rect 37186 4870 37198 4922
rect 37198 4870 37212 4922
rect 37236 4870 37250 4922
rect 37250 4870 37262 4922
rect 37262 4870 37292 4922
rect 37316 4870 37326 4922
rect 37326 4870 37372 4922
rect 37076 4868 37132 4870
rect 37156 4868 37212 4870
rect 37236 4868 37292 4870
rect 37316 4868 37372 4870
rect 37646 4664 37702 4720
rect 35438 4528 35494 4584
rect 29852 3290 29908 3292
rect 29932 3290 29988 3292
rect 30012 3290 30068 3292
rect 30092 3290 30148 3292
rect 29852 3238 29898 3290
rect 29898 3238 29908 3290
rect 29932 3238 29962 3290
rect 29962 3238 29974 3290
rect 29974 3238 29988 3290
rect 30012 3238 30026 3290
rect 30026 3238 30038 3290
rect 30038 3238 30068 3290
rect 30092 3238 30102 3290
rect 30102 3238 30148 3290
rect 29852 3236 29908 3238
rect 29932 3236 29988 3238
rect 30012 3236 30068 3238
rect 30092 3236 30148 3238
rect 30470 3340 30472 3360
rect 30472 3340 30524 3360
rect 30524 3340 30526 3360
rect 30470 3304 30526 3340
rect 29852 2202 29908 2204
rect 29932 2202 29988 2204
rect 30012 2202 30068 2204
rect 30092 2202 30148 2204
rect 29852 2150 29898 2202
rect 29898 2150 29908 2202
rect 29932 2150 29962 2202
rect 29962 2150 29974 2202
rect 29974 2150 29988 2202
rect 30012 2150 30026 2202
rect 30026 2150 30038 2202
rect 30038 2150 30068 2202
rect 30092 2150 30102 2202
rect 30102 2150 30148 2202
rect 29852 2148 29908 2150
rect 29932 2148 29988 2150
rect 30012 2148 30068 2150
rect 30092 2148 30148 2150
rect 32770 3848 32826 3904
rect 34426 3576 34482 3632
rect 34058 3340 34060 3360
rect 34060 3340 34112 3360
rect 34112 3340 34114 3360
rect 34058 3304 34114 3340
rect 37462 4392 37518 4448
rect 35898 3848 35954 3904
rect 35990 3596 36046 3632
rect 35990 3576 35992 3596
rect 35992 3576 36044 3596
rect 36044 3576 36046 3596
rect 36082 3440 36138 3496
rect 37076 3834 37132 3836
rect 37156 3834 37212 3836
rect 37236 3834 37292 3836
rect 37316 3834 37372 3836
rect 37076 3782 37122 3834
rect 37122 3782 37132 3834
rect 37156 3782 37186 3834
rect 37186 3782 37198 3834
rect 37198 3782 37212 3834
rect 37236 3782 37250 3834
rect 37250 3782 37262 3834
rect 37262 3782 37292 3834
rect 37316 3782 37326 3834
rect 37326 3782 37372 3834
rect 37076 3780 37132 3782
rect 37156 3780 37212 3782
rect 37236 3780 37292 3782
rect 37316 3780 37372 3782
rect 36358 3032 36414 3088
rect 37076 2746 37132 2748
rect 37156 2746 37212 2748
rect 37236 2746 37292 2748
rect 37316 2746 37372 2748
rect 37076 2694 37122 2746
rect 37122 2694 37132 2746
rect 37156 2694 37186 2746
rect 37186 2694 37198 2746
rect 37198 2694 37212 2746
rect 37236 2694 37250 2746
rect 37250 2694 37262 2746
rect 37262 2694 37292 2746
rect 37316 2694 37326 2746
rect 37326 2694 37372 2746
rect 37076 2692 37132 2694
rect 37156 2692 37212 2694
rect 37236 2692 37292 2694
rect 37316 2692 37372 2694
rect 37738 3576 37794 3632
rect 39854 5480 39910 5536
rect 40682 5480 40738 5536
rect 40222 5092 40278 5128
rect 40222 5072 40224 5092
rect 40224 5072 40276 5092
rect 40276 5072 40278 5092
rect 38934 4664 38990 4720
rect 38934 4428 38936 4448
rect 38936 4428 38988 4448
rect 38988 4428 38990 4448
rect 38934 4392 38990 4428
rect 40130 4936 40186 4992
rect 42614 5208 42670 5264
rect 38658 3712 38714 3768
rect 38842 3712 38898 3768
rect 38750 1808 38806 1864
rect 40590 3848 40646 3904
rect 39762 3440 39818 3496
rect 43442 5616 43498 5672
rect 44300 5466 44356 5468
rect 44380 5466 44436 5468
rect 44460 5466 44516 5468
rect 44540 5466 44596 5468
rect 44300 5414 44346 5466
rect 44346 5414 44356 5466
rect 44380 5414 44410 5466
rect 44410 5414 44422 5466
rect 44422 5414 44436 5466
rect 44460 5414 44474 5466
rect 44474 5414 44486 5466
rect 44486 5414 44516 5466
rect 44540 5414 44550 5466
rect 44550 5414 44596 5466
rect 44300 5412 44356 5414
rect 44380 5412 44436 5414
rect 44460 5412 44516 5414
rect 44540 5412 44596 5414
rect 44362 5208 44418 5264
rect 44730 5228 44786 5264
rect 44730 5208 44732 5228
rect 44732 5208 44784 5228
rect 44784 5208 44786 5228
rect 44730 4936 44786 4992
rect 43074 3884 43076 3904
rect 43076 3884 43128 3904
rect 43128 3884 43130 3904
rect 43074 3848 43130 3884
rect 42890 3032 42946 3088
rect 44300 4378 44356 4380
rect 44380 4378 44436 4380
rect 44460 4378 44516 4380
rect 44540 4378 44596 4380
rect 44300 4326 44346 4378
rect 44346 4326 44356 4378
rect 44380 4326 44410 4378
rect 44410 4326 44422 4378
rect 44422 4326 44436 4378
rect 44460 4326 44474 4378
rect 44474 4326 44486 4378
rect 44486 4326 44516 4378
rect 44540 4326 44550 4378
rect 44550 4326 44596 4378
rect 44300 4324 44356 4326
rect 44380 4324 44436 4326
rect 44460 4324 44516 4326
rect 44540 4324 44596 4326
rect 44086 3984 44142 4040
rect 44270 3984 44326 4040
rect 44086 3440 44142 3496
rect 44638 3596 44694 3632
rect 44638 3576 44640 3596
rect 44640 3576 44692 3596
rect 44692 3576 44694 3596
rect 44300 3290 44356 3292
rect 44380 3290 44436 3292
rect 44460 3290 44516 3292
rect 44540 3290 44596 3292
rect 44300 3238 44346 3290
rect 44346 3238 44356 3290
rect 44380 3238 44410 3290
rect 44410 3238 44422 3290
rect 44422 3238 44436 3290
rect 44460 3238 44474 3290
rect 44474 3238 44486 3290
rect 44486 3238 44516 3290
rect 44540 3238 44550 3290
rect 44550 3238 44596 3290
rect 44300 3236 44356 3238
rect 44380 3236 44436 3238
rect 44460 3236 44516 3238
rect 44540 3236 44596 3238
rect 45190 3440 45246 3496
rect 44300 2202 44356 2204
rect 44380 2202 44436 2204
rect 44460 2202 44516 2204
rect 44540 2202 44596 2204
rect 44300 2150 44346 2202
rect 44346 2150 44356 2202
rect 44380 2150 44410 2202
rect 44410 2150 44422 2202
rect 44422 2150 44436 2202
rect 44460 2150 44474 2202
rect 44474 2150 44486 2202
rect 44486 2150 44516 2202
rect 44540 2150 44550 2202
rect 44550 2150 44596 2202
rect 44300 2148 44356 2150
rect 44380 2148 44436 2150
rect 44460 2148 44516 2150
rect 44540 2148 44596 2150
rect 46570 2896 46626 2952
rect 47122 5208 47178 5264
rect 48594 4700 48596 4720
rect 48596 4700 48648 4720
rect 48648 4700 48650 4720
rect 48594 4664 48650 4700
rect 49054 3984 49110 4040
rect 47582 3712 47638 3768
rect 47030 3576 47086 3632
rect 46938 3340 46940 3360
rect 46940 3340 46992 3360
rect 46992 3340 46994 3360
rect 46938 3304 46994 3340
rect 47122 2352 47178 2408
rect 50066 3304 50122 3360
rect 50158 2488 50214 2544
rect 51524 6010 51580 6012
rect 51604 6010 51660 6012
rect 51684 6010 51740 6012
rect 51764 6010 51820 6012
rect 51524 5958 51570 6010
rect 51570 5958 51580 6010
rect 51604 5958 51634 6010
rect 51634 5958 51646 6010
rect 51646 5958 51660 6010
rect 51684 5958 51698 6010
rect 51698 5958 51710 6010
rect 51710 5958 51740 6010
rect 51764 5958 51774 6010
rect 51774 5958 51820 6010
rect 51524 5956 51580 5958
rect 51604 5956 51660 5958
rect 51684 5956 51740 5958
rect 51764 5956 51820 5958
rect 51262 3848 51318 3904
rect 51170 3032 51226 3088
rect 51524 4922 51580 4924
rect 51604 4922 51660 4924
rect 51684 4922 51740 4924
rect 51764 4922 51820 4924
rect 51524 4870 51570 4922
rect 51570 4870 51580 4922
rect 51604 4870 51634 4922
rect 51634 4870 51646 4922
rect 51646 4870 51660 4922
rect 51684 4870 51698 4922
rect 51698 4870 51710 4922
rect 51710 4870 51740 4922
rect 51764 4870 51774 4922
rect 51774 4870 51820 4922
rect 51524 4868 51580 4870
rect 51604 4868 51660 4870
rect 51684 4868 51740 4870
rect 51764 4868 51820 4870
rect 51524 3834 51580 3836
rect 51604 3834 51660 3836
rect 51684 3834 51740 3836
rect 51764 3834 51820 3836
rect 51524 3782 51570 3834
rect 51570 3782 51580 3834
rect 51604 3782 51634 3834
rect 51634 3782 51646 3834
rect 51646 3782 51660 3834
rect 51684 3782 51698 3834
rect 51698 3782 51710 3834
rect 51710 3782 51740 3834
rect 51764 3782 51774 3834
rect 51774 3782 51820 3834
rect 51524 3780 51580 3782
rect 51604 3780 51660 3782
rect 51684 3780 51740 3782
rect 51764 3780 51820 3782
rect 51524 2746 51580 2748
rect 51604 2746 51660 2748
rect 51684 2746 51740 2748
rect 51764 2746 51820 2748
rect 51524 2694 51570 2746
rect 51570 2694 51580 2746
rect 51604 2694 51634 2746
rect 51634 2694 51646 2746
rect 51646 2694 51660 2746
rect 51684 2694 51698 2746
rect 51698 2694 51710 2746
rect 51710 2694 51740 2746
rect 51764 2694 51774 2746
rect 51774 2694 51820 2746
rect 51524 2692 51580 2694
rect 51604 2692 51660 2694
rect 51684 2692 51740 2694
rect 51764 2692 51820 2694
rect 52090 4528 52146 4584
rect 54482 3576 54538 3632
rect 55494 5072 55550 5128
rect 55862 3440 55918 3496
<< metal3 >>
rect 15394 7648 15710 7649
rect 15394 7584 15400 7648
rect 15464 7584 15480 7648
rect 15544 7584 15560 7648
rect 15624 7584 15640 7648
rect 15704 7584 15710 7648
rect 15394 7583 15710 7584
rect 29842 7648 30158 7649
rect 29842 7584 29848 7648
rect 29912 7584 29928 7648
rect 29992 7584 30008 7648
rect 30072 7584 30088 7648
rect 30152 7584 30158 7648
rect 29842 7583 30158 7584
rect 44290 7648 44606 7649
rect 44290 7584 44296 7648
rect 44360 7584 44376 7648
rect 44440 7584 44456 7648
rect 44520 7584 44536 7648
rect 44600 7584 44606 7648
rect 44290 7583 44606 7584
rect 8170 7104 8486 7105
rect 8170 7040 8176 7104
rect 8240 7040 8256 7104
rect 8320 7040 8336 7104
rect 8400 7040 8416 7104
rect 8480 7040 8486 7104
rect 8170 7039 8486 7040
rect 22618 7104 22934 7105
rect 22618 7040 22624 7104
rect 22688 7040 22704 7104
rect 22768 7040 22784 7104
rect 22848 7040 22864 7104
rect 22928 7040 22934 7104
rect 22618 7039 22934 7040
rect 37066 7104 37382 7105
rect 37066 7040 37072 7104
rect 37136 7040 37152 7104
rect 37216 7040 37232 7104
rect 37296 7040 37312 7104
rect 37376 7040 37382 7104
rect 37066 7039 37382 7040
rect 51514 7104 51830 7105
rect 51514 7040 51520 7104
rect 51584 7040 51600 7104
rect 51664 7040 51680 7104
rect 51744 7040 51760 7104
rect 51824 7040 51830 7104
rect 51514 7039 51830 7040
rect 15394 6560 15710 6561
rect 15394 6496 15400 6560
rect 15464 6496 15480 6560
rect 15544 6496 15560 6560
rect 15624 6496 15640 6560
rect 15704 6496 15710 6560
rect 15394 6495 15710 6496
rect 29842 6560 30158 6561
rect 29842 6496 29848 6560
rect 29912 6496 29928 6560
rect 29992 6496 30008 6560
rect 30072 6496 30088 6560
rect 30152 6496 30158 6560
rect 29842 6495 30158 6496
rect 44290 6560 44606 6561
rect 44290 6496 44296 6560
rect 44360 6496 44376 6560
rect 44440 6496 44456 6560
rect 44520 6496 44536 6560
rect 44600 6496 44606 6560
rect 44290 6495 44606 6496
rect 8170 6016 8486 6017
rect 8170 5952 8176 6016
rect 8240 5952 8256 6016
rect 8320 5952 8336 6016
rect 8400 5952 8416 6016
rect 8480 5952 8486 6016
rect 8170 5951 8486 5952
rect 22618 6016 22934 6017
rect 22618 5952 22624 6016
rect 22688 5952 22704 6016
rect 22768 5952 22784 6016
rect 22848 5952 22864 6016
rect 22928 5952 22934 6016
rect 22618 5951 22934 5952
rect 37066 6016 37382 6017
rect 37066 5952 37072 6016
rect 37136 5952 37152 6016
rect 37216 5952 37232 6016
rect 37296 5952 37312 6016
rect 37376 5952 37382 6016
rect 37066 5951 37382 5952
rect 51514 6016 51830 6017
rect 51514 5952 51520 6016
rect 51584 5952 51600 6016
rect 51664 5952 51680 6016
rect 51744 5952 51760 6016
rect 51824 5952 51830 6016
rect 51514 5951 51830 5952
rect 31017 5810 31083 5813
rect 34697 5810 34763 5813
rect 31017 5808 34763 5810
rect 31017 5752 31022 5808
rect 31078 5752 34702 5808
rect 34758 5752 34763 5808
rect 31017 5750 34763 5752
rect 31017 5747 31083 5750
rect 34697 5747 34763 5750
rect 32121 5674 32187 5677
rect 43437 5674 43503 5677
rect 32121 5672 43503 5674
rect 32121 5616 32126 5672
rect 32182 5616 43442 5672
rect 43498 5616 43503 5672
rect 32121 5614 43503 5616
rect 32121 5611 32187 5614
rect 43437 5611 43503 5614
rect 33961 5538 34027 5541
rect 36445 5538 36511 5541
rect 33961 5536 36511 5538
rect 33961 5480 33966 5536
rect 34022 5480 36450 5536
rect 36506 5480 36511 5536
rect 33961 5478 36511 5480
rect 33961 5475 34027 5478
rect 36445 5475 36511 5478
rect 39849 5538 39915 5541
rect 40677 5538 40743 5541
rect 39849 5536 40743 5538
rect 39849 5480 39854 5536
rect 39910 5480 40682 5536
rect 40738 5480 40743 5536
rect 39849 5478 40743 5480
rect 39849 5475 39915 5478
rect 40677 5475 40743 5478
rect 15394 5472 15710 5473
rect 15394 5408 15400 5472
rect 15464 5408 15480 5472
rect 15544 5408 15560 5472
rect 15624 5408 15640 5472
rect 15704 5408 15710 5472
rect 15394 5407 15710 5408
rect 29842 5472 30158 5473
rect 29842 5408 29848 5472
rect 29912 5408 29928 5472
rect 29992 5408 30008 5472
rect 30072 5408 30088 5472
rect 30152 5408 30158 5472
rect 29842 5407 30158 5408
rect 44290 5472 44606 5473
rect 44290 5408 44296 5472
rect 44360 5408 44376 5472
rect 44440 5408 44456 5472
rect 44520 5408 44536 5472
rect 44600 5408 44606 5472
rect 44290 5407 44606 5408
rect 13445 5266 13511 5269
rect 30373 5266 30439 5269
rect 13445 5264 30439 5266
rect 13445 5208 13450 5264
rect 13506 5208 30378 5264
rect 30434 5208 30439 5264
rect 13445 5206 30439 5208
rect 13445 5203 13511 5206
rect 30373 5203 30439 5206
rect 42609 5266 42675 5269
rect 44357 5266 44423 5269
rect 42609 5264 44423 5266
rect 42609 5208 42614 5264
rect 42670 5208 44362 5264
rect 44418 5208 44423 5264
rect 42609 5206 44423 5208
rect 42609 5203 42675 5206
rect 44357 5203 44423 5206
rect 44725 5266 44791 5269
rect 47117 5266 47183 5269
rect 44725 5264 47183 5266
rect 44725 5208 44730 5264
rect 44786 5208 47122 5264
rect 47178 5208 47183 5264
rect 44725 5206 47183 5208
rect 44725 5203 44791 5206
rect 47117 5203 47183 5206
rect 5349 5130 5415 5133
rect 11053 5130 11119 5133
rect 5349 5128 11119 5130
rect 5349 5072 5354 5128
rect 5410 5072 11058 5128
rect 11114 5072 11119 5128
rect 5349 5070 11119 5072
rect 5349 5067 5415 5070
rect 11053 5067 11119 5070
rect 33869 5130 33935 5133
rect 36721 5130 36787 5133
rect 40217 5130 40283 5133
rect 55489 5130 55555 5133
rect 33869 5128 55555 5130
rect 33869 5072 33874 5128
rect 33930 5072 36726 5128
rect 36782 5072 40222 5128
rect 40278 5072 55494 5128
rect 55550 5072 55555 5128
rect 33869 5070 55555 5072
rect 33869 5067 33935 5070
rect 36721 5067 36787 5070
rect 40217 5067 40283 5070
rect 55489 5067 55555 5070
rect 23013 4994 23079 4997
rect 30281 4994 30347 4997
rect 23013 4992 30347 4994
rect 23013 4936 23018 4992
rect 23074 4936 30286 4992
rect 30342 4936 30347 4992
rect 23013 4934 30347 4936
rect 23013 4931 23079 4934
rect 30281 4931 30347 4934
rect 40125 4994 40191 4997
rect 44725 4994 44791 4997
rect 40125 4992 44791 4994
rect 40125 4936 40130 4992
rect 40186 4936 44730 4992
rect 44786 4936 44791 4992
rect 40125 4934 44791 4936
rect 40125 4931 40191 4934
rect 44725 4931 44791 4934
rect 8170 4928 8486 4929
rect 8170 4864 8176 4928
rect 8240 4864 8256 4928
rect 8320 4864 8336 4928
rect 8400 4864 8416 4928
rect 8480 4864 8486 4928
rect 8170 4863 8486 4864
rect 22618 4928 22934 4929
rect 22618 4864 22624 4928
rect 22688 4864 22704 4928
rect 22768 4864 22784 4928
rect 22848 4864 22864 4928
rect 22928 4864 22934 4928
rect 22618 4863 22934 4864
rect 37066 4928 37382 4929
rect 37066 4864 37072 4928
rect 37136 4864 37152 4928
rect 37216 4864 37232 4928
rect 37296 4864 37312 4928
rect 37376 4864 37382 4928
rect 37066 4863 37382 4864
rect 51514 4928 51830 4929
rect 51514 4864 51520 4928
rect 51584 4864 51600 4928
rect 51664 4864 51680 4928
rect 51744 4864 51760 4928
rect 51824 4864 51830 4928
rect 51514 4863 51830 4864
rect 9673 4722 9739 4725
rect 12617 4722 12683 4725
rect 9673 4720 12683 4722
rect 9673 4664 9678 4720
rect 9734 4664 12622 4720
rect 12678 4664 12683 4720
rect 9673 4662 12683 4664
rect 9673 4659 9739 4662
rect 12617 4659 12683 4662
rect 12934 4660 12940 4724
rect 13004 4722 13010 4724
rect 18137 4722 18203 4725
rect 13004 4720 18203 4722
rect 13004 4664 18142 4720
rect 18198 4664 18203 4720
rect 13004 4662 18203 4664
rect 13004 4660 13010 4662
rect 18137 4659 18203 4662
rect 28257 4722 28323 4725
rect 37641 4722 37707 4725
rect 28257 4720 37707 4722
rect 28257 4664 28262 4720
rect 28318 4664 37646 4720
rect 37702 4664 37707 4720
rect 28257 4662 37707 4664
rect 28257 4659 28323 4662
rect 37641 4659 37707 4662
rect 38929 4722 38995 4725
rect 48589 4722 48655 4725
rect 38929 4720 48655 4722
rect 38929 4664 38934 4720
rect 38990 4664 48594 4720
rect 48650 4664 48655 4720
rect 38929 4662 48655 4664
rect 38929 4659 38995 4662
rect 48589 4659 48655 4662
rect 8293 4586 8359 4589
rect 17585 4586 17651 4589
rect 8293 4584 17651 4586
rect 8293 4528 8298 4584
rect 8354 4528 17590 4584
rect 17646 4528 17651 4584
rect 8293 4526 17651 4528
rect 8293 4523 8359 4526
rect 17585 4523 17651 4526
rect 32581 4586 32647 4589
rect 35433 4586 35499 4589
rect 52085 4586 52151 4589
rect 32581 4584 52151 4586
rect 32581 4528 32586 4584
rect 32642 4528 35438 4584
rect 35494 4528 52090 4584
rect 52146 4528 52151 4584
rect 32581 4526 52151 4528
rect 32581 4523 32647 4526
rect 35433 4523 35499 4526
rect 52085 4523 52151 4526
rect 6269 4450 6335 4453
rect 12985 4450 13051 4453
rect 6269 4448 13051 4450
rect 6269 4392 6274 4448
rect 6330 4392 12990 4448
rect 13046 4392 13051 4448
rect 6269 4390 13051 4392
rect 6269 4387 6335 4390
rect 12985 4387 13051 4390
rect 30281 4450 30347 4453
rect 37457 4450 37523 4453
rect 38929 4450 38995 4453
rect 30281 4448 38995 4450
rect 30281 4392 30286 4448
rect 30342 4392 37462 4448
rect 37518 4392 38934 4448
rect 38990 4392 38995 4448
rect 30281 4390 38995 4392
rect 30281 4387 30347 4390
rect 37457 4387 37523 4390
rect 38929 4387 38995 4390
rect 15394 4384 15710 4385
rect 15394 4320 15400 4384
rect 15464 4320 15480 4384
rect 15544 4320 15560 4384
rect 15624 4320 15640 4384
rect 15704 4320 15710 4384
rect 15394 4319 15710 4320
rect 29842 4384 30158 4385
rect 29842 4320 29848 4384
rect 29912 4320 29928 4384
rect 29992 4320 30008 4384
rect 30072 4320 30088 4384
rect 30152 4320 30158 4384
rect 29842 4319 30158 4320
rect 44290 4384 44606 4385
rect 44290 4320 44296 4384
rect 44360 4320 44376 4384
rect 44440 4320 44456 4384
rect 44520 4320 44536 4384
rect 44600 4320 44606 4384
rect 44290 4319 44606 4320
rect 6821 4314 6887 4317
rect 6821 4312 15210 4314
rect 6821 4256 6826 4312
rect 6882 4256 15210 4312
rect 6821 4254 15210 4256
rect 6821 4251 6887 4254
rect 7649 4178 7715 4181
rect 13997 4178 14063 4181
rect 7649 4176 14063 4178
rect 7649 4120 7654 4176
rect 7710 4120 14002 4176
rect 14058 4120 14063 4176
rect 7649 4118 14063 4120
rect 15150 4178 15210 4254
rect 15653 4178 15719 4181
rect 15150 4176 15719 4178
rect 15150 4120 15658 4176
rect 15714 4120 15719 4176
rect 15150 4118 15719 4120
rect 7649 4115 7715 4118
rect 13997 4115 14063 4118
rect 15653 4115 15719 4118
rect 19057 4178 19123 4181
rect 24945 4178 25011 4181
rect 19057 4176 25011 4178
rect 19057 4120 19062 4176
rect 19118 4120 24950 4176
rect 25006 4120 25011 4176
rect 19057 4118 25011 4120
rect 19057 4115 19123 4118
rect 24945 4115 25011 4118
rect 17861 4042 17927 4045
rect 20713 4042 20779 4045
rect 17861 4040 20779 4042
rect 17861 3984 17866 4040
rect 17922 3984 20718 4040
rect 20774 3984 20779 4040
rect 17861 3982 20779 3984
rect 17861 3979 17927 3982
rect 20713 3979 20779 3982
rect 24853 4042 24919 4045
rect 25497 4042 25563 4045
rect 25773 4042 25839 4045
rect 44081 4042 44147 4045
rect 24853 4040 44147 4042
rect 24853 3984 24858 4040
rect 24914 3984 25502 4040
rect 25558 3984 25778 4040
rect 25834 3984 44086 4040
rect 44142 3984 44147 4040
rect 24853 3982 44147 3984
rect 24853 3979 24919 3982
rect 25497 3979 25563 3982
rect 25773 3979 25839 3982
rect 44081 3979 44147 3982
rect 44265 4042 44331 4045
rect 49049 4042 49115 4045
rect 44265 4040 49115 4042
rect 44265 3984 44270 4040
rect 44326 3984 49054 4040
rect 49110 3984 49115 4040
rect 44265 3982 49115 3984
rect 44265 3979 44331 3982
rect 49049 3979 49115 3982
rect 12157 3906 12223 3909
rect 19333 3906 19399 3909
rect 12157 3904 19399 3906
rect 12157 3848 12162 3904
rect 12218 3848 19338 3904
rect 19394 3848 19399 3904
rect 12157 3846 19399 3848
rect 12157 3843 12223 3846
rect 19333 3843 19399 3846
rect 32765 3906 32831 3909
rect 35893 3906 35959 3909
rect 32765 3904 35959 3906
rect 32765 3848 32770 3904
rect 32826 3848 35898 3904
rect 35954 3848 35959 3904
rect 32765 3846 35959 3848
rect 32765 3843 32831 3846
rect 35893 3843 35959 3846
rect 40585 3906 40651 3909
rect 43069 3906 43135 3909
rect 51257 3906 51323 3909
rect 40585 3904 51323 3906
rect 40585 3848 40590 3904
rect 40646 3848 43074 3904
rect 43130 3848 51262 3904
rect 51318 3848 51323 3904
rect 40585 3846 51323 3848
rect 40585 3843 40651 3846
rect 43069 3843 43135 3846
rect 51257 3843 51323 3846
rect 8170 3840 8486 3841
rect 8170 3776 8176 3840
rect 8240 3776 8256 3840
rect 8320 3776 8336 3840
rect 8400 3776 8416 3840
rect 8480 3776 8486 3840
rect 8170 3775 8486 3776
rect 22618 3840 22934 3841
rect 22618 3776 22624 3840
rect 22688 3776 22704 3840
rect 22768 3776 22784 3840
rect 22848 3776 22864 3840
rect 22928 3776 22934 3840
rect 22618 3775 22934 3776
rect 37066 3840 37382 3841
rect 37066 3776 37072 3840
rect 37136 3776 37152 3840
rect 37216 3776 37232 3840
rect 37296 3776 37312 3840
rect 37376 3776 37382 3840
rect 37066 3775 37382 3776
rect 51514 3840 51830 3841
rect 51514 3776 51520 3840
rect 51584 3776 51600 3840
rect 51664 3776 51680 3840
rect 51744 3776 51760 3840
rect 51824 3776 51830 3840
rect 51514 3775 51830 3776
rect 12934 3708 12940 3772
rect 13004 3770 13010 3772
rect 13077 3770 13143 3773
rect 38653 3770 38719 3773
rect 13004 3768 13143 3770
rect 13004 3712 13082 3768
rect 13138 3712 13143 3768
rect 13004 3710 13143 3712
rect 13004 3708 13010 3710
rect 13077 3707 13143 3710
rect 37598 3768 38719 3770
rect 37598 3712 38658 3768
rect 38714 3712 38719 3768
rect 37598 3710 38719 3712
rect 4429 3634 4495 3637
rect 12341 3634 12407 3637
rect 13905 3634 13971 3637
rect 34421 3634 34487 3637
rect 35985 3634 36051 3637
rect 37598 3634 37658 3710
rect 38653 3707 38719 3710
rect 38837 3770 38903 3773
rect 47577 3770 47643 3773
rect 38837 3768 47643 3770
rect 38837 3712 38842 3768
rect 38898 3712 47582 3768
rect 47638 3712 47643 3768
rect 38837 3710 47643 3712
rect 38837 3707 38903 3710
rect 47577 3707 47643 3710
rect 4429 3632 16590 3634
rect 4429 3576 4434 3632
rect 4490 3576 12346 3632
rect 12402 3576 13910 3632
rect 13966 3576 16590 3632
rect 4429 3574 16590 3576
rect 4429 3571 4495 3574
rect 12341 3571 12407 3574
rect 13905 3571 13971 3574
rect 5441 3498 5507 3501
rect 13353 3498 13419 3501
rect 5441 3496 13419 3498
rect 5441 3440 5446 3496
rect 5502 3440 13358 3496
rect 13414 3440 13419 3496
rect 5441 3438 13419 3440
rect 16530 3498 16590 3574
rect 34421 3632 37658 3634
rect 34421 3576 34426 3632
rect 34482 3576 35990 3632
rect 36046 3576 37658 3632
rect 34421 3574 37658 3576
rect 37733 3634 37799 3637
rect 44633 3634 44699 3637
rect 37733 3632 44699 3634
rect 37733 3576 37738 3632
rect 37794 3576 44638 3632
rect 44694 3576 44699 3632
rect 37733 3574 44699 3576
rect 34421 3571 34487 3574
rect 35985 3571 36051 3574
rect 37733 3571 37799 3574
rect 44633 3571 44699 3574
rect 47025 3634 47091 3637
rect 54477 3634 54543 3637
rect 47025 3632 54543 3634
rect 47025 3576 47030 3632
rect 47086 3576 54482 3632
rect 54538 3576 54543 3632
rect 47025 3574 54543 3576
rect 47025 3571 47091 3574
rect 54477 3571 54543 3574
rect 19701 3498 19767 3501
rect 16530 3496 19767 3498
rect 16530 3440 19706 3496
rect 19762 3440 19767 3496
rect 16530 3438 19767 3440
rect 5441 3435 5507 3438
rect 13353 3435 13419 3438
rect 19701 3435 19767 3438
rect 26049 3498 26115 3501
rect 36077 3498 36143 3501
rect 39757 3498 39823 3501
rect 26049 3496 39823 3498
rect 26049 3440 26054 3496
rect 26110 3440 36082 3496
rect 36138 3440 39762 3496
rect 39818 3440 39823 3496
rect 26049 3438 39823 3440
rect 26049 3435 26115 3438
rect 36077 3435 36143 3438
rect 39757 3435 39823 3438
rect 44081 3498 44147 3501
rect 45185 3498 45251 3501
rect 55857 3498 55923 3501
rect 44081 3496 45018 3498
rect 44081 3440 44086 3496
rect 44142 3440 45018 3496
rect 44081 3438 45018 3440
rect 44081 3435 44147 3438
rect 3141 3362 3207 3365
rect 9673 3362 9739 3365
rect 3141 3360 9739 3362
rect 3141 3304 3146 3360
rect 3202 3304 9678 3360
rect 9734 3304 9739 3360
rect 3141 3302 9739 3304
rect 3141 3299 3207 3302
rect 9673 3299 9739 3302
rect 30465 3362 30531 3365
rect 34053 3362 34119 3365
rect 30465 3360 34119 3362
rect 30465 3304 30470 3360
rect 30526 3304 34058 3360
rect 34114 3304 34119 3360
rect 30465 3302 34119 3304
rect 44958 3362 45018 3438
rect 45185 3496 55923 3498
rect 45185 3440 45190 3496
rect 45246 3440 55862 3496
rect 55918 3440 55923 3496
rect 45185 3438 55923 3440
rect 45185 3435 45251 3438
rect 55857 3435 55923 3438
rect 46933 3362 46999 3365
rect 50061 3362 50127 3365
rect 44958 3360 50127 3362
rect 44958 3304 46938 3360
rect 46994 3304 50066 3360
rect 50122 3304 50127 3360
rect 44958 3302 50127 3304
rect 30465 3299 30531 3302
rect 34053 3299 34119 3302
rect 46933 3299 46999 3302
rect 50061 3299 50127 3302
rect 15394 3296 15710 3297
rect 15394 3232 15400 3296
rect 15464 3232 15480 3296
rect 15544 3232 15560 3296
rect 15624 3232 15640 3296
rect 15704 3232 15710 3296
rect 15394 3231 15710 3232
rect 29842 3296 30158 3297
rect 29842 3232 29848 3296
rect 29912 3232 29928 3296
rect 29992 3232 30008 3296
rect 30072 3232 30088 3296
rect 30152 3232 30158 3296
rect 29842 3231 30158 3232
rect 44290 3296 44606 3297
rect 44290 3232 44296 3296
rect 44360 3232 44376 3296
rect 44440 3232 44456 3296
rect 44520 3232 44536 3296
rect 44600 3232 44606 3296
rect 44290 3231 44606 3232
rect 8753 3226 8819 3229
rect 13261 3226 13327 3229
rect 8753 3224 13327 3226
rect 8753 3168 8758 3224
rect 8814 3168 13266 3224
rect 13322 3168 13327 3224
rect 8753 3166 13327 3168
rect 8753 3163 8819 3166
rect 13261 3163 13327 3166
rect 21725 3226 21791 3229
rect 28257 3226 28323 3229
rect 21725 3224 28323 3226
rect 21725 3168 21730 3224
rect 21786 3168 28262 3224
rect 28318 3168 28323 3224
rect 21725 3166 28323 3168
rect 21725 3163 21791 3166
rect 28257 3163 28323 3166
rect 8753 3090 8819 3093
rect 19793 3090 19859 3093
rect 8753 3088 19859 3090
rect 8753 3032 8758 3088
rect 8814 3032 19798 3088
rect 19854 3032 19859 3088
rect 8753 3030 19859 3032
rect 8753 3027 8819 3030
rect 19793 3027 19859 3030
rect 19977 3090 20043 3093
rect 27245 3090 27311 3093
rect 19977 3088 27311 3090
rect 19977 3032 19982 3088
rect 20038 3032 27250 3088
rect 27306 3032 27311 3088
rect 19977 3030 27311 3032
rect 19977 3027 20043 3030
rect 27245 3027 27311 3030
rect 36353 3090 36419 3093
rect 42885 3090 42951 3093
rect 51165 3090 51231 3093
rect 36353 3088 51231 3090
rect 36353 3032 36358 3088
rect 36414 3032 42890 3088
rect 42946 3032 51170 3088
rect 51226 3032 51231 3088
rect 36353 3030 51231 3032
rect 36353 3027 36419 3030
rect 42885 3027 42951 3030
rect 51165 3027 51231 3030
rect 18597 2954 18663 2957
rect 21725 2954 21791 2957
rect 18597 2952 21791 2954
rect 18597 2896 18602 2952
rect 18658 2896 21730 2952
rect 21786 2896 21791 2952
rect 18597 2894 21791 2896
rect 18597 2891 18663 2894
rect 21725 2891 21791 2894
rect 26693 2954 26759 2957
rect 46565 2954 46631 2957
rect 26693 2952 46631 2954
rect 26693 2896 26698 2952
rect 26754 2896 46570 2952
rect 46626 2896 46631 2952
rect 26693 2894 46631 2896
rect 26693 2891 26759 2894
rect 46565 2891 46631 2894
rect 10777 2818 10843 2821
rect 15285 2818 15351 2821
rect 10777 2816 15351 2818
rect 10777 2760 10782 2816
rect 10838 2760 15290 2816
rect 15346 2760 15351 2816
rect 10777 2758 15351 2760
rect 10777 2755 10843 2758
rect 15285 2755 15351 2758
rect 8170 2752 8486 2753
rect 8170 2688 8176 2752
rect 8240 2688 8256 2752
rect 8320 2688 8336 2752
rect 8400 2688 8416 2752
rect 8480 2688 8486 2752
rect 8170 2687 8486 2688
rect 22618 2752 22934 2753
rect 22618 2688 22624 2752
rect 22688 2688 22704 2752
rect 22768 2688 22784 2752
rect 22848 2688 22864 2752
rect 22928 2688 22934 2752
rect 22618 2687 22934 2688
rect 37066 2752 37382 2753
rect 37066 2688 37072 2752
rect 37136 2688 37152 2752
rect 37216 2688 37232 2752
rect 37296 2688 37312 2752
rect 37376 2688 37382 2752
rect 37066 2687 37382 2688
rect 51514 2752 51830 2753
rect 51514 2688 51520 2752
rect 51584 2688 51600 2752
rect 51664 2688 51680 2752
rect 51744 2688 51760 2752
rect 51824 2688 51830 2752
rect 51514 2687 51830 2688
rect 4061 2546 4127 2549
rect 12934 2546 12940 2548
rect 4061 2544 12940 2546
rect 4061 2488 4066 2544
rect 4122 2488 12940 2544
rect 4061 2486 12940 2488
rect 4061 2483 4127 2486
rect 12934 2484 12940 2486
rect 13004 2484 13010 2548
rect 26877 2546 26943 2549
rect 50153 2546 50219 2549
rect 26877 2544 50219 2546
rect 26877 2488 26882 2544
rect 26938 2488 50158 2544
rect 50214 2488 50219 2544
rect 26877 2486 50219 2488
rect 26877 2483 26943 2486
rect 50153 2483 50219 2486
rect 27245 2410 27311 2413
rect 47117 2410 47183 2413
rect 27245 2408 47183 2410
rect 27245 2352 27250 2408
rect 27306 2352 47122 2408
rect 47178 2352 47183 2408
rect 27245 2350 47183 2352
rect 27245 2347 27311 2350
rect 47117 2347 47183 2350
rect 15394 2208 15710 2209
rect 15394 2144 15400 2208
rect 15464 2144 15480 2208
rect 15544 2144 15560 2208
rect 15624 2144 15640 2208
rect 15704 2144 15710 2208
rect 15394 2143 15710 2144
rect 29842 2208 30158 2209
rect 29842 2144 29848 2208
rect 29912 2144 29928 2208
rect 29992 2144 30008 2208
rect 30072 2144 30088 2208
rect 30152 2144 30158 2208
rect 29842 2143 30158 2144
rect 44290 2208 44606 2209
rect 44290 2144 44296 2208
rect 44360 2144 44376 2208
rect 44440 2144 44456 2208
rect 44520 2144 44536 2208
rect 44600 2144 44606 2208
rect 44290 2143 44606 2144
rect 7281 2002 7347 2005
rect 23473 2002 23539 2005
rect 7281 2000 23539 2002
rect 7281 1944 7286 2000
rect 7342 1944 23478 2000
rect 23534 1944 23539 2000
rect 7281 1942 23539 1944
rect 7281 1939 7347 1942
rect 23473 1939 23539 1942
rect 12157 1866 12223 1869
rect 38745 1866 38811 1869
rect 12157 1864 38811 1866
rect 12157 1808 12162 1864
rect 12218 1808 38750 1864
rect 38806 1808 38811 1864
rect 12157 1806 38811 1808
rect 12157 1803 12223 1806
rect 38745 1803 38811 1806
rect 9397 1730 9463 1733
rect 28349 1730 28415 1733
rect 9397 1728 28415 1730
rect 9397 1672 9402 1728
rect 9458 1672 28354 1728
rect 28410 1672 28415 1728
rect 9397 1670 28415 1672
rect 9397 1667 9463 1670
rect 28349 1667 28415 1670
<< via3 >>
rect 15400 7644 15464 7648
rect 15400 7588 15404 7644
rect 15404 7588 15460 7644
rect 15460 7588 15464 7644
rect 15400 7584 15464 7588
rect 15480 7644 15544 7648
rect 15480 7588 15484 7644
rect 15484 7588 15540 7644
rect 15540 7588 15544 7644
rect 15480 7584 15544 7588
rect 15560 7644 15624 7648
rect 15560 7588 15564 7644
rect 15564 7588 15620 7644
rect 15620 7588 15624 7644
rect 15560 7584 15624 7588
rect 15640 7644 15704 7648
rect 15640 7588 15644 7644
rect 15644 7588 15700 7644
rect 15700 7588 15704 7644
rect 15640 7584 15704 7588
rect 29848 7644 29912 7648
rect 29848 7588 29852 7644
rect 29852 7588 29908 7644
rect 29908 7588 29912 7644
rect 29848 7584 29912 7588
rect 29928 7644 29992 7648
rect 29928 7588 29932 7644
rect 29932 7588 29988 7644
rect 29988 7588 29992 7644
rect 29928 7584 29992 7588
rect 30008 7644 30072 7648
rect 30008 7588 30012 7644
rect 30012 7588 30068 7644
rect 30068 7588 30072 7644
rect 30008 7584 30072 7588
rect 30088 7644 30152 7648
rect 30088 7588 30092 7644
rect 30092 7588 30148 7644
rect 30148 7588 30152 7644
rect 30088 7584 30152 7588
rect 44296 7644 44360 7648
rect 44296 7588 44300 7644
rect 44300 7588 44356 7644
rect 44356 7588 44360 7644
rect 44296 7584 44360 7588
rect 44376 7644 44440 7648
rect 44376 7588 44380 7644
rect 44380 7588 44436 7644
rect 44436 7588 44440 7644
rect 44376 7584 44440 7588
rect 44456 7644 44520 7648
rect 44456 7588 44460 7644
rect 44460 7588 44516 7644
rect 44516 7588 44520 7644
rect 44456 7584 44520 7588
rect 44536 7644 44600 7648
rect 44536 7588 44540 7644
rect 44540 7588 44596 7644
rect 44596 7588 44600 7644
rect 44536 7584 44600 7588
rect 8176 7100 8240 7104
rect 8176 7044 8180 7100
rect 8180 7044 8236 7100
rect 8236 7044 8240 7100
rect 8176 7040 8240 7044
rect 8256 7100 8320 7104
rect 8256 7044 8260 7100
rect 8260 7044 8316 7100
rect 8316 7044 8320 7100
rect 8256 7040 8320 7044
rect 8336 7100 8400 7104
rect 8336 7044 8340 7100
rect 8340 7044 8396 7100
rect 8396 7044 8400 7100
rect 8336 7040 8400 7044
rect 8416 7100 8480 7104
rect 8416 7044 8420 7100
rect 8420 7044 8476 7100
rect 8476 7044 8480 7100
rect 8416 7040 8480 7044
rect 22624 7100 22688 7104
rect 22624 7044 22628 7100
rect 22628 7044 22684 7100
rect 22684 7044 22688 7100
rect 22624 7040 22688 7044
rect 22704 7100 22768 7104
rect 22704 7044 22708 7100
rect 22708 7044 22764 7100
rect 22764 7044 22768 7100
rect 22704 7040 22768 7044
rect 22784 7100 22848 7104
rect 22784 7044 22788 7100
rect 22788 7044 22844 7100
rect 22844 7044 22848 7100
rect 22784 7040 22848 7044
rect 22864 7100 22928 7104
rect 22864 7044 22868 7100
rect 22868 7044 22924 7100
rect 22924 7044 22928 7100
rect 22864 7040 22928 7044
rect 37072 7100 37136 7104
rect 37072 7044 37076 7100
rect 37076 7044 37132 7100
rect 37132 7044 37136 7100
rect 37072 7040 37136 7044
rect 37152 7100 37216 7104
rect 37152 7044 37156 7100
rect 37156 7044 37212 7100
rect 37212 7044 37216 7100
rect 37152 7040 37216 7044
rect 37232 7100 37296 7104
rect 37232 7044 37236 7100
rect 37236 7044 37292 7100
rect 37292 7044 37296 7100
rect 37232 7040 37296 7044
rect 37312 7100 37376 7104
rect 37312 7044 37316 7100
rect 37316 7044 37372 7100
rect 37372 7044 37376 7100
rect 37312 7040 37376 7044
rect 51520 7100 51584 7104
rect 51520 7044 51524 7100
rect 51524 7044 51580 7100
rect 51580 7044 51584 7100
rect 51520 7040 51584 7044
rect 51600 7100 51664 7104
rect 51600 7044 51604 7100
rect 51604 7044 51660 7100
rect 51660 7044 51664 7100
rect 51600 7040 51664 7044
rect 51680 7100 51744 7104
rect 51680 7044 51684 7100
rect 51684 7044 51740 7100
rect 51740 7044 51744 7100
rect 51680 7040 51744 7044
rect 51760 7100 51824 7104
rect 51760 7044 51764 7100
rect 51764 7044 51820 7100
rect 51820 7044 51824 7100
rect 51760 7040 51824 7044
rect 15400 6556 15464 6560
rect 15400 6500 15404 6556
rect 15404 6500 15460 6556
rect 15460 6500 15464 6556
rect 15400 6496 15464 6500
rect 15480 6556 15544 6560
rect 15480 6500 15484 6556
rect 15484 6500 15540 6556
rect 15540 6500 15544 6556
rect 15480 6496 15544 6500
rect 15560 6556 15624 6560
rect 15560 6500 15564 6556
rect 15564 6500 15620 6556
rect 15620 6500 15624 6556
rect 15560 6496 15624 6500
rect 15640 6556 15704 6560
rect 15640 6500 15644 6556
rect 15644 6500 15700 6556
rect 15700 6500 15704 6556
rect 15640 6496 15704 6500
rect 29848 6556 29912 6560
rect 29848 6500 29852 6556
rect 29852 6500 29908 6556
rect 29908 6500 29912 6556
rect 29848 6496 29912 6500
rect 29928 6556 29992 6560
rect 29928 6500 29932 6556
rect 29932 6500 29988 6556
rect 29988 6500 29992 6556
rect 29928 6496 29992 6500
rect 30008 6556 30072 6560
rect 30008 6500 30012 6556
rect 30012 6500 30068 6556
rect 30068 6500 30072 6556
rect 30008 6496 30072 6500
rect 30088 6556 30152 6560
rect 30088 6500 30092 6556
rect 30092 6500 30148 6556
rect 30148 6500 30152 6556
rect 30088 6496 30152 6500
rect 44296 6556 44360 6560
rect 44296 6500 44300 6556
rect 44300 6500 44356 6556
rect 44356 6500 44360 6556
rect 44296 6496 44360 6500
rect 44376 6556 44440 6560
rect 44376 6500 44380 6556
rect 44380 6500 44436 6556
rect 44436 6500 44440 6556
rect 44376 6496 44440 6500
rect 44456 6556 44520 6560
rect 44456 6500 44460 6556
rect 44460 6500 44516 6556
rect 44516 6500 44520 6556
rect 44456 6496 44520 6500
rect 44536 6556 44600 6560
rect 44536 6500 44540 6556
rect 44540 6500 44596 6556
rect 44596 6500 44600 6556
rect 44536 6496 44600 6500
rect 8176 6012 8240 6016
rect 8176 5956 8180 6012
rect 8180 5956 8236 6012
rect 8236 5956 8240 6012
rect 8176 5952 8240 5956
rect 8256 6012 8320 6016
rect 8256 5956 8260 6012
rect 8260 5956 8316 6012
rect 8316 5956 8320 6012
rect 8256 5952 8320 5956
rect 8336 6012 8400 6016
rect 8336 5956 8340 6012
rect 8340 5956 8396 6012
rect 8396 5956 8400 6012
rect 8336 5952 8400 5956
rect 8416 6012 8480 6016
rect 8416 5956 8420 6012
rect 8420 5956 8476 6012
rect 8476 5956 8480 6012
rect 8416 5952 8480 5956
rect 22624 6012 22688 6016
rect 22624 5956 22628 6012
rect 22628 5956 22684 6012
rect 22684 5956 22688 6012
rect 22624 5952 22688 5956
rect 22704 6012 22768 6016
rect 22704 5956 22708 6012
rect 22708 5956 22764 6012
rect 22764 5956 22768 6012
rect 22704 5952 22768 5956
rect 22784 6012 22848 6016
rect 22784 5956 22788 6012
rect 22788 5956 22844 6012
rect 22844 5956 22848 6012
rect 22784 5952 22848 5956
rect 22864 6012 22928 6016
rect 22864 5956 22868 6012
rect 22868 5956 22924 6012
rect 22924 5956 22928 6012
rect 22864 5952 22928 5956
rect 37072 6012 37136 6016
rect 37072 5956 37076 6012
rect 37076 5956 37132 6012
rect 37132 5956 37136 6012
rect 37072 5952 37136 5956
rect 37152 6012 37216 6016
rect 37152 5956 37156 6012
rect 37156 5956 37212 6012
rect 37212 5956 37216 6012
rect 37152 5952 37216 5956
rect 37232 6012 37296 6016
rect 37232 5956 37236 6012
rect 37236 5956 37292 6012
rect 37292 5956 37296 6012
rect 37232 5952 37296 5956
rect 37312 6012 37376 6016
rect 37312 5956 37316 6012
rect 37316 5956 37372 6012
rect 37372 5956 37376 6012
rect 37312 5952 37376 5956
rect 51520 6012 51584 6016
rect 51520 5956 51524 6012
rect 51524 5956 51580 6012
rect 51580 5956 51584 6012
rect 51520 5952 51584 5956
rect 51600 6012 51664 6016
rect 51600 5956 51604 6012
rect 51604 5956 51660 6012
rect 51660 5956 51664 6012
rect 51600 5952 51664 5956
rect 51680 6012 51744 6016
rect 51680 5956 51684 6012
rect 51684 5956 51740 6012
rect 51740 5956 51744 6012
rect 51680 5952 51744 5956
rect 51760 6012 51824 6016
rect 51760 5956 51764 6012
rect 51764 5956 51820 6012
rect 51820 5956 51824 6012
rect 51760 5952 51824 5956
rect 15400 5468 15464 5472
rect 15400 5412 15404 5468
rect 15404 5412 15460 5468
rect 15460 5412 15464 5468
rect 15400 5408 15464 5412
rect 15480 5468 15544 5472
rect 15480 5412 15484 5468
rect 15484 5412 15540 5468
rect 15540 5412 15544 5468
rect 15480 5408 15544 5412
rect 15560 5468 15624 5472
rect 15560 5412 15564 5468
rect 15564 5412 15620 5468
rect 15620 5412 15624 5468
rect 15560 5408 15624 5412
rect 15640 5468 15704 5472
rect 15640 5412 15644 5468
rect 15644 5412 15700 5468
rect 15700 5412 15704 5468
rect 15640 5408 15704 5412
rect 29848 5468 29912 5472
rect 29848 5412 29852 5468
rect 29852 5412 29908 5468
rect 29908 5412 29912 5468
rect 29848 5408 29912 5412
rect 29928 5468 29992 5472
rect 29928 5412 29932 5468
rect 29932 5412 29988 5468
rect 29988 5412 29992 5468
rect 29928 5408 29992 5412
rect 30008 5468 30072 5472
rect 30008 5412 30012 5468
rect 30012 5412 30068 5468
rect 30068 5412 30072 5468
rect 30008 5408 30072 5412
rect 30088 5468 30152 5472
rect 30088 5412 30092 5468
rect 30092 5412 30148 5468
rect 30148 5412 30152 5468
rect 30088 5408 30152 5412
rect 44296 5468 44360 5472
rect 44296 5412 44300 5468
rect 44300 5412 44356 5468
rect 44356 5412 44360 5468
rect 44296 5408 44360 5412
rect 44376 5468 44440 5472
rect 44376 5412 44380 5468
rect 44380 5412 44436 5468
rect 44436 5412 44440 5468
rect 44376 5408 44440 5412
rect 44456 5468 44520 5472
rect 44456 5412 44460 5468
rect 44460 5412 44516 5468
rect 44516 5412 44520 5468
rect 44456 5408 44520 5412
rect 44536 5468 44600 5472
rect 44536 5412 44540 5468
rect 44540 5412 44596 5468
rect 44596 5412 44600 5468
rect 44536 5408 44600 5412
rect 8176 4924 8240 4928
rect 8176 4868 8180 4924
rect 8180 4868 8236 4924
rect 8236 4868 8240 4924
rect 8176 4864 8240 4868
rect 8256 4924 8320 4928
rect 8256 4868 8260 4924
rect 8260 4868 8316 4924
rect 8316 4868 8320 4924
rect 8256 4864 8320 4868
rect 8336 4924 8400 4928
rect 8336 4868 8340 4924
rect 8340 4868 8396 4924
rect 8396 4868 8400 4924
rect 8336 4864 8400 4868
rect 8416 4924 8480 4928
rect 8416 4868 8420 4924
rect 8420 4868 8476 4924
rect 8476 4868 8480 4924
rect 8416 4864 8480 4868
rect 22624 4924 22688 4928
rect 22624 4868 22628 4924
rect 22628 4868 22684 4924
rect 22684 4868 22688 4924
rect 22624 4864 22688 4868
rect 22704 4924 22768 4928
rect 22704 4868 22708 4924
rect 22708 4868 22764 4924
rect 22764 4868 22768 4924
rect 22704 4864 22768 4868
rect 22784 4924 22848 4928
rect 22784 4868 22788 4924
rect 22788 4868 22844 4924
rect 22844 4868 22848 4924
rect 22784 4864 22848 4868
rect 22864 4924 22928 4928
rect 22864 4868 22868 4924
rect 22868 4868 22924 4924
rect 22924 4868 22928 4924
rect 22864 4864 22928 4868
rect 37072 4924 37136 4928
rect 37072 4868 37076 4924
rect 37076 4868 37132 4924
rect 37132 4868 37136 4924
rect 37072 4864 37136 4868
rect 37152 4924 37216 4928
rect 37152 4868 37156 4924
rect 37156 4868 37212 4924
rect 37212 4868 37216 4924
rect 37152 4864 37216 4868
rect 37232 4924 37296 4928
rect 37232 4868 37236 4924
rect 37236 4868 37292 4924
rect 37292 4868 37296 4924
rect 37232 4864 37296 4868
rect 37312 4924 37376 4928
rect 37312 4868 37316 4924
rect 37316 4868 37372 4924
rect 37372 4868 37376 4924
rect 37312 4864 37376 4868
rect 51520 4924 51584 4928
rect 51520 4868 51524 4924
rect 51524 4868 51580 4924
rect 51580 4868 51584 4924
rect 51520 4864 51584 4868
rect 51600 4924 51664 4928
rect 51600 4868 51604 4924
rect 51604 4868 51660 4924
rect 51660 4868 51664 4924
rect 51600 4864 51664 4868
rect 51680 4924 51744 4928
rect 51680 4868 51684 4924
rect 51684 4868 51740 4924
rect 51740 4868 51744 4924
rect 51680 4864 51744 4868
rect 51760 4924 51824 4928
rect 51760 4868 51764 4924
rect 51764 4868 51820 4924
rect 51820 4868 51824 4924
rect 51760 4864 51824 4868
rect 12940 4660 13004 4724
rect 15400 4380 15464 4384
rect 15400 4324 15404 4380
rect 15404 4324 15460 4380
rect 15460 4324 15464 4380
rect 15400 4320 15464 4324
rect 15480 4380 15544 4384
rect 15480 4324 15484 4380
rect 15484 4324 15540 4380
rect 15540 4324 15544 4380
rect 15480 4320 15544 4324
rect 15560 4380 15624 4384
rect 15560 4324 15564 4380
rect 15564 4324 15620 4380
rect 15620 4324 15624 4380
rect 15560 4320 15624 4324
rect 15640 4380 15704 4384
rect 15640 4324 15644 4380
rect 15644 4324 15700 4380
rect 15700 4324 15704 4380
rect 15640 4320 15704 4324
rect 29848 4380 29912 4384
rect 29848 4324 29852 4380
rect 29852 4324 29908 4380
rect 29908 4324 29912 4380
rect 29848 4320 29912 4324
rect 29928 4380 29992 4384
rect 29928 4324 29932 4380
rect 29932 4324 29988 4380
rect 29988 4324 29992 4380
rect 29928 4320 29992 4324
rect 30008 4380 30072 4384
rect 30008 4324 30012 4380
rect 30012 4324 30068 4380
rect 30068 4324 30072 4380
rect 30008 4320 30072 4324
rect 30088 4380 30152 4384
rect 30088 4324 30092 4380
rect 30092 4324 30148 4380
rect 30148 4324 30152 4380
rect 30088 4320 30152 4324
rect 44296 4380 44360 4384
rect 44296 4324 44300 4380
rect 44300 4324 44356 4380
rect 44356 4324 44360 4380
rect 44296 4320 44360 4324
rect 44376 4380 44440 4384
rect 44376 4324 44380 4380
rect 44380 4324 44436 4380
rect 44436 4324 44440 4380
rect 44376 4320 44440 4324
rect 44456 4380 44520 4384
rect 44456 4324 44460 4380
rect 44460 4324 44516 4380
rect 44516 4324 44520 4380
rect 44456 4320 44520 4324
rect 44536 4380 44600 4384
rect 44536 4324 44540 4380
rect 44540 4324 44596 4380
rect 44596 4324 44600 4380
rect 44536 4320 44600 4324
rect 8176 3836 8240 3840
rect 8176 3780 8180 3836
rect 8180 3780 8236 3836
rect 8236 3780 8240 3836
rect 8176 3776 8240 3780
rect 8256 3836 8320 3840
rect 8256 3780 8260 3836
rect 8260 3780 8316 3836
rect 8316 3780 8320 3836
rect 8256 3776 8320 3780
rect 8336 3836 8400 3840
rect 8336 3780 8340 3836
rect 8340 3780 8396 3836
rect 8396 3780 8400 3836
rect 8336 3776 8400 3780
rect 8416 3836 8480 3840
rect 8416 3780 8420 3836
rect 8420 3780 8476 3836
rect 8476 3780 8480 3836
rect 8416 3776 8480 3780
rect 22624 3836 22688 3840
rect 22624 3780 22628 3836
rect 22628 3780 22684 3836
rect 22684 3780 22688 3836
rect 22624 3776 22688 3780
rect 22704 3836 22768 3840
rect 22704 3780 22708 3836
rect 22708 3780 22764 3836
rect 22764 3780 22768 3836
rect 22704 3776 22768 3780
rect 22784 3836 22848 3840
rect 22784 3780 22788 3836
rect 22788 3780 22844 3836
rect 22844 3780 22848 3836
rect 22784 3776 22848 3780
rect 22864 3836 22928 3840
rect 22864 3780 22868 3836
rect 22868 3780 22924 3836
rect 22924 3780 22928 3836
rect 22864 3776 22928 3780
rect 37072 3836 37136 3840
rect 37072 3780 37076 3836
rect 37076 3780 37132 3836
rect 37132 3780 37136 3836
rect 37072 3776 37136 3780
rect 37152 3836 37216 3840
rect 37152 3780 37156 3836
rect 37156 3780 37212 3836
rect 37212 3780 37216 3836
rect 37152 3776 37216 3780
rect 37232 3836 37296 3840
rect 37232 3780 37236 3836
rect 37236 3780 37292 3836
rect 37292 3780 37296 3836
rect 37232 3776 37296 3780
rect 37312 3836 37376 3840
rect 37312 3780 37316 3836
rect 37316 3780 37372 3836
rect 37372 3780 37376 3836
rect 37312 3776 37376 3780
rect 51520 3836 51584 3840
rect 51520 3780 51524 3836
rect 51524 3780 51580 3836
rect 51580 3780 51584 3836
rect 51520 3776 51584 3780
rect 51600 3836 51664 3840
rect 51600 3780 51604 3836
rect 51604 3780 51660 3836
rect 51660 3780 51664 3836
rect 51600 3776 51664 3780
rect 51680 3836 51744 3840
rect 51680 3780 51684 3836
rect 51684 3780 51740 3836
rect 51740 3780 51744 3836
rect 51680 3776 51744 3780
rect 51760 3836 51824 3840
rect 51760 3780 51764 3836
rect 51764 3780 51820 3836
rect 51820 3780 51824 3836
rect 51760 3776 51824 3780
rect 12940 3708 13004 3772
rect 15400 3292 15464 3296
rect 15400 3236 15404 3292
rect 15404 3236 15460 3292
rect 15460 3236 15464 3292
rect 15400 3232 15464 3236
rect 15480 3292 15544 3296
rect 15480 3236 15484 3292
rect 15484 3236 15540 3292
rect 15540 3236 15544 3292
rect 15480 3232 15544 3236
rect 15560 3292 15624 3296
rect 15560 3236 15564 3292
rect 15564 3236 15620 3292
rect 15620 3236 15624 3292
rect 15560 3232 15624 3236
rect 15640 3292 15704 3296
rect 15640 3236 15644 3292
rect 15644 3236 15700 3292
rect 15700 3236 15704 3292
rect 15640 3232 15704 3236
rect 29848 3292 29912 3296
rect 29848 3236 29852 3292
rect 29852 3236 29908 3292
rect 29908 3236 29912 3292
rect 29848 3232 29912 3236
rect 29928 3292 29992 3296
rect 29928 3236 29932 3292
rect 29932 3236 29988 3292
rect 29988 3236 29992 3292
rect 29928 3232 29992 3236
rect 30008 3292 30072 3296
rect 30008 3236 30012 3292
rect 30012 3236 30068 3292
rect 30068 3236 30072 3292
rect 30008 3232 30072 3236
rect 30088 3292 30152 3296
rect 30088 3236 30092 3292
rect 30092 3236 30148 3292
rect 30148 3236 30152 3292
rect 30088 3232 30152 3236
rect 44296 3292 44360 3296
rect 44296 3236 44300 3292
rect 44300 3236 44356 3292
rect 44356 3236 44360 3292
rect 44296 3232 44360 3236
rect 44376 3292 44440 3296
rect 44376 3236 44380 3292
rect 44380 3236 44436 3292
rect 44436 3236 44440 3292
rect 44376 3232 44440 3236
rect 44456 3292 44520 3296
rect 44456 3236 44460 3292
rect 44460 3236 44516 3292
rect 44516 3236 44520 3292
rect 44456 3232 44520 3236
rect 44536 3292 44600 3296
rect 44536 3236 44540 3292
rect 44540 3236 44596 3292
rect 44596 3236 44600 3292
rect 44536 3232 44600 3236
rect 8176 2748 8240 2752
rect 8176 2692 8180 2748
rect 8180 2692 8236 2748
rect 8236 2692 8240 2748
rect 8176 2688 8240 2692
rect 8256 2748 8320 2752
rect 8256 2692 8260 2748
rect 8260 2692 8316 2748
rect 8316 2692 8320 2748
rect 8256 2688 8320 2692
rect 8336 2748 8400 2752
rect 8336 2692 8340 2748
rect 8340 2692 8396 2748
rect 8396 2692 8400 2748
rect 8336 2688 8400 2692
rect 8416 2748 8480 2752
rect 8416 2692 8420 2748
rect 8420 2692 8476 2748
rect 8476 2692 8480 2748
rect 8416 2688 8480 2692
rect 22624 2748 22688 2752
rect 22624 2692 22628 2748
rect 22628 2692 22684 2748
rect 22684 2692 22688 2748
rect 22624 2688 22688 2692
rect 22704 2748 22768 2752
rect 22704 2692 22708 2748
rect 22708 2692 22764 2748
rect 22764 2692 22768 2748
rect 22704 2688 22768 2692
rect 22784 2748 22848 2752
rect 22784 2692 22788 2748
rect 22788 2692 22844 2748
rect 22844 2692 22848 2748
rect 22784 2688 22848 2692
rect 22864 2748 22928 2752
rect 22864 2692 22868 2748
rect 22868 2692 22924 2748
rect 22924 2692 22928 2748
rect 22864 2688 22928 2692
rect 37072 2748 37136 2752
rect 37072 2692 37076 2748
rect 37076 2692 37132 2748
rect 37132 2692 37136 2748
rect 37072 2688 37136 2692
rect 37152 2748 37216 2752
rect 37152 2692 37156 2748
rect 37156 2692 37212 2748
rect 37212 2692 37216 2748
rect 37152 2688 37216 2692
rect 37232 2748 37296 2752
rect 37232 2692 37236 2748
rect 37236 2692 37292 2748
rect 37292 2692 37296 2748
rect 37232 2688 37296 2692
rect 37312 2748 37376 2752
rect 37312 2692 37316 2748
rect 37316 2692 37372 2748
rect 37372 2692 37376 2748
rect 37312 2688 37376 2692
rect 51520 2748 51584 2752
rect 51520 2692 51524 2748
rect 51524 2692 51580 2748
rect 51580 2692 51584 2748
rect 51520 2688 51584 2692
rect 51600 2748 51664 2752
rect 51600 2692 51604 2748
rect 51604 2692 51660 2748
rect 51660 2692 51664 2748
rect 51600 2688 51664 2692
rect 51680 2748 51744 2752
rect 51680 2692 51684 2748
rect 51684 2692 51740 2748
rect 51740 2692 51744 2748
rect 51680 2688 51744 2692
rect 51760 2748 51824 2752
rect 51760 2692 51764 2748
rect 51764 2692 51820 2748
rect 51820 2692 51824 2748
rect 51760 2688 51824 2692
rect 12940 2484 13004 2548
rect 15400 2204 15464 2208
rect 15400 2148 15404 2204
rect 15404 2148 15460 2204
rect 15460 2148 15464 2204
rect 15400 2144 15464 2148
rect 15480 2204 15544 2208
rect 15480 2148 15484 2204
rect 15484 2148 15540 2204
rect 15540 2148 15544 2204
rect 15480 2144 15544 2148
rect 15560 2204 15624 2208
rect 15560 2148 15564 2204
rect 15564 2148 15620 2204
rect 15620 2148 15624 2204
rect 15560 2144 15624 2148
rect 15640 2204 15704 2208
rect 15640 2148 15644 2204
rect 15644 2148 15700 2204
rect 15700 2148 15704 2204
rect 15640 2144 15704 2148
rect 29848 2204 29912 2208
rect 29848 2148 29852 2204
rect 29852 2148 29908 2204
rect 29908 2148 29912 2204
rect 29848 2144 29912 2148
rect 29928 2204 29992 2208
rect 29928 2148 29932 2204
rect 29932 2148 29988 2204
rect 29988 2148 29992 2204
rect 29928 2144 29992 2148
rect 30008 2204 30072 2208
rect 30008 2148 30012 2204
rect 30012 2148 30068 2204
rect 30068 2148 30072 2204
rect 30008 2144 30072 2148
rect 30088 2204 30152 2208
rect 30088 2148 30092 2204
rect 30092 2148 30148 2204
rect 30148 2148 30152 2204
rect 30088 2144 30152 2148
rect 44296 2204 44360 2208
rect 44296 2148 44300 2204
rect 44300 2148 44356 2204
rect 44356 2148 44360 2204
rect 44296 2144 44360 2148
rect 44376 2204 44440 2208
rect 44376 2148 44380 2204
rect 44380 2148 44436 2204
rect 44436 2148 44440 2204
rect 44376 2144 44440 2148
rect 44456 2204 44520 2208
rect 44456 2148 44460 2204
rect 44460 2148 44516 2204
rect 44516 2148 44520 2204
rect 44456 2144 44520 2148
rect 44536 2204 44600 2208
rect 44536 2148 44540 2204
rect 44540 2148 44596 2204
rect 44596 2148 44600 2204
rect 44536 2144 44600 2148
<< metal4 >>
rect 8168 7104 8488 7664
rect 8168 7040 8176 7104
rect 8240 7040 8256 7104
rect 8320 7040 8336 7104
rect 8400 7040 8416 7104
rect 8480 7040 8488 7104
rect 8168 6016 8488 7040
rect 8168 5952 8176 6016
rect 8240 5952 8256 6016
rect 8320 5952 8336 6016
rect 8400 5952 8416 6016
rect 8480 5952 8488 6016
rect 8168 4928 8488 5952
rect 8168 4864 8176 4928
rect 8240 4864 8256 4928
rect 8320 4864 8336 4928
rect 8400 4864 8416 4928
rect 8480 4864 8488 4928
rect 8168 3840 8488 4864
rect 15392 7648 15712 7664
rect 15392 7584 15400 7648
rect 15464 7584 15480 7648
rect 15544 7584 15560 7648
rect 15624 7584 15640 7648
rect 15704 7584 15712 7648
rect 15392 6560 15712 7584
rect 15392 6496 15400 6560
rect 15464 6496 15480 6560
rect 15544 6496 15560 6560
rect 15624 6496 15640 6560
rect 15704 6496 15712 6560
rect 15392 5472 15712 6496
rect 15392 5408 15400 5472
rect 15464 5408 15480 5472
rect 15544 5408 15560 5472
rect 15624 5408 15640 5472
rect 15704 5408 15712 5472
rect 12939 4724 13005 4725
rect 12939 4660 12940 4724
rect 13004 4660 13005 4724
rect 12939 4659 13005 4660
rect 8168 3776 8176 3840
rect 8240 3776 8256 3840
rect 8320 3776 8336 3840
rect 8400 3776 8416 3840
rect 8480 3776 8488 3840
rect 8168 2752 8488 3776
rect 12942 3773 13002 4659
rect 15392 4384 15712 5408
rect 15392 4320 15400 4384
rect 15464 4320 15480 4384
rect 15544 4320 15560 4384
rect 15624 4320 15640 4384
rect 15704 4320 15712 4384
rect 12939 3772 13005 3773
rect 12939 3708 12940 3772
rect 13004 3708 13005 3772
rect 12939 3707 13005 3708
rect 8168 2688 8176 2752
rect 8240 2688 8256 2752
rect 8320 2688 8336 2752
rect 8400 2688 8416 2752
rect 8480 2688 8488 2752
rect 8168 2128 8488 2688
rect 12942 2549 13002 3707
rect 15392 3296 15712 4320
rect 15392 3232 15400 3296
rect 15464 3232 15480 3296
rect 15544 3232 15560 3296
rect 15624 3232 15640 3296
rect 15704 3232 15712 3296
rect 12939 2548 13005 2549
rect 12939 2484 12940 2548
rect 13004 2484 13005 2548
rect 12939 2483 13005 2484
rect 15392 2208 15712 3232
rect 15392 2144 15400 2208
rect 15464 2144 15480 2208
rect 15544 2144 15560 2208
rect 15624 2144 15640 2208
rect 15704 2144 15712 2208
rect 15392 2128 15712 2144
rect 22616 7104 22936 7664
rect 22616 7040 22624 7104
rect 22688 7040 22704 7104
rect 22768 7040 22784 7104
rect 22848 7040 22864 7104
rect 22928 7040 22936 7104
rect 22616 6016 22936 7040
rect 22616 5952 22624 6016
rect 22688 5952 22704 6016
rect 22768 5952 22784 6016
rect 22848 5952 22864 6016
rect 22928 5952 22936 6016
rect 22616 4928 22936 5952
rect 22616 4864 22624 4928
rect 22688 4864 22704 4928
rect 22768 4864 22784 4928
rect 22848 4864 22864 4928
rect 22928 4864 22936 4928
rect 22616 3840 22936 4864
rect 22616 3776 22624 3840
rect 22688 3776 22704 3840
rect 22768 3776 22784 3840
rect 22848 3776 22864 3840
rect 22928 3776 22936 3840
rect 22616 2752 22936 3776
rect 22616 2688 22624 2752
rect 22688 2688 22704 2752
rect 22768 2688 22784 2752
rect 22848 2688 22864 2752
rect 22928 2688 22936 2752
rect 22616 2128 22936 2688
rect 29840 7648 30160 7664
rect 29840 7584 29848 7648
rect 29912 7584 29928 7648
rect 29992 7584 30008 7648
rect 30072 7584 30088 7648
rect 30152 7584 30160 7648
rect 29840 6560 30160 7584
rect 29840 6496 29848 6560
rect 29912 6496 29928 6560
rect 29992 6496 30008 6560
rect 30072 6496 30088 6560
rect 30152 6496 30160 6560
rect 29840 5472 30160 6496
rect 29840 5408 29848 5472
rect 29912 5408 29928 5472
rect 29992 5408 30008 5472
rect 30072 5408 30088 5472
rect 30152 5408 30160 5472
rect 29840 4384 30160 5408
rect 29840 4320 29848 4384
rect 29912 4320 29928 4384
rect 29992 4320 30008 4384
rect 30072 4320 30088 4384
rect 30152 4320 30160 4384
rect 29840 3296 30160 4320
rect 29840 3232 29848 3296
rect 29912 3232 29928 3296
rect 29992 3232 30008 3296
rect 30072 3232 30088 3296
rect 30152 3232 30160 3296
rect 29840 2208 30160 3232
rect 29840 2144 29848 2208
rect 29912 2144 29928 2208
rect 29992 2144 30008 2208
rect 30072 2144 30088 2208
rect 30152 2144 30160 2208
rect 29840 2128 30160 2144
rect 37064 7104 37384 7664
rect 37064 7040 37072 7104
rect 37136 7040 37152 7104
rect 37216 7040 37232 7104
rect 37296 7040 37312 7104
rect 37376 7040 37384 7104
rect 37064 6016 37384 7040
rect 37064 5952 37072 6016
rect 37136 5952 37152 6016
rect 37216 5952 37232 6016
rect 37296 5952 37312 6016
rect 37376 5952 37384 6016
rect 37064 4928 37384 5952
rect 37064 4864 37072 4928
rect 37136 4864 37152 4928
rect 37216 4864 37232 4928
rect 37296 4864 37312 4928
rect 37376 4864 37384 4928
rect 37064 3840 37384 4864
rect 37064 3776 37072 3840
rect 37136 3776 37152 3840
rect 37216 3776 37232 3840
rect 37296 3776 37312 3840
rect 37376 3776 37384 3840
rect 37064 2752 37384 3776
rect 37064 2688 37072 2752
rect 37136 2688 37152 2752
rect 37216 2688 37232 2752
rect 37296 2688 37312 2752
rect 37376 2688 37384 2752
rect 37064 2128 37384 2688
rect 44288 7648 44608 7664
rect 44288 7584 44296 7648
rect 44360 7584 44376 7648
rect 44440 7584 44456 7648
rect 44520 7584 44536 7648
rect 44600 7584 44608 7648
rect 44288 6560 44608 7584
rect 44288 6496 44296 6560
rect 44360 6496 44376 6560
rect 44440 6496 44456 6560
rect 44520 6496 44536 6560
rect 44600 6496 44608 6560
rect 44288 5472 44608 6496
rect 44288 5408 44296 5472
rect 44360 5408 44376 5472
rect 44440 5408 44456 5472
rect 44520 5408 44536 5472
rect 44600 5408 44608 5472
rect 44288 4384 44608 5408
rect 44288 4320 44296 4384
rect 44360 4320 44376 4384
rect 44440 4320 44456 4384
rect 44520 4320 44536 4384
rect 44600 4320 44608 4384
rect 44288 3296 44608 4320
rect 44288 3232 44296 3296
rect 44360 3232 44376 3296
rect 44440 3232 44456 3296
rect 44520 3232 44536 3296
rect 44600 3232 44608 3296
rect 44288 2208 44608 3232
rect 44288 2144 44296 2208
rect 44360 2144 44376 2208
rect 44440 2144 44456 2208
rect 44520 2144 44536 2208
rect 44600 2144 44608 2208
rect 44288 2128 44608 2144
rect 51512 7104 51832 7664
rect 51512 7040 51520 7104
rect 51584 7040 51600 7104
rect 51664 7040 51680 7104
rect 51744 7040 51760 7104
rect 51824 7040 51832 7104
rect 51512 6016 51832 7040
rect 51512 5952 51520 6016
rect 51584 5952 51600 6016
rect 51664 5952 51680 6016
rect 51744 5952 51760 6016
rect 51824 5952 51832 6016
rect 51512 4928 51832 5952
rect 51512 4864 51520 4928
rect 51584 4864 51600 4928
rect 51664 4864 51680 4928
rect 51744 4864 51760 4928
rect 51824 4864 51832 4928
rect 51512 3840 51832 4864
rect 51512 3776 51520 3840
rect 51584 3776 51600 3840
rect 51664 3776 51680 3840
rect 51744 3776 51760 3840
rect 51824 3776 51832 3840
rect 51512 2752 51832 3776
rect 51512 2688 51520 2752
rect 51584 2688 51600 2752
rect 51664 2688 51680 2752
rect 51744 2688 51760 2752
rect 51824 2688 51832 2752
rect 51512 2128 51832 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 31096 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__B
timestamp 1649977179
transform -1 0 30544 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A0
timestamp 1649977179
transform -1 0 38272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A0
timestamp 1649977179
transform -1 0 41952 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A1
timestamp 1649977179
transform 1 0 39192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1649977179
transform -1 0 35512 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__B
timestamp 1649977179
transform 1 0 38916 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A0
timestamp 1649977179
transform 1 0 46920 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A1
timestamp 1649977179
transform 1 0 46920 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__S
timestamp 1649977179
transform -1 0 44528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A0
timestamp 1649977179
transform 1 0 55292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A1
timestamp 1649977179
transform -1 0 58052 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__S
timestamp 1649977179
transform -1 0 56488 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A_N
timestamp 1649977179
transform 1 0 49496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__B
timestamp 1649977179
transform 1 0 48116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__C
timestamp 1649977179
transform 1 0 47012 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A0
timestamp 1649977179
transform 1 0 57132 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A1
timestamp 1649977179
transform -1 0 56856 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__S
timestamp 1649977179
transform -1 0 55936 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A_N
timestamp 1649977179
transform -1 0 26588 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__B
timestamp 1649977179
transform -1 0 24564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__C
timestamp 1649977179
transform 1 0 24564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A1
timestamp 1649977179
transform -1 0 34224 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A
timestamp 1649977179
transform -1 0 57408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__B_N
timestamp 1649977179
transform -1 0 56028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1649977179
transform 1 0 29716 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1649977179
transform 1 0 43056 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__B
timestamp 1649977179
transform 1 0 38180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__B
timestamp 1649977179
transform 1 0 35696 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__C_N
timestamp 1649977179
transform -1 0 34684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__B1
timestamp 1649977179
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1649977179
transform -1 0 46092 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__B
timestamp 1649977179
transform -1 0 45724 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__B
timestamp 1649977179
transform 1 0 31280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__C
timestamp 1649977179
transform -1 0 30544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__B1
timestamp 1649977179
transform 1 0 32568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__B
timestamp 1649977179
transform -1 0 32752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__164__A
timestamp 1649977179
transform -1 0 33396 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__166__A
timestamp 1649977179
transform -1 0 56304 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__168__A
timestamp 1649977179
transform -1 0 50692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__A
timestamp 1649977179
transform -1 0 50048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__B
timestamp 1649977179
transform -1 0 54832 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__C
timestamp 1649977179
transform 1 0 55016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A
timestamp 1649977179
transform -1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A2
timestamp 1649977179
transform 1 0 22724 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A1
timestamp 1649977179
transform 1 0 22816 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__C1
timestamp 1649977179
transform 1 0 4692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__A1
timestamp 1649977179
transform 1 0 22172 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__210__C1
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1649977179
transform -1 0 21620 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__212__A
timestamp 1649977179
transform -1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A0
timestamp 1649977179
transform -1 0 2116 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__A
timestamp 1649977179
transform 1 0 3128 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A0
timestamp 1649977179
transform -1 0 20240 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__219__A
timestamp 1649977179
transform -1 0 20792 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__221__A0
timestamp 1649977179
transform -1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A
timestamp 1649977179
transform -1 0 10580 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__A
timestamp 1649977179
transform 1 0 42504 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__225__A
timestamp 1649977179
transform 1 0 40480 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A
timestamp 1649977179
transform -1 0 34224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__227__A
timestamp 1649977179
transform -1 0 41952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A
timestamp 1649977179
transform -1 0 52900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__229__A
timestamp 1649977179
transform -1 0 51980 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__A
timestamp 1649977179
transform 1 0 38364 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A
timestamp 1649977179
transform 1 0 49496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__237__A
timestamp 1649977179
transform -1 0 28060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__CLK
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__239__CLK
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__CLK
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__241__CLK
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__CLK
timestamp 1649977179
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__243__CLK
timestamp 1649977179
transform 1 0 23828 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__CLK
timestamp 1649977179
transform 1 0 20608 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__CLK
timestamp 1649977179
transform 1 0 25116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__246__CLK
timestamp 1649977179
transform 1 0 6440 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__CLK
timestamp 1649977179
transform 1 0 21160 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__248__CLK
timestamp 1649977179
transform -1 0 10120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__250__CLK
timestamp 1649977179
transform 1 0 33764 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__CLK
timestamp 1649977179
transform 1 0 26312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__252__CLK
timestamp 1649977179
transform -1 0 33580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__CLK
timestamp 1649977179
transform -1 0 52256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__254__CLK
timestamp 1649977179
transform -1 0 53820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__CLK
timestamp 1649977179
transform -1 0 49680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__256__CLK
timestamp 1649977179
transform 1 0 47564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__CLK
timestamp 1649977179
transform 1 0 40388 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__258__CLK
timestamp 1649977179
transform 1 0 41676 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__CLK
timestamp 1649977179
transform 1 0 35604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__260__CLK
timestamp 1649977179
transform 1 0 46460 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__CLK
timestamp 1649977179
transform 1 0 25668 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__264__GATE_N
timestamp 1649977179
transform -1 0 52256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__D
timestamp 1649977179
transform 1 0 36616 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__GATE_N
timestamp 1649977179
transform -1 0 35236 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__GATE_N
timestamp 1649977179
transform 1 0 41584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_wb_clk_i_A
timestamp 1649977179
transform -1 0 28980 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 3036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 7268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 2208 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 14444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 15916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 8832 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 7176 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 1932 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 2668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 7820 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 6532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output19_A
timestamp 1649977179
transform -1 0 23460 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output20_A
timestamp 1649977179
transform -1 0 23552 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output24_A
timestamp 1649977179
transform -1 0 22448 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output25_A
timestamp 1649977179
transform -1 0 23368 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output26_A
timestamp 1649977179
transform -1 0 19412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output27_A
timestamp 1649977179
transform 1 0 36616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output30_A
timestamp 1649977179
transform -1 0 25852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_A
timestamp 1649977179
transform -1 0 27876 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output32_A
timestamp 1649977179
transform -1 0 7176 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater36_A
timestamp 1649977179
transform -1 0 51244 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10
timestamp 1649977179
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40
timestamp 1649977179
transform 1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6808 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68
timestamp 1649977179
transform 1 0 7360 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79
timestamp 1649977179
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_122
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1649977179
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143
timestamp 1649977179
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_178
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_199
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_213
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_220
timestamp 1649977179
transform 1 0 21344 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_232
timestamp 1649977179
transform 1 0 22448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1649977179
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_248
timestamp 1649977179
transform 1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1649977179
transform 1 0 26220 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_279
timestamp 1649977179
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_297
timestamp 1649977179
transform 1 0 28428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_313
timestamp 1649977179
transform 1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1649977179
transform 1 0 30544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_324
timestamp 1649977179
transform 1 0 30912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_328
timestamp 1649977179
transform 1 0 31280 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_340
timestamp 1649977179
transform 1 0 32384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1649977179
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_354
timestamp 1649977179
transform 1 0 33672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_368
timestamp 1649977179
transform 1 0 34960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_382
timestamp 1649977179
transform 1 0 36248 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1649977179
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_396
timestamp 1649977179
transform 1 0 37536 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_410
timestamp 1649977179
transform 1 0 38824 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1649977179
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_424
timestamp 1649977179
transform 1 0 40112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_431
timestamp 1649977179
transform 1 0 40756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_438
timestamp 1649977179
transform 1 0 41400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1649977179
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_452
timestamp 1649977179
transform 1 0 42688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_459
timestamp 1649977179
transform 1 0 43332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_466
timestamp 1649977179
transform 1 0 43976 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1649977179
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_480
timestamp 1649977179
transform 1 0 45264 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_487
timestamp 1649977179
transform 1 0 45908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_494
timestamp 1649977179
transform 1 0 46552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1649977179
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_508
timestamp 1649977179
transform 1 0 47840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_515
timestamp 1649977179
transform 1 0 48484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_522
timestamp 1649977179
transform 1 0 49128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_528
timestamp 1649977179
transform 1 0 49680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_536
timestamp 1649977179
transform 1 0 50416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_543
timestamp 1649977179
transform 1 0 51060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_550
timestamp 1649977179
transform 1 0 51704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_556
timestamp 1649977179
transform 1 0 52256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_564
timestamp 1649977179
transform 1 0 52992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_571
timestamp 1649977179
transform 1 0 53636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_578
timestamp 1649977179
transform 1 0 54280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_584
timestamp 1649977179
transform 1 0 54832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_595
timestamp 1649977179
transform 1 0 55844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_602
timestamp 1649977179
transform 1 0 56488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_609
timestamp 1649977179
transform 1 0 57132 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_615
timestamp 1649977179
transform 1 0 57684 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_620
timestamp 1649977179
transform 1 0 58144 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_624
timestamp 1649977179
transform 1 0 58512 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1649977179
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1649977179
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_28
timestamp 1649977179
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_65
timestamp 1649977179
transform 1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_74
timestamp 1649977179
transform 1 0 7912 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_84
timestamp 1649977179
transform 1 0 8832 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_90
timestamp 1649977179
transform 1 0 9384 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_94
timestamp 1649977179
transform 1 0 9752 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_101
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1649977179
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_122
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_136
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_174
timestamp 1649977179
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_188
timestamp 1649977179
transform 1 0 18400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1649977179
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_215
timestamp 1649977179
transform 1 0 20884 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_230
timestamp 1649977179
transform 1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_238
timestamp 1649977179
transform 1 0 23000 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_262
timestamp 1649977179
transform 1 0 25208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_270
timestamp 1649977179
transform 1 0 25944 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_275
timestamp 1649977179
transform 1 0 26404 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_285
timestamp 1649977179
transform 1 0 27324 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_291
timestamp 1649977179
transform 1 0 27876 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1649977179
transform 1 0 28244 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_319
timestamp 1649977179
transform 1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_340
timestamp 1649977179
transform 1 0 32384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_347
timestamp 1649977179
transform 1 0 33028 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_373
timestamp 1649977179
transform 1 0 35420 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_380
timestamp 1649977179
transform 1 0 36064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1649977179
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1649977179
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_396
timestamp 1649977179
transform 1 0 37536 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1649977179
transform 1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_410
timestamp 1649977179
transform 1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_417
timestamp 1649977179
transform 1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_424
timestamp 1649977179
transform 1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_431
timestamp 1649977179
transform 1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_438
timestamp 1649977179
transform 1 0 41400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1649977179
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_452
timestamp 1649977179
transform 1 0 42688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_459
timestamp 1649977179
transform 1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_466
timestamp 1649977179
transform 1 0 43976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_473
timestamp 1649977179
transform 1 0 44620 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_480
timestamp 1649977179
transform 1 0 45264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_487
timestamp 1649977179
transform 1 0 45908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_494
timestamp 1649977179
transform 1 0 46552 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_500
timestamp 1649977179
transform 1 0 47104 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_508
timestamp 1649977179
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_515
timestamp 1649977179
transform 1 0 48484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_522
timestamp 1649977179
transform 1 0 49128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_528
timestamp 1649977179
transform 1 0 49680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_537
timestamp 1649977179
transform 1 0 50508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_544
timestamp 1649977179
transform 1 0 51152 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_551
timestamp 1649977179
transform 1 0 51796 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1649977179
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_564
timestamp 1649977179
transform 1 0 52992 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_571
timestamp 1649977179
transform 1 0 53636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_589
timestamp 1649977179
transform 1 0 55292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_602
timestamp 1649977179
transform 1 0 56488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_609
timestamp 1649977179
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_615
timestamp 1649977179
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_620
timestamp 1649977179
transform 1 0 58144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_624
timestamp 1649977179
transform 1 0 58512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_5
timestamp 1649977179
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1649977179
transform 1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_38
timestamp 1649977179
transform 1 0 4600 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_44
timestamp 1649977179
transform 1 0 5152 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1649977179
transform 1 0 5520 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1649977179
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_66
timestamp 1649977179
transform 1 0 7176 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_73
timestamp 1649977179
transform 1 0 7820 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_88
timestamp 1649977179
transform 1 0 9200 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_96
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_100
timestamp 1649977179
transform 1 0 10304 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_105
timestamp 1649977179
transform 1 0 10764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_112
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_125
timestamp 1649977179
transform 1 0 12604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1649977179
transform 1 0 14812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1649977179
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_171
timestamp 1649977179
transform 1 0 16836 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_182
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1649977179
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_210
timestamp 1649977179
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1649977179
transform 1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_227
timestamp 1649977179
transform 1 0 21988 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_235
timestamp 1649977179
transform 1 0 22724 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_240
timestamp 1649977179
transform 1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1649977179
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_264
timestamp 1649977179
transform 1 0 25392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_272
timestamp 1649977179
transform 1 0 26128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_280
timestamp 1649977179
transform 1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1649977179
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_312
timestamp 1649977179
transform 1 0 29808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_325
timestamp 1649977179
transform 1 0 31004 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_332
timestamp 1649977179
transform 1 0 31648 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_336
timestamp 1649977179
transform 1 0 32016 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_340
timestamp 1649977179
transform 1 0 32384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_347
timestamp 1649977179
transform 1 0 33028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_354
timestamp 1649977179
transform 1 0 33672 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1649977179
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_368
timestamp 1649977179
transform 1 0 34960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_374
timestamp 1649977179
transform 1 0 35512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_387
timestamp 1649977179
transform 1 0 36708 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_394
timestamp 1649977179
transform 1 0 37352 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_416
timestamp 1649977179
transform 1 0 39376 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_424
timestamp 1649977179
transform 1 0 40112 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_431
timestamp 1649977179
transform 1 0 40756 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_438
timestamp 1649977179
transform 1 0 41400 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_454
timestamp 1649977179
transform 1 0 42872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_461
timestamp 1649977179
transform 1 0 43516 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_468
timestamp 1649977179
transform 1 0 44160 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_486
timestamp 1649977179
transform 1 0 45816 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_501
timestamp 1649977179
transform 1 0 47196 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_525
timestamp 1649977179
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_531
timestamp 1649977179
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_545
timestamp 1649977179
transform 1 0 51244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_552
timestamp 1649977179
transform 1 0 51888 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_577
timestamp 1649977179
transform 1 0 54188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_584
timestamp 1649977179
transform 1 0 54832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_598
timestamp 1649977179
transform 1 0 56120 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_605
timestamp 1649977179
transform 1 0 56764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_612
timestamp 1649977179
transform 1 0 57408 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_619
timestamp 1649977179
transform 1 0 58052 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp 1649977179
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_12
timestamp 1649977179
transform 1 0 2208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_20
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1649977179
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_76
timestamp 1649977179
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_96
timestamp 1649977179
transform 1 0 9936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_102
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_121
timestamp 1649977179
transform 1 0 12236 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_127
timestamp 1649977179
transform 1 0 12788 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_134
timestamp 1649977179
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_141
timestamp 1649977179
transform 1 0 14076 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_148
timestamp 1649977179
transform 1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp 1649977179
transform 1 0 15364 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1649977179
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_178
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1649977179
transform 1 0 18400 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_212
timestamp 1649977179
transform 1 0 20608 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_216
timestamp 1649977179
transform 1 0 20976 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_233
timestamp 1649977179
transform 1 0 22540 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_245
timestamp 1649977179
transform 1 0 23644 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_266
timestamp 1649977179
transform 1 0 25576 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_272
timestamp 1649977179
transform 1 0 26128 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_276
timestamp 1649977179
transform 1 0 26496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_284
timestamp 1649977179
transform 1 0 27232 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_290
timestamp 1649977179
transform 1 0 27784 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_294
timestamp 1649977179
transform 1 0 28152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_318
timestamp 1649977179
transform 1 0 30360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_325
timestamp 1649977179
transform 1 0 31004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_331
timestamp 1649977179
transform 1 0 31556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_345
timestamp 1649977179
transform 1 0 32844 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_371
timestamp 1649977179
transform 1 0 35236 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_381
timestamp 1649977179
transform 1 0 36156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1649977179
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_399
timestamp 1649977179
transform 1 0 37812 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_406
timestamp 1649977179
transform 1 0 38456 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_412
timestamp 1649977179
transform 1 0 39008 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_416
timestamp 1649977179
transform 1 0 39376 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_442
timestamp 1649977179
transform 1 0 41768 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_449
timestamp 1649977179
transform 1 0 42412 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_453
timestamp 1649977179
transform 1 0 42780 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_458
timestamp 1649977179
transform 1 0 43240 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_467
timestamp 1649977179
transform 1 0 44068 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_474
timestamp 1649977179
transform 1 0 44712 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_481
timestamp 1649977179
transform 1 0 45356 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_488
timestamp 1649977179
transform 1 0 46000 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1649977179
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1649977179
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_525
timestamp 1649977179
transform 1 0 49404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_532
timestamp 1649977179
transform 1 0 50048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_539
timestamp 1649977179
transform 1 0 50692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_546
timestamp 1649977179
transform 1 0 51336 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1649977179
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1649977179
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_582
timestamp 1649977179
transform 1 0 54648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_588
timestamp 1649977179
transform 1 0 55200 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_605
timestamp 1649977179
transform 1 0 56764 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_611
timestamp 1649977179
transform 1 0 57316 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1649977179
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_619
timestamp 1649977179
transform 1 0 58052 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_19
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_52
timestamp 1649977179
transform 1 0 5888 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_60
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_66
timestamp 1649977179
transform 1 0 7176 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_73
timestamp 1649977179
transform 1 0 7820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_90
timestamp 1649977179
transform 1 0 9384 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1649977179
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_127
timestamp 1649977179
transform 1 0 12788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_136
timestamp 1649977179
transform 1 0 13616 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 1649977179
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_155
timestamp 1649977179
transform 1 0 15364 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_162
timestamp 1649977179
transform 1 0 16008 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_173
timestamp 1649977179
transform 1 0 17020 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_181
timestamp 1649977179
transform 1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1649977179
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_213
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_223
timestamp 1649977179
transform 1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_227
timestamp 1649977179
transform 1 0 21988 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_236
timestamp 1649977179
transform 1 0 22816 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1649977179
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_261
timestamp 1649977179
transform 1 0 25116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_296
timestamp 1649977179
transform 1 0 28336 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_300
timestamp 1649977179
transform 1 0 28704 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_304
timestamp 1649977179
transform 1 0 29072 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_316
timestamp 1649977179
transform 1 0 30176 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_338
timestamp 1649977179
transform 1 0 32200 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_344
timestamp 1649977179
transform 1 0 32752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1649977179
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_369
timestamp 1649977179
transform 1 0 35052 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_390
timestamp 1649977179
transform 1 0 36984 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_396
timestamp 1649977179
transform 1 0 37536 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_407
timestamp 1649977179
transform 1 0 38548 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1649977179
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1649977179
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_424
timestamp 1649977179
transform 1 0 40112 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_430
timestamp 1649977179
transform 1 0 40664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_454
timestamp 1649977179
transform 1 0 42872 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_4_463
timestamp 1649977179
transform 1 0 43700 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_472
timestamp 1649977179
transform 1 0 44528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_480
timestamp 1649977179
transform 1 0 45264 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_509
timestamp 1649977179
transform 1 0 47932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_515
timestamp 1649977179
transform 1 0 48484 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_528
timestamp 1649977179
transform 1 0 49680 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_536
timestamp 1649977179
transform 1 0 50416 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_542
timestamp 1649977179
transform 1 0 50968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_546
timestamp 1649977179
transform 1 0 51336 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_4_566
timestamp 1649977179
transform 1 0 53176 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_584
timestamp 1649977179
transform 1 0 54832 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_594
timestamp 1649977179
transform 1 0 55752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_600
timestamp 1649977179
transform 1 0 56304 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_606
timestamp 1649977179
transform 1 0 56856 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_612
timestamp 1649977179
transform 1 0 57408 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_624
timestamp 1649977179
transform 1 0 58512 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_21
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_24
timestamp 1649977179
transform 1 0 3312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_40
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1649977179
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_59
timestamp 1649977179
transform 1 0 6532 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_66
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_73
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_80
timestamp 1649977179
transform 1 0 8464 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_87
timestamp 1649977179
transform 1 0 9108 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1649977179
transform 1 0 9752 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_101
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1649977179
transform 1 0 11960 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_135
timestamp 1649977179
transform 1 0 13524 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_139
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_143
timestamp 1649977179
transform 1 0 14260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_150
timestamp 1649977179
transform 1 0 14904 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_157
timestamp 1649977179
transform 1 0 15548 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_171
timestamp 1649977179
transform 1 0 16836 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_178
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_188
timestamp 1649977179
transform 1 0 18400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_196
timestamp 1649977179
transform 1 0 19136 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_204
timestamp 1649977179
transform 1 0 19872 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_208
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_214
timestamp 1649977179
transform 1 0 20792 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_231
timestamp 1649977179
transform 1 0 22356 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_243
timestamp 1649977179
transform 1 0 23460 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_255
timestamp 1649977179
transform 1 0 24564 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_262
timestamp 1649977179
transform 1 0 25208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_269
timestamp 1649977179
transform 1 0 25852 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1649977179
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_297
timestamp 1649977179
transform 1 0 28428 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_304
timestamp 1649977179
transform 1 0 29072 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_312
timestamp 1649977179
transform 1 0 29808 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_323
timestamp 1649977179
transform 1 0 30820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_327
timestamp 1649977179
transform 1 0 31188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_330
timestamp 1649977179
transform 1 0 31464 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_340
timestamp 1649977179
transform 1 0 32384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_362
timestamp 1649977179
transform 1 0 34408 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_372
timestamp 1649977179
transform 1 0 35328 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_376
timestamp 1649977179
transform 1 0 35696 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_382
timestamp 1649977179
transform 1 0 36248 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1649977179
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_398
timestamp 1649977179
transform 1 0 37720 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_404
timestamp 1649977179
transform 1 0 38272 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_412
timestamp 1649977179
transform 1 0 39008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_418
timestamp 1649977179
transform 1 0 39560 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_429
timestamp 1649977179
transform 1 0 40572 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_433
timestamp 1649977179
transform 1 0 40940 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_437
timestamp 1649977179
transform 1 0 41308 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_443
timestamp 1649977179
transform 1 0 41860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1649977179
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_456
timestamp 1649977179
transform 1 0 43056 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_463
timestamp 1649977179
transform 1 0 43700 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_471
timestamp 1649977179
transform 1 0 44436 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_475
timestamp 1649977179
transform 1 0 44804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_485
timestamp 1649977179
transform 1 0 45724 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_493
timestamp 1649977179
transform 1 0 46460 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1649977179
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_508
timestamp 1649977179
transform 1 0 47840 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_512
timestamp 1649977179
transform 1 0 48208 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_518
timestamp 1649977179
transform 1 0 48760 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_525
timestamp 1649977179
transform 1 0 49404 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_532
timestamp 1649977179
transform 1 0 50048 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_538
timestamp 1649977179
transform 1 0 50600 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_542
timestamp 1649977179
transform 1 0 50968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_549
timestamp 1649977179
transform 1 0 51612 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_556
timestamp 1649977179
transform 1 0 52256 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_564
timestamp 1649977179
transform 1 0 52992 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_571
timestamp 1649977179
transform 1 0 53636 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_578
timestamp 1649977179
transform 1 0 54280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_586
timestamp 1649977179
transform 1 0 55016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_590
timestamp 1649977179
transform 1 0 55384 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_596
timestamp 1649977179
transform 1 0 55936 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_602
timestamp 1649977179
transform 1 0 56488 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_614
timestamp 1649977179
transform 1 0 57592 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1649977179
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_49
timestamp 1649977179
transform 1 0 5612 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_54
timestamp 1649977179
transform 1 0 6072 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_60
timestamp 1649977179
transform 1 0 6624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_64
timestamp 1649977179
transform 1 0 6992 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_67
timestamp 1649977179
transform 1 0 7268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_73
timestamp 1649977179
transform 1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 1649977179
transform 1 0 9292 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1649977179
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_101
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_110
timestamp 1649977179
transform 1 0 11224 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_118
timestamp 1649977179
transform 1 0 11960 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_122
timestamp 1649977179
transform 1 0 12328 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_131
timestamp 1649977179
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_145
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_152
timestamp 1649977179
transform 1 0 15088 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_158
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_161
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_168
timestamp 1649977179
transform 1 0 16560 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_172
timestamp 1649977179
transform 1 0 16928 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_176
timestamp 1649977179
transform 1 0 17296 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_188
timestamp 1649977179
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_205
timestamp 1649977179
transform 1 0 19964 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_208
timestamp 1649977179
transform 1 0 20240 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_214
timestamp 1649977179
transform 1 0 20792 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_223
timestamp 1649977179
transform 1 0 21620 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_229
timestamp 1649977179
transform 1 0 22172 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_232
timestamp 1649977179
transform 1 0 22448 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_238
timestamp 1649977179
transform 1 0 23000 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_244
timestamp 1649977179
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_257
timestamp 1649977179
transform 1 0 24748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_263
timestamp 1649977179
transform 1 0 25300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_269
timestamp 1649977179
transform 1 0 25852 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_276
timestamp 1649977179
transform 1 0 26496 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_283
timestamp 1649977179
transform 1 0 27140 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_290
timestamp 1649977179
transform 1 0 27784 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_297
timestamp 1649977179
transform 1 0 28428 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1649977179
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_313
timestamp 1649977179
transform 1 0 29900 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_317
timestamp 1649977179
transform 1 0 30268 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_320
timestamp 1649977179
transform 1 0 30544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_328
timestamp 1649977179
transform 1 0 31280 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_338
timestamp 1649977179
transform 1 0 32200 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_344
timestamp 1649977179
transform 1 0 32752 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_350
timestamp 1649977179
transform 1 0 33304 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_355
timestamp 1649977179
transform 1 0 33764 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_372
timestamp 1649977179
transform 1 0 35328 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_378
timestamp 1649977179
transform 1 0 35880 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_385
timestamp 1649977179
transform 1 0 36524 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_391
timestamp 1649977179
transform 1 0 37076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_399
timestamp 1649977179
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_405
timestamp 1649977179
transform 1 0 38364 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_417
timestamp 1649977179
transform 1 0 39468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_423
timestamp 1649977179
transform 1 0 40020 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_429
timestamp 1649977179
transform 1 0 40572 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_437
timestamp 1649977179
transform 1 0 41308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_442
timestamp 1649977179
transform 1 0 41768 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_452
timestamp 1649977179
transform 1 0 42688 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_458
timestamp 1649977179
transform 1 0 43240 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_470
timestamp 1649977179
transform 1 0 44344 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_477
timestamp 1649977179
transform 1 0 44988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_483
timestamp 1649977179
transform 1 0 45540 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_489
timestamp 1649977179
transform 1 0 46092 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_495
timestamp 1649977179
transform 1 0 46644 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_501
timestamp 1649977179
transform 1 0 47196 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_507
timestamp 1649977179
transform 1 0 47748 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1649977179
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_525
timestamp 1649977179
transform 1 0 49404 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_528
timestamp 1649977179
transform 1 0 49680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_533
timestamp 1649977179
transform 1 0 50140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_538
timestamp 1649977179
transform 1 0 50600 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_545
timestamp 1649977179
transform 1 0 51244 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_549
timestamp 1649977179
transform 1 0 51612 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_553
timestamp 1649977179
transform 1 0 51980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_560
timestamp 1649977179
transform 1 0 52624 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_567
timestamp 1649977179
transform 1 0 53268 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_573
timestamp 1649977179
transform 1 0 53820 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_585
timestamp 1649977179
transform 1 0 54924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_591
timestamp 1649977179
transform 1 0 55476 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_597
timestamp 1649977179
transform 1 0 56028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_609
timestamp 1649977179
transform 1 0 57132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_621
timestamp 1649977179
transform 1 0 58236 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_78
timestamp 1649977179
transform 1 0 8280 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_84
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_90
timestamp 1649977179
transform 1 0 9384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_96
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_100
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_103
timestamp 1649977179
transform 1 0 10580 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_119
timestamp 1649977179
transform 1 0 12052 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_131
timestamp 1649977179
transform 1 0 13156 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_143
timestamp 1649977179
transform 1 0 14260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_155
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_211
timestamp 1649977179
transform 1 0 20516 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_214
timestamp 1649977179
transform 1 0 20792 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_220
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_242
timestamp 1649977179
transform 1 0 23368 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_254
timestamp 1649977179
transform 1 0 24472 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_266
timestamp 1649977179
transform 1 0 25576 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_269
timestamp 1649977179
transform 1 0 25852 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1649977179
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_283
timestamp 1649977179
transform 1 0 27140 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_320
timestamp 1649977179
transform 1 0 30544 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_326
timestamp 1649977179
transform 1 0 31096 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_334
timestamp 1649977179
transform 1 0 31832 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_351
timestamp 1649977179
transform 1 0 33396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_357
timestamp 1649977179
transform 1 0 33948 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_365
timestamp 1649977179
transform 1 0 34684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_371
timestamp 1649977179
transform 1 0 35236 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_377
timestamp 1649977179
transform 1 0 35788 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_389
timestamp 1649977179
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1649977179
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1649977179
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1649977179
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1649977179
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1649977179
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1649977179
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_473
timestamp 1649977179
transform 1 0 44620 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_481
timestamp 1649977179
transform 1 0 45356 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1649977179
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1649977179
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1649977179
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1649977179
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_517
timestamp 1649977179
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_529
timestamp 1649977179
transform 1 0 49772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_532
timestamp 1649977179
transform 1 0 50048 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_536
timestamp 1649977179
transform 1 0 50416 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_539
timestamp 1649977179
transform 1 0 50692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_545
timestamp 1649977179
transform 1 0 51244 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_553
timestamp 1649977179
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_559
timestamp 1649977179
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_563
timestamp 1649977179
transform 1 0 52900 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_575
timestamp 1649977179
transform 1 0 54004 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_587
timestamp 1649977179
transform 1 0 55108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_599
timestamp 1649977179
transform 1 0 56212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_611
timestamp 1649977179
transform 1 0 57316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1649977179
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_617
timestamp 1649977179
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_60
timestamp 1649977179
transform 1 0 6624 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_72
timestamp 1649977179
transform 1 0 7728 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1649977179
transform 1 0 9660 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_98
timestamp 1649977179
transform 1 0 10120 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_110
timestamp 1649977179
transform 1 0 11224 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_115
timestamp 1649977179
transform 1 0 11684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_127
timestamp 1649977179
transform 1 0 12788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_145
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_157
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_169
timestamp 1649977179
transform 1 0 16652 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_175
timestamp 1649977179
transform 1 0 17204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_187
timestamp 1649977179
transform 1 0 18308 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_220
timestamp 1649977179
transform 1 0 21344 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_232
timestamp 1649977179
transform 1 0 22448 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_244
timestamp 1649977179
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_256
timestamp 1649977179
transform 1 0 24656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_268
timestamp 1649977179
transform 1 0 25760 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1649977179
transform 1 0 26312 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_281
timestamp 1649977179
transform 1 0 26956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_285
timestamp 1649977179
transform 1 0 27324 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_291
timestamp 1649977179
transform 1 0 27876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_303
timestamp 1649977179
transform 1 0 28980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_8_353
timestamp 1649977179
transform 1 0 33580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1649977179
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_381
timestamp 1649977179
transform 1 0 36156 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_385
timestamp 1649977179
transform 1 0 36524 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_397
timestamp 1649977179
transform 1 0 37628 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_409
timestamp 1649977179
transform 1 0 38732 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_417
timestamp 1649977179
transform 1 0 39468 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_424
timestamp 1649977179
transform 1 0 40112 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_436
timestamp 1649977179
transform 1 0 41216 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_448
timestamp 1649977179
transform 1 0 42320 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_460
timestamp 1649977179
transform 1 0 43424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_465
timestamp 1649977179
transform 1 0 43884 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_473
timestamp 1649977179
transform 1 0 44620 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1649977179
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_489
timestamp 1649977179
transform 1 0 46092 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_495
timestamp 1649977179
transform 1 0 46644 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_507
timestamp 1649977179
transform 1 0 47748 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_519
timestamp 1649977179
transform 1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_525
timestamp 1649977179
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1649977179
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_533
timestamp 1649977179
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_545
timestamp 1649977179
transform 1 0 51244 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_553
timestamp 1649977179
transform 1 0 51980 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_556
timestamp 1649977179
transform 1 0 52256 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_568
timestamp 1649977179
transform 1 0 53360 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_576
timestamp 1649977179
transform 1 0 54096 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_580
timestamp 1649977179
transform 1 0 54464 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_589
timestamp 1649977179
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_601
timestamp 1649977179
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_613
timestamp 1649977179
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_29
timestamp 1649977179
transform 1 0 3772 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_38
timestamp 1649977179
transform 1 0 4600 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_45
timestamp 1649977179
transform 1 0 5244 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_52
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_66
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_73
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_80
timestamp 1649977179
transform 1 0 8464 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_85
timestamp 1649977179
transform 1 0 8924 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_90
timestamp 1649977179
transform 1 0 9384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_94
timestamp 1649977179
transform 1 0 9752 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_98
timestamp 1649977179
transform 1 0 10120 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_120
timestamp 1649977179
transform 1 0 12144 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_124
timestamp 1649977179
transform 1 0 12512 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_128
timestamp 1649977179
transform 1 0 12880 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_135
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_139
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_141
timestamp 1649977179
transform 1 0 14076 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_150
timestamp 1649977179
transform 1 0 14904 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_157
timestamp 1649977179
transform 1 0 15548 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_178
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_185
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_192
timestamp 1649977179
transform 1 0 18768 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_197
timestamp 1649977179
transform 1 0 19228 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_203
timestamp 1649977179
transform 1 0 19780 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_210
timestamp 1649977179
transform 1 0 20424 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_216
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_229
timestamp 1649977179
transform 1 0 22172 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_233
timestamp 1649977179
transform 1 0 22540 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_240
timestamp 1649977179
transform 1 0 23184 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_244
timestamp 1649977179
transform 1 0 23552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_248
timestamp 1649977179
transform 1 0 23920 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_253
timestamp 1649977179
transform 1 0 24380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_262
timestamp 1649977179
transform 1 0 25208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_269
timestamp 1649977179
transform 1 0 25852 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1649977179
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_290
timestamp 1649977179
transform 1 0 27784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_297
timestamp 1649977179
transform 1 0 28428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_304
timestamp 1649977179
transform 1 0 29072 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_309
timestamp 1649977179
transform 1 0 29532 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_315
timestamp 1649977179
transform 1 0 30084 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_319
timestamp 1649977179
transform 1 0 30452 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_323
timestamp 1649977179
transform 1 0 30820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_330
timestamp 1649977179
transform 1 0 31464 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_340
timestamp 1649977179
transform 1 0 32384 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_347
timestamp 1649977179
transform 1 0 33028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_351
timestamp 1649977179
transform 1 0 33396 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_355
timestamp 1649977179
transform 1 0 33764 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_363
timestamp 1649977179
transform 1 0 34500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_368
timestamp 1649977179
transform 1 0 34960 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_375
timestamp 1649977179
transform 1 0 35604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_382
timestamp 1649977179
transform 1 0 36248 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_390
timestamp 1649977179
transform 1 0 36984 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_396
timestamp 1649977179
transform 1 0 37536 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1649977179
transform 1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_410
timestamp 1649977179
transform 1 0 38824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_418
timestamp 1649977179
transform 1 0 39560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_424
timestamp 1649977179
transform 1 0 40112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_431
timestamp 1649977179
transform 1 0 40756 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_438
timestamp 1649977179
transform 1 0 41400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_446
timestamp 1649977179
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_452
timestamp 1649977179
transform 1 0 42688 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_459
timestamp 1649977179
transform 1 0 43332 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_466
timestamp 1649977179
transform 1 0 43976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_474
timestamp 1649977179
transform 1 0 44712 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_480
timestamp 1649977179
transform 1 0 45264 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_487
timestamp 1649977179
transform 1 0 45908 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_494
timestamp 1649977179
transform 1 0 46552 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_502
timestamp 1649977179
transform 1 0 47288 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_508
timestamp 1649977179
transform 1 0 47840 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_515
timestamp 1649977179
transform 1 0 48484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_522
timestamp 1649977179
transform 1 0 49128 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_530
timestamp 1649977179
transform 1 0 49864 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_536
timestamp 1649977179
transform 1 0 50416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_543
timestamp 1649977179
transform 1 0 51060 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_550
timestamp 1649977179
transform 1 0 51704 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_558
timestamp 1649977179
transform 1 0 52440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_564
timestamp 1649977179
transform 1 0 52992 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_571
timestamp 1649977179
transform 1 0 53636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_578
timestamp 1649977179
transform 1 0 54280 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_586
timestamp 1649977179
transform 1 0 55016 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_592
timestamp 1649977179
transform 1 0 55568 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_599
timestamp 1649977179
transform 1 0 56212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_606
timestamp 1649977179
transform 1 0 56856 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_614
timestamp 1649977179
transform 1 0 57592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_617
timestamp 1649977179
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_20 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_21
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1649977179
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1649977179
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1649977179
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1649977179
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1649977179
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1649977179
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1649977179
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1649977179
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 24288 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 34592 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 39744 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 44896 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 50048 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 55200 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__or3b_2  _117_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _118_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 36708 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _119_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 40112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _120_
timestamp 1649977179
transform -1 0 39376 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1649977179
transform -1 0 43516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _122_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 32476 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _123_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _124_
timestamp 1649977179
transform -1 0 45816 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform -1 0 46000 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _126_
timestamp 1649977179
transform 1 0 55660 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1649977179
transform 1 0 53360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _128_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 46552 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _129_
timestamp 1649977179
transform 1 0 55292 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1649977179
transform -1 0 51612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _131_
timestamp 1649977179
transform -1 0 31648 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1649977179
transform -1 0 31648 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _133_
timestamp 1649977179
transform -1 0 25208 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1649977179
transform -1 0 26496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _135_
timestamp 1649977179
transform -1 0 26220 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _136_
timestamp 1649977179
transform -1 0 31004 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1649977179
transform -1 0 31004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _138_
timestamp 1649977179
transform -1 0 25392 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1649977179
transform 1 0 24932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _140_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 55292 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1649977179
transform 1 0 57776 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _142_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 41308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _143_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 35788 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _144_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 30820 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_2  _145_
timestamp 1649977179
transform 1 0 42412 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _146_
timestamp 1649977179
transform 1 0 44252 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _147_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 39560 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _148_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37168 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _149_
timestamp 1649977179
transform -1 0 35328 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _150_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 39928 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _151_
timestamp 1649977179
transform -1 0 45540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _152_
timestamp 1649977179
transform 1 0 46552 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1649977179
transform -1 0 49404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _154_
timestamp 1649977179
transform -1 0 44804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _155_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12328 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_1  _156_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30912 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _157_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 32200 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _158_
timestamp 1649977179
transform 1 0 43424 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _159_
timestamp 1649977179
transform 1 0 36248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _160_
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _161_
timestamp 1649977179
transform 1 0 33396 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _162_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 34776 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _163_
timestamp 1649977179
transform -1 0 45724 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _164_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 33212 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1649977179
transform 1 0 27508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _166_
timestamp 1649977179
transform 1 0 55292 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1649977179
transform -1 0 55384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _168_
timestamp 1649977179
transform 1 0 50692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 51336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _170_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 48300 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1649977179
transform -1 0 50416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _172_
timestamp 1649977179
transform 1 0 50048 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _173_
timestamp 1649977179
transform 1 0 57132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _174_
timestamp 1649977179
transform 1 0 33948 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1649977179
transform 1 0 35788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _176_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4692 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _177_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12696 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1649977179
transform -1 0 13340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _179_
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _180_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16192 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _181_
timestamp 1649977179
transform -1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _182_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14352 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1649977179
transform -1 0 18400 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _185_
timestamp 1649977179
transform -1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 1649977179
transform -1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _187_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp 1649977179
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1649977179
transform 1 0 9568 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _190_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23920 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _191_
timestamp 1649977179
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _192_
timestamp 1649977179
transform 1 0 18768 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _193_
timestamp 1649977179
transform 1 0 17848 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _194_
timestamp 1649977179
transform 1 0 22080 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _195_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5888 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _196_
timestamp 1649977179
transform -1 0 17756 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _197_
timestamp 1649977179
transform 1 0 18216 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _198_
timestamp 1649977179
transform -1 0 25116 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _199_
timestamp 1649977179
transform 1 0 5060 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _200_
timestamp 1649977179
transform -1 0 6624 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _201_
timestamp 1649977179
transform -1 0 12788 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _202_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_2  _203_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _204_
timestamp 1649977179
transform -1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _205_
timestamp 1649977179
transform -1 0 13432 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _206_
timestamp 1649977179
transform 1 0 2576 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _207_
timestamp 1649977179
transform 1 0 4876 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _208_
timestamp 1649977179
transform 1 0 15732 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _209_
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _210_
timestamp 1649977179
transform -1 0 22540 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _211_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21620 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _212_
timestamp 1649977179
transform -1 0 10764 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _213_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _214_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _215_
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _216_
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1649977179
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1649977179
transform -1 0 20424 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _219_
timestamp 1649977179
transform -1 0 21252 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _220_
timestamp 1649977179
transform -1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _221_
timestamp 1649977179
transform 1 0 11776 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _222_
timestamp 1649977179
transform -1 0 11040 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _224_
timestamp 1649977179
transform 1 0 42872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 1649977179
transform -1 0 40112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _226_
timestamp 1649977179
transform -1 0 32384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _227_
timestamp 1649977179
transform -1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _228_
timestamp 1649977179
transform 1 0 52716 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _229_
timestamp 1649977179
transform 1 0 51980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _230_
timestamp 1649977179
transform 1 0 37628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1649977179
transform 1 0 46552 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _232_
timestamp 1649977179
transform 1 0 43792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _233_
timestamp 1649977179
transform 1 0 39100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _234_
timestamp 1649977179
transform -1 0 45264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _235_
timestamp 1649977179
transform -1 0 37720 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _236_
timestamp 1649977179
transform 1 0 49772 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1649977179
transform -1 0 28336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _238_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 30728 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _239_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _240_
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _241_
timestamp 1649977179
transform 1 0 10396 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _242_
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _243_
timestamp 1649977179
transform 1 0 24104 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _244_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18768 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _245_
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _246_
timestamp 1649977179
transform 1 0 4140 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _247_
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _248_
timestamp 1649977179
transform -1 0 9936 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtp_1  _249_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 55292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dfrtp_1  _250_
timestamp 1649977179
transform 1 0 33396 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _251_
timestamp 1649977179
transform 1 0 27232 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _252_
timestamp 1649977179
transform 1 0 33580 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _253_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 52256 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _254_
timestamp 1649977179
transform 1 0 52716 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _255_
timestamp 1649977179
transform -1 0 49404 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _256_
timestamp 1649977179
transform -1 0 49404 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _257_
timestamp 1649977179
transform -1 0 41768 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _258_
timestamp 1649977179
transform -1 0 42872 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _259_
timestamp 1649977179
transform 1 0 35144 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _260_
timestamp 1649977179
transform 1 0 46000 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _261_
timestamp 1649977179
transform 1 0 25852 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtn_2  _262_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 55568 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _263_ dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 53728 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _264_
timestamp 1649977179
transform -1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _265_
timestamp 1649977179
transform -1 0 34224 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _266_
timestamp 1649977179
transform -1 0 53176 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _267_
timestamp 1649977179
transform -1 0 42872 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _268_
timestamp 1649977179
transform -1 0 49680 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 28520 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1649977179
transform -1 0 25208 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1649977179
transform 1 0 28612 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 14720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 4140 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 9752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 3680 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 5520 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 7176 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1649977179
transform -1 0 23644 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1649977179
transform -1 0 23184 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1649977179
transform -1 0 22264 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1649977179
transform -1 0 23000 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1649977179
transform -1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1649977179
transform -1 0 22448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1649977179
transform -1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1649977179
transform 1 0 23552 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1649977179
transform -1 0 29900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1649977179
transform -1 0 26128 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1649977179
transform 1 0 26036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1649977179
transform -1 0 26864 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1649977179
transform -1 0 27324 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1649977179
transform -1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1649977179
transform -1 0 8832 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1649977179
transform -1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater36
timestamp 1649977179
transform 1 0 51060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_37 dependencies/pdks/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4600 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_38
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_39
timestamp 1649977179
transform 1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_40
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_41
timestamp 1649977179
transform -1 0 10120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_42
timestamp 1649977179
transform -1 0 11684 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_43
timestamp 1649977179
transform -1 0 12880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_44
timestamp 1649977179
transform -1 0 14444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_45
timestamp 1649977179
transform 1 0 15272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_46
timestamp 1649977179
transform -1 0 17204 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_47
timestamp 1649977179
transform 1 0 17848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_48
timestamp 1649977179
transform -1 0 19780 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_49
timestamp 1649977179
transform -1 0 21344 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_50
timestamp 1649977179
transform -1 0 22540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_51
timestamp 1649977179
transform -1 0 23920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_52
timestamp 1649977179
transform 1 0 24932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_53
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_54
timestamp 1649977179
transform 1 0 27508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_55
timestamp 1649977179
transform 1 0 28796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_56
timestamp 1649977179
transform -1 0 30820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_57
timestamp 1649977179
transform -1 0 32384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_58
timestamp 1649977179
transform -1 0 33764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_59
timestamp 1649977179
transform -1 0 35604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_60
timestamp 1649977179
transform -1 0 36524 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_61
timestamp 1649977179
transform -1 0 38180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_62
timestamp 1649977179
transform -1 0 40112 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_63
timestamp 1649977179
transform -1 0 40756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_64
timestamp 1649977179
transform -1 0 42688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_65
timestamp 1649977179
transform -1 0 43976 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_66
timestamp 1649977179
transform -1 0 45264 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_67
timestamp 1649977179
transform -1 0 46552 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_68
timestamp 1649977179
transform -1 0 47840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_69
timestamp 1649977179
transform -1 0 49128 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_70
timestamp 1649977179
transform -1 0 50416 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_71
timestamp 1649977179
transform -1 0 51704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_72
timestamp 1649977179
transform -1 0 53636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_73
timestamp 1649977179
transform -1 0 54464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_74
timestamp 1649977179
transform -1 0 56212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_75
timestamp 1649977179
transform -1 0 5244 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_76
timestamp 1649977179
transform -1 0 6624 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_77
timestamp 1649977179
transform -1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_78
timestamp 1649977179
transform -1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_79
timestamp 1649977179
transform -1 0 10764 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_80
timestamp 1649977179
transform -1 0 12144 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_81
timestamp 1649977179
transform -1 0 13524 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_82
timestamp 1649977179
transform -1 0 14904 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_83
timestamp 1649977179
transform -1 0 16192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_84
timestamp 1649977179
transform -1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_85
timestamp 1649977179
transform 1 0 18492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_86
timestamp 1649977179
transform -1 0 20424 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_87
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_88
timestamp 1649977179
transform -1 0 23184 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_89
timestamp 1649977179
transform -1 0 24656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_90
timestamp 1649977179
transform -1 0 25852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_91
timestamp 1649977179
transform -1 0 27324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_92
timestamp 1649977179
transform 1 0 28152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_93
timestamp 1649977179
transform -1 0 30084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_94
timestamp 1649977179
transform -1 0 31464 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_95
timestamp 1649977179
transform -1 0 33028 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_96
timestamp 1649977179
transform -1 0 34960 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_97
timestamp 1649977179
transform -1 0 36248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_98
timestamp 1649977179
transform -1 0 37536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_99
timestamp 1649977179
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_100
timestamp 1649977179
transform -1 0 40112 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_101
timestamp 1649977179
transform -1 0 41400 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_102
timestamp 1649977179
transform -1 0 43332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_103
timestamp 1649977179
transform -1 0 43884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_104
timestamp 1649977179
transform -1 0 45908 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_105
timestamp 1649977179
transform -1 0 46644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_106
timestamp 1649977179
transform -1 0 48484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_107
timestamp 1649977179
transform -1 0 49404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_108
timestamp 1649977179
transform -1 0 51060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_109
timestamp 1649977179
transform -1 0 52992 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_110
timestamp 1649977179
transform -1 0 54280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_111
timestamp 1649977179
transform -1 0 55568 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_112
timestamp 1649977179
transform -1 0 56856 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_113
timestamp 1649977179
transform -1 0 57132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_114
timestamp 1649977179
transform -1 0 58144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_115
timestamp 1649977179
transform -1 0 54280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_116
timestamp 1649977179
transform -1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_117
timestamp 1649977179
transform 1 0 16744 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_118
timestamp 1649977179
transform 1 0 15272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_119
timestamp 1649977179
transform 1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_120
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_121
timestamp 1649977179
transform 1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_122
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_123
timestamp 1649977179
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_124
timestamp 1649977179
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_125
timestamp 1649977179
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_126
timestamp 1649977179
transform -1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_127
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_128
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_129
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_130
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_131
timestamp 1649977179
transform -1 0 21620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_132
timestamp 1649977179
transform 1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_133
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_134
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_135
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_136
timestamp 1649977179
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_137
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_138
timestamp 1649977179
transform -1 0 27140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_139
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_140
timestamp 1649977179
transform -1 0 28428 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_141
timestamp 1649977179
transform 1 0 26220 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_142
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_143
timestamp 1649977179
transform 1 0 25576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_144
timestamp 1649977179
transform -1 0 29072 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_145
timestamp 1649977179
transform -1 0 29072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_146
timestamp 1649977179
transform -1 0 29808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_147
timestamp 1649977179
transform -1 0 30544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_148
timestamp 1649977179
transform 1 0 27968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_149
timestamp 1649977179
transform 1 0 27876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_150
timestamp 1649977179
transform -1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_151
timestamp 1649977179
transform 1 0 28796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_152
timestamp 1649977179
transform -1 0 32384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_153
timestamp 1649977179
transform -1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_154
timestamp 1649977179
transform -1 0 33028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_155
timestamp 1649977179
transform -1 0 33028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_156
timestamp 1649977179
transform -1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_157
timestamp 1649977179
transform -1 0 33672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_158
timestamp 1649977179
transform -1 0 35604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_159
timestamp 1649977179
transform -1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_160
timestamp 1649977179
transform -1 0 36248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_161
timestamp 1649977179
transform -1 0 33672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_162
timestamp 1649977179
transform -1 0 36708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_163
timestamp 1649977179
transform -1 0 37536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_164
timestamp 1649977179
transform -1 0 34960 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_165
timestamp 1649977179
transform -1 0 36064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_166
timestamp 1649977179
transform -1 0 38180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_167
timestamp 1649977179
transform -1 0 37536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_168
timestamp 1649977179
transform -1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_169
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_170
timestamp 1649977179
transform -1 0 36800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_171
timestamp 1649977179
transform -1 0 40112 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_172
timestamp 1649977179
transform -1 0 37352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_173
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_174
timestamp 1649977179
transform -1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_175
timestamp 1649977179
transform -1 0 37996 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_176
timestamp 1649977179
transform -1 0 40756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_177
timestamp 1649977179
transform -1 0 38456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_178
timestamp 1649977179
transform -1 0 41400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_179
timestamp 1649977179
transform -1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_180
timestamp 1649977179
transform -1 0 42688 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_181
timestamp 1649977179
transform -1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_182
timestamp 1649977179
transform -1 0 40756 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_183
timestamp 1649977179
transform -1 0 42688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_184
timestamp 1649977179
transform -1 0 41400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_185
timestamp 1649977179
transform -1 0 43332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_186
timestamp 1649977179
transform -1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_187
timestamp 1649977179
transform -1 0 43976 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_188
timestamp 1649977179
transform -1 0 43976 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_189
timestamp 1649977179
transform -1 0 45264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_190
timestamp 1649977179
transform -1 0 44620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_191
timestamp 1649977179
transform -1 0 45908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_192
timestamp 1649977179
transform -1 0 45264 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_193
timestamp 1649977179
transform -1 0 46552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_194
timestamp 1649977179
transform -1 0 44160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_195
timestamp 1649977179
transform -1 0 45908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_196
timestamp 1649977179
transform -1 0 47840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_197
timestamp 1649977179
transform -1 0 46552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_198
timestamp 1649977179
transform -1 0 43700 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_199
timestamp 1649977179
transform -1 0 44712 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_200
timestamp 1649977179
transform -1 0 47840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_201
timestamp 1649977179
transform -1 0 45356 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_202
timestamp 1649977179
transform -1 0 48484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_203
timestamp 1649977179
transform -1 0 49128 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_204
timestamp 1649977179
transform -1 0 48484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_205
timestamp 1649977179
transform -1 0 51060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_206
timestamp 1649977179
transform -1 0 49128 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_207
timestamp 1649977179
transform -1 0 50416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_208
timestamp 1649977179
transform -1 0 51152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_209
timestamp 1649977179
transform -1 0 51704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_210
timestamp 1649977179
transform -1 0 47840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_211
timestamp 1649977179
transform -1 0 52992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_212
timestamp 1649977179
transform -1 0 51796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_213
timestamp 1649977179
transform -1 0 52992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_214
timestamp 1649977179
transform -1 0 50692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_215
timestamp 1649977179
transform -1 0 51888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_216
timestamp 1649977179
transform -1 0 53636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_217
timestamp 1649977179
transform -1 0 53636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_218
timestamp 1649977179
transform -1 0 54832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_219
timestamp 1649977179
transform -1 0 50048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_220
timestamp 1649977179
transform -1 0 56488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_221
timestamp 1649977179
transform -1 0 54280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_222
timestamp 1649977179
transform -1 0 51980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_223
timestamp 1649977179
transform -1 0 50600 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_224
timestamp 1649977179
transform -1 0 51244 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_225
timestamp 1649977179
transform -1 0 57132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_226
timestamp 1649977179
transform -1 0 56764 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_227
timestamp 1649977179
transform -1 0 58144 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_228
timestamp 1649977179
transform -1 0 51980 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_229
timestamp 1649977179
transform -1 0 52624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_230
timestamp 1649977179
transform -1 0 53268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_231
timestamp 1649977179
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_232
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_233
timestamp 1649977179
transform 1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_234
timestamp 1649977179
transform -1 0 10396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_235
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_236
timestamp 1649977179
transform 1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_237
timestamp 1649977179
transform -1 0 11224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_238
timestamp 1649977179
transform 1 0 4508 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_239
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_240
timestamp 1649977179
transform 1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_241
timestamp 1649977179
transform -1 0 12328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_242
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_243
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_244
timestamp 1649977179
transform -1 0 13156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_245
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_246
timestamp 1649977179
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_247
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_248
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_249
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_250
timestamp 1649977179
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_251
timestamp 1649977179
transform -1 0 15088 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_252
timestamp 1649977179
transform 1 0 14628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_253
timestamp 1649977179
transform 1 0 10120 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_254
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_255
timestamp 1649977179
transform 1 0 13800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_256
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_257
timestamp 1649977179
transform 1 0 14444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_258
timestamp 1649977179
transform 1 0 15088 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rlbp_macro_259
timestamp 1649977179
transform -1 0 17296 0 1 5440
box -38 -48 314 592
<< labels >>
flabel metal2 s 3974 9200 4030 10000 0 FreeSans 224 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 17774 9200 17830 10000 0 FreeSans 224 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 19154 9200 19210 10000 0 FreeSans 224 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 20534 9200 20590 10000 0 FreeSans 224 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 21914 9200 21970 10000 0 FreeSans 224 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal2 s 23294 9200 23350 10000 0 FreeSans 224 90 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 24674 9200 24730 10000 0 FreeSans 224 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 26054 9200 26110 10000 0 FreeSans 224 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 27434 9200 27490 10000 0 FreeSans 224 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 28814 9200 28870 10000 0 FreeSans 224 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 30194 9200 30250 10000 0 FreeSans 224 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal2 s 5354 9200 5410 10000 0 FreeSans 224 90 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 31574 9200 31630 10000 0 FreeSans 224 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 32954 9200 33010 10000 0 FreeSans 224 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 34334 9200 34390 10000 0 FreeSans 224 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 35714 9200 35770 10000 0 FreeSans 224 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal2 s 37094 9200 37150 10000 0 FreeSans 224 90 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 38474 9200 38530 10000 0 FreeSans 224 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal2 s 39854 9200 39910 10000 0 FreeSans 224 90 0 0 io_in[26]
port 18 nsew signal input
flabel metal2 s 41234 9200 41290 10000 0 FreeSans 224 90 0 0 io_in[27]
port 19 nsew signal input
flabel metal2 s 42614 9200 42670 10000 0 FreeSans 224 90 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 43994 9200 44050 10000 0 FreeSans 224 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 6734 9200 6790 10000 0 FreeSans 224 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal2 s 45374 9200 45430 10000 0 FreeSans 224 90 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 46754 9200 46810 10000 0 FreeSans 224 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 48134 9200 48190 10000 0 FreeSans 224 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 49514 9200 49570 10000 0 FreeSans 224 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 50894 9200 50950 10000 0 FreeSans 224 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal2 s 52274 9200 52330 10000 0 FreeSans 224 90 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 53654 9200 53710 10000 0 FreeSans 224 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal2 s 55034 9200 55090 10000 0 FreeSans 224 90 0 0 io_in[37]
port 30 nsew signal input
flabel metal2 s 8114 9200 8170 10000 0 FreeSans 224 90 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 9494 9200 9550 10000 0 FreeSans 224 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 10874 9200 10930 10000 0 FreeSans 224 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 12254 9200 12310 10000 0 FreeSans 224 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 13634 9200 13690 10000 0 FreeSans 224 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 15014 9200 15070 10000 0 FreeSans 224 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal2 s 16394 9200 16450 10000 0 FreeSans 224 90 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 4434 9200 4490 10000 0 FreeSans 224 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal2 s 18234 9200 18290 10000 0 FreeSans 224 90 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal2 s 19614 9200 19670 10000 0 FreeSans 224 90 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal2 s 20994 9200 21050 10000 0 FreeSans 224 90 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal2 s 22374 9200 22430 10000 0 FreeSans 224 90 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal2 s 23754 9200 23810 10000 0 FreeSans 224 90 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 25134 9200 25190 10000 0 FreeSans 224 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 26514 9200 26570 10000 0 FreeSans 224 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 27894 9200 27950 10000 0 FreeSans 224 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 29274 9200 29330 10000 0 FreeSans 224 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 30654 9200 30710 10000 0 FreeSans 224 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 5814 9200 5870 10000 0 FreeSans 224 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 32034 9200 32090 10000 0 FreeSans 224 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 33414 9200 33470 10000 0 FreeSans 224 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 34794 9200 34850 10000 0 FreeSans 224 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 36174 9200 36230 10000 0 FreeSans 224 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal2 s 37554 9200 37610 10000 0 FreeSans 224 90 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 38934 9200 38990 10000 0 FreeSans 224 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 40314 9200 40370 10000 0 FreeSans 224 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal2 s 41694 9200 41750 10000 0 FreeSans 224 90 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal2 s 43074 9200 43130 10000 0 FreeSans 224 90 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal2 s 44454 9200 44510 10000 0 FreeSans 224 90 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 7194 9200 7250 10000 0 FreeSans 224 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 45834 9200 45890 10000 0 FreeSans 224 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal2 s 47214 9200 47270 10000 0 FreeSans 224 90 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal2 s 48594 9200 48650 10000 0 FreeSans 224 90 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal2 s 49974 9200 50030 10000 0 FreeSans 224 90 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal2 s 51354 9200 51410 10000 0 FreeSans 224 90 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal2 s 52734 9200 52790 10000 0 FreeSans 224 90 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 54114 9200 54170 10000 0 FreeSans 224 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal2 s 55494 9200 55550 10000 0 FreeSans 224 90 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal2 s 8574 9200 8630 10000 0 FreeSans 224 90 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 9954 9200 10010 10000 0 FreeSans 224 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal2 s 11334 9200 11390 10000 0 FreeSans 224 90 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal2 s 12714 9200 12770 10000 0 FreeSans 224 90 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal2 s 14094 9200 14150 10000 0 FreeSans 224 90 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal2 s 15474 9200 15530 10000 0 FreeSans 224 90 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 16854 9200 16910 10000 0 FreeSans 224 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal2 s 4894 9200 4950 10000 0 FreeSans 224 90 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal2 s 18694 9200 18750 10000 0 FreeSans 224 90 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal2 s 20074 9200 20130 10000 0 FreeSans 224 90 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal2 s 21454 9200 21510 10000 0 FreeSans 224 90 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal2 s 22834 9200 22890 10000 0 FreeSans 224 90 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 24214 9200 24270 10000 0 FreeSans 224 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 25594 9200 25650 10000 0 FreeSans 224 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 26974 9200 27030 10000 0 FreeSans 224 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 28354 9200 28410 10000 0 FreeSans 224 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 29734 9200 29790 10000 0 FreeSans 224 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 31114 9200 31170 10000 0 FreeSans 224 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 6274 9200 6330 10000 0 FreeSans 224 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 32494 9200 32550 10000 0 FreeSans 224 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 33874 9200 33930 10000 0 FreeSans 224 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 35254 9200 35310 10000 0 FreeSans 224 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 36634 9200 36690 10000 0 FreeSans 224 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal2 s 38014 9200 38070 10000 0 FreeSans 224 90 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 39394 9200 39450 10000 0 FreeSans 224 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 40774 9200 40830 10000 0 FreeSans 224 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 42154 9200 42210 10000 0 FreeSans 224 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 43534 9200 43590 10000 0 FreeSans 224 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 44914 9200 44970 10000 0 FreeSans 224 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal2 s 7654 9200 7710 10000 0 FreeSans 224 90 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal2 s 46294 9200 46350 10000 0 FreeSans 224 90 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal2 s 47674 9200 47730 10000 0 FreeSans 224 90 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 49054 9200 49110 10000 0 FreeSans 224 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 50434 9200 50490 10000 0 FreeSans 224 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal2 s 51814 9200 51870 10000 0 FreeSans 224 90 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal2 s 53194 9200 53250 10000 0 FreeSans 224 90 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 54574 9200 54630 10000 0 FreeSans 224 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 55954 9200 56010 10000 0 FreeSans 224 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 9034 9200 9090 10000 0 FreeSans 224 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 10414 9200 10470 10000 0 FreeSans 224 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 11794 9200 11850 10000 0 FreeSans 224 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 13174 9200 13230 10000 0 FreeSans 224 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal2 s 14554 9200 14610 10000 0 FreeSans 224 90 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal2 s 15934 9200 15990 10000 0 FreeSans 224 90 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal2 s 17314 9200 17370 10000 0 FreeSans 224 90 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 52366 0 52422 800 0 FreeSans 224 90 0 0 irq[0]
port 114 nsew signal tristate
flabel metal2 s 52458 0 52514 800 0 FreeSans 224 90 0 0 irq[1]
port 115 nsew signal tristate
flabel metal2 s 52550 0 52606 800 0 FreeSans 224 90 0 0 irq[2]
port 116 nsew signal tristate
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 la_data_in[0]
port 117 nsew signal input
flabel metal2 s 44638 0 44694 800 0 FreeSans 224 90 0 0 la_data_in[100]
port 118 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 la_data_in[101]
port 119 nsew signal input
flabel metal2 s 45190 0 45246 800 0 FreeSans 224 90 0 0 la_data_in[102]
port 120 nsew signal input
flabel metal2 s 45466 0 45522 800 0 FreeSans 224 90 0 0 la_data_in[103]
port 121 nsew signal input
flabel metal2 s 45742 0 45798 800 0 FreeSans 224 90 0 0 la_data_in[104]
port 122 nsew signal input
flabel metal2 s 46018 0 46074 800 0 FreeSans 224 90 0 0 la_data_in[105]
port 123 nsew signal input
flabel metal2 s 46294 0 46350 800 0 FreeSans 224 90 0 0 la_data_in[106]
port 124 nsew signal input
flabel metal2 s 46570 0 46626 800 0 FreeSans 224 90 0 0 la_data_in[107]
port 125 nsew signal input
flabel metal2 s 46846 0 46902 800 0 FreeSans 224 90 0 0 la_data_in[108]
port 126 nsew signal input
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 la_data_in[109]
port 127 nsew signal input
flabel metal2 s 19798 0 19854 800 0 FreeSans 224 90 0 0 la_data_in[10]
port 128 nsew signal input
flabel metal2 s 47398 0 47454 800 0 FreeSans 224 90 0 0 la_data_in[110]
port 129 nsew signal input
flabel metal2 s 47674 0 47730 800 0 FreeSans 224 90 0 0 la_data_in[111]
port 130 nsew signal input
flabel metal2 s 47950 0 48006 800 0 FreeSans 224 90 0 0 la_data_in[112]
port 131 nsew signal input
flabel metal2 s 48226 0 48282 800 0 FreeSans 224 90 0 0 la_data_in[113]
port 132 nsew signal input
flabel metal2 s 48502 0 48558 800 0 FreeSans 224 90 0 0 la_data_in[114]
port 133 nsew signal input
flabel metal2 s 48778 0 48834 800 0 FreeSans 224 90 0 0 la_data_in[115]
port 134 nsew signal input
flabel metal2 s 49054 0 49110 800 0 FreeSans 224 90 0 0 la_data_in[116]
port 135 nsew signal input
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 la_data_in[117]
port 136 nsew signal input
flabel metal2 s 49606 0 49662 800 0 FreeSans 224 90 0 0 la_data_in[118]
port 137 nsew signal input
flabel metal2 s 49882 0 49938 800 0 FreeSans 224 90 0 0 la_data_in[119]
port 138 nsew signal input
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 la_data_in[11]
port 139 nsew signal input
flabel metal2 s 50158 0 50214 800 0 FreeSans 224 90 0 0 la_data_in[120]
port 140 nsew signal input
flabel metal2 s 50434 0 50490 800 0 FreeSans 224 90 0 0 la_data_in[121]
port 141 nsew signal input
flabel metal2 s 50710 0 50766 800 0 FreeSans 224 90 0 0 la_data_in[122]
port 142 nsew signal input
flabel metal2 s 50986 0 51042 800 0 FreeSans 224 90 0 0 la_data_in[123]
port 143 nsew signal input
flabel metal2 s 51262 0 51318 800 0 FreeSans 224 90 0 0 la_data_in[124]
port 144 nsew signal input
flabel metal2 s 51538 0 51594 800 0 FreeSans 224 90 0 0 la_data_in[125]
port 145 nsew signal input
flabel metal2 s 51814 0 51870 800 0 FreeSans 224 90 0 0 la_data_in[126]
port 146 nsew signal input
flabel metal2 s 52090 0 52146 800 0 FreeSans 224 90 0 0 la_data_in[127]
port 147 nsew signal input
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 la_data_in[12]
port 148 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 la_data_in[13]
port 149 nsew signal input
flabel metal2 s 20902 0 20958 800 0 FreeSans 224 90 0 0 la_data_in[14]
port 150 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 la_data_in[15]
port 151 nsew signal input
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 la_data_in[16]
port 152 nsew signal input
flabel metal2 s 21730 0 21786 800 0 FreeSans 224 90 0 0 la_data_in[17]
port 153 nsew signal input
flabel metal2 s 22006 0 22062 800 0 FreeSans 224 90 0 0 la_data_in[18]
port 154 nsew signal input
flabel metal2 s 22282 0 22338 800 0 FreeSans 224 90 0 0 la_data_in[19]
port 155 nsew signal input
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 la_data_in[1]
port 156 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 la_data_in[20]
port 157 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 la_data_in[21]
port 158 nsew signal input
flabel metal2 s 23110 0 23166 800 0 FreeSans 224 90 0 0 la_data_in[22]
port 159 nsew signal input
flabel metal2 s 23386 0 23442 800 0 FreeSans 224 90 0 0 la_data_in[23]
port 160 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 la_data_in[24]
port 161 nsew signal input
flabel metal2 s 23938 0 23994 800 0 FreeSans 224 90 0 0 la_data_in[25]
port 162 nsew signal input
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 la_data_in[26]
port 163 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 la_data_in[27]
port 164 nsew signal input
flabel metal2 s 24766 0 24822 800 0 FreeSans 224 90 0 0 la_data_in[28]
port 165 nsew signal input
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 la_data_in[29]
port 166 nsew signal input
flabel metal2 s 17590 0 17646 800 0 FreeSans 224 90 0 0 la_data_in[2]
port 167 nsew signal input
flabel metal2 s 25318 0 25374 800 0 FreeSans 224 90 0 0 la_data_in[30]
port 168 nsew signal input
flabel metal2 s 25594 0 25650 800 0 FreeSans 224 90 0 0 la_data_in[31]
port 169 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 la_data_in[32]
port 170 nsew signal input
flabel metal2 s 26146 0 26202 800 0 FreeSans 224 90 0 0 la_data_in[33]
port 171 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 la_data_in[34]
port 172 nsew signal input
flabel metal2 s 26698 0 26754 800 0 FreeSans 224 90 0 0 la_data_in[35]
port 173 nsew signal input
flabel metal2 s 26974 0 27030 800 0 FreeSans 224 90 0 0 la_data_in[36]
port 174 nsew signal input
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 la_data_in[37]
port 175 nsew signal input
flabel metal2 s 27526 0 27582 800 0 FreeSans 224 90 0 0 la_data_in[38]
port 176 nsew signal input
flabel metal2 s 27802 0 27858 800 0 FreeSans 224 90 0 0 la_data_in[39]
port 177 nsew signal input
flabel metal2 s 17866 0 17922 800 0 FreeSans 224 90 0 0 la_data_in[3]
port 178 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 la_data_in[40]
port 179 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 la_data_in[41]
port 180 nsew signal input
flabel metal2 s 28630 0 28686 800 0 FreeSans 224 90 0 0 la_data_in[42]
port 181 nsew signal input
flabel metal2 s 28906 0 28962 800 0 FreeSans 224 90 0 0 la_data_in[43]
port 182 nsew signal input
flabel metal2 s 29182 0 29238 800 0 FreeSans 224 90 0 0 la_data_in[44]
port 183 nsew signal input
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 la_data_in[45]
port 184 nsew signal input
flabel metal2 s 29734 0 29790 800 0 FreeSans 224 90 0 0 la_data_in[46]
port 185 nsew signal input
flabel metal2 s 30010 0 30066 800 0 FreeSans 224 90 0 0 la_data_in[47]
port 186 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 la_data_in[48]
port 187 nsew signal input
flabel metal2 s 30562 0 30618 800 0 FreeSans 224 90 0 0 la_data_in[49]
port 188 nsew signal input
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 la_data_in[4]
port 189 nsew signal input
flabel metal2 s 30838 0 30894 800 0 FreeSans 224 90 0 0 la_data_in[50]
port 190 nsew signal input
flabel metal2 s 31114 0 31170 800 0 FreeSans 224 90 0 0 la_data_in[51]
port 191 nsew signal input
flabel metal2 s 31390 0 31446 800 0 FreeSans 224 90 0 0 la_data_in[52]
port 192 nsew signal input
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 la_data_in[53]
port 193 nsew signal input
flabel metal2 s 31942 0 31998 800 0 FreeSans 224 90 0 0 la_data_in[54]
port 194 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_data_in[55]
port 195 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 la_data_in[56]
port 196 nsew signal input
flabel metal2 s 32770 0 32826 800 0 FreeSans 224 90 0 0 la_data_in[57]
port 197 nsew signal input
flabel metal2 s 33046 0 33102 800 0 FreeSans 224 90 0 0 la_data_in[58]
port 198 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 la_data_in[59]
port 199 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 la_data_in[5]
port 200 nsew signal input
flabel metal2 s 33598 0 33654 800 0 FreeSans 224 90 0 0 la_data_in[60]
port 201 nsew signal input
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 la_data_in[61]
port 202 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 la_data_in[62]
port 203 nsew signal input
flabel metal2 s 34426 0 34482 800 0 FreeSans 224 90 0 0 la_data_in[63]
port 204 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 la_data_in[64]
port 205 nsew signal input
flabel metal2 s 34978 0 35034 800 0 FreeSans 224 90 0 0 la_data_in[65]
port 206 nsew signal input
flabel metal2 s 35254 0 35310 800 0 FreeSans 224 90 0 0 la_data_in[66]
port 207 nsew signal input
flabel metal2 s 35530 0 35586 800 0 FreeSans 224 90 0 0 la_data_in[67]
port 208 nsew signal input
flabel metal2 s 35806 0 35862 800 0 FreeSans 224 90 0 0 la_data_in[68]
port 209 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_data_in[69]
port 210 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_data_in[6]
port 211 nsew signal input
flabel metal2 s 36358 0 36414 800 0 FreeSans 224 90 0 0 la_data_in[70]
port 212 nsew signal input
flabel metal2 s 36634 0 36690 800 0 FreeSans 224 90 0 0 la_data_in[71]
port 213 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 la_data_in[72]
port 214 nsew signal input
flabel metal2 s 37186 0 37242 800 0 FreeSans 224 90 0 0 la_data_in[73]
port 215 nsew signal input
flabel metal2 s 37462 0 37518 800 0 FreeSans 224 90 0 0 la_data_in[74]
port 216 nsew signal input
flabel metal2 s 37738 0 37794 800 0 FreeSans 224 90 0 0 la_data_in[75]
port 217 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 la_data_in[76]
port 218 nsew signal input
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 la_data_in[77]
port 219 nsew signal input
flabel metal2 s 38566 0 38622 800 0 FreeSans 224 90 0 0 la_data_in[78]
port 220 nsew signal input
flabel metal2 s 38842 0 38898 800 0 FreeSans 224 90 0 0 la_data_in[79]
port 221 nsew signal input
flabel metal2 s 18970 0 19026 800 0 FreeSans 224 90 0 0 la_data_in[7]
port 222 nsew signal input
flabel metal2 s 39118 0 39174 800 0 FreeSans 224 90 0 0 la_data_in[80]
port 223 nsew signal input
flabel metal2 s 39394 0 39450 800 0 FreeSans 224 90 0 0 la_data_in[81]
port 224 nsew signal input
flabel metal2 s 39670 0 39726 800 0 FreeSans 224 90 0 0 la_data_in[82]
port 225 nsew signal input
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 la_data_in[83]
port 226 nsew signal input
flabel metal2 s 40222 0 40278 800 0 FreeSans 224 90 0 0 la_data_in[84]
port 227 nsew signal input
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 la_data_in[85]
port 228 nsew signal input
flabel metal2 s 40774 0 40830 800 0 FreeSans 224 90 0 0 la_data_in[86]
port 229 nsew signal input
flabel metal2 s 41050 0 41106 800 0 FreeSans 224 90 0 0 la_data_in[87]
port 230 nsew signal input
flabel metal2 s 41326 0 41382 800 0 FreeSans 224 90 0 0 la_data_in[88]
port 231 nsew signal input
flabel metal2 s 41602 0 41658 800 0 FreeSans 224 90 0 0 la_data_in[89]
port 232 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 la_data_in[8]
port 233 nsew signal input
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 la_data_in[90]
port 234 nsew signal input
flabel metal2 s 42154 0 42210 800 0 FreeSans 224 90 0 0 la_data_in[91]
port 235 nsew signal input
flabel metal2 s 42430 0 42486 800 0 FreeSans 224 90 0 0 la_data_in[92]
port 236 nsew signal input
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 la_data_in[93]
port 237 nsew signal input
flabel metal2 s 42982 0 43038 800 0 FreeSans 224 90 0 0 la_data_in[94]
port 238 nsew signal input
flabel metal2 s 43258 0 43314 800 0 FreeSans 224 90 0 0 la_data_in[95]
port 239 nsew signal input
flabel metal2 s 43534 0 43590 800 0 FreeSans 224 90 0 0 la_data_in[96]
port 240 nsew signal input
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 la_data_in[97]
port 241 nsew signal input
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 la_data_in[98]
port 242 nsew signal input
flabel metal2 s 44362 0 44418 800 0 FreeSans 224 90 0 0 la_data_in[99]
port 243 nsew signal input
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 la_data_in[9]
port 244 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 la_data_out[0]
port 245 nsew signal tristate
flabel metal2 s 44730 0 44786 800 0 FreeSans 224 90 0 0 la_data_out[100]
port 246 nsew signal tristate
flabel metal2 s 45006 0 45062 800 0 FreeSans 224 90 0 0 la_data_out[101]
port 247 nsew signal tristate
flabel metal2 s 45282 0 45338 800 0 FreeSans 224 90 0 0 la_data_out[102]
port 248 nsew signal tristate
flabel metal2 s 45558 0 45614 800 0 FreeSans 224 90 0 0 la_data_out[103]
port 249 nsew signal tristate
flabel metal2 s 45834 0 45890 800 0 FreeSans 224 90 0 0 la_data_out[104]
port 250 nsew signal tristate
flabel metal2 s 46110 0 46166 800 0 FreeSans 224 90 0 0 la_data_out[105]
port 251 nsew signal tristate
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 la_data_out[106]
port 252 nsew signal tristate
flabel metal2 s 46662 0 46718 800 0 FreeSans 224 90 0 0 la_data_out[107]
port 253 nsew signal tristate
flabel metal2 s 46938 0 46994 800 0 FreeSans 224 90 0 0 la_data_out[108]
port 254 nsew signal tristate
flabel metal2 s 47214 0 47270 800 0 FreeSans 224 90 0 0 la_data_out[109]
port 255 nsew signal tristate
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 la_data_out[10]
port 256 nsew signal tristate
flabel metal2 s 47490 0 47546 800 0 FreeSans 224 90 0 0 la_data_out[110]
port 257 nsew signal tristate
flabel metal2 s 47766 0 47822 800 0 FreeSans 224 90 0 0 la_data_out[111]
port 258 nsew signal tristate
flabel metal2 s 48042 0 48098 800 0 FreeSans 224 90 0 0 la_data_out[112]
port 259 nsew signal tristate
flabel metal2 s 48318 0 48374 800 0 FreeSans 224 90 0 0 la_data_out[113]
port 260 nsew signal tristate
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 la_data_out[114]
port 261 nsew signal tristate
flabel metal2 s 48870 0 48926 800 0 FreeSans 224 90 0 0 la_data_out[115]
port 262 nsew signal tristate
flabel metal2 s 49146 0 49202 800 0 FreeSans 224 90 0 0 la_data_out[116]
port 263 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 la_data_out[117]
port 264 nsew signal tristate
flabel metal2 s 49698 0 49754 800 0 FreeSans 224 90 0 0 la_data_out[118]
port 265 nsew signal tristate
flabel metal2 s 49974 0 50030 800 0 FreeSans 224 90 0 0 la_data_out[119]
port 266 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 la_data_out[11]
port 267 nsew signal tristate
flabel metal2 s 50250 0 50306 800 0 FreeSans 224 90 0 0 la_data_out[120]
port 268 nsew signal tristate
flabel metal2 s 50526 0 50582 800 0 FreeSans 224 90 0 0 la_data_out[121]
port 269 nsew signal tristate
flabel metal2 s 50802 0 50858 800 0 FreeSans 224 90 0 0 la_data_out[122]
port 270 nsew signal tristate
flabel metal2 s 51078 0 51134 800 0 FreeSans 224 90 0 0 la_data_out[123]
port 271 nsew signal tristate
flabel metal2 s 51354 0 51410 800 0 FreeSans 224 90 0 0 la_data_out[124]
port 272 nsew signal tristate
flabel metal2 s 51630 0 51686 800 0 FreeSans 224 90 0 0 la_data_out[125]
port 273 nsew signal tristate
flabel metal2 s 51906 0 51962 800 0 FreeSans 224 90 0 0 la_data_out[126]
port 274 nsew signal tristate
flabel metal2 s 52182 0 52238 800 0 FreeSans 224 90 0 0 la_data_out[127]
port 275 nsew signal tristate
flabel metal2 s 20442 0 20498 800 0 FreeSans 224 90 0 0 la_data_out[12]
port 276 nsew signal tristate
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 la_data_out[13]
port 277 nsew signal tristate
flabel metal2 s 20994 0 21050 800 0 FreeSans 224 90 0 0 la_data_out[14]
port 278 nsew signal tristate
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 la_data_out[15]
port 279 nsew signal tristate
flabel metal2 s 21546 0 21602 800 0 FreeSans 224 90 0 0 la_data_out[16]
port 280 nsew signal tristate
flabel metal2 s 21822 0 21878 800 0 FreeSans 224 90 0 0 la_data_out[17]
port 281 nsew signal tristate
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 la_data_out[18]
port 282 nsew signal tristate
flabel metal2 s 22374 0 22430 800 0 FreeSans 224 90 0 0 la_data_out[19]
port 283 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 la_data_out[1]
port 284 nsew signal tristate
flabel metal2 s 22650 0 22706 800 0 FreeSans 224 90 0 0 la_data_out[20]
port 285 nsew signal tristate
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 la_data_out[21]
port 286 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 la_data_out[22]
port 287 nsew signal tristate
flabel metal2 s 23478 0 23534 800 0 FreeSans 224 90 0 0 la_data_out[23]
port 288 nsew signal tristate
flabel metal2 s 23754 0 23810 800 0 FreeSans 224 90 0 0 la_data_out[24]
port 289 nsew signal tristate
flabel metal2 s 24030 0 24086 800 0 FreeSans 224 90 0 0 la_data_out[25]
port 290 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 la_data_out[26]
port 291 nsew signal tristate
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 la_data_out[27]
port 292 nsew signal tristate
flabel metal2 s 24858 0 24914 800 0 FreeSans 224 90 0 0 la_data_out[28]
port 293 nsew signal tristate
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 la_data_out[29]
port 294 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 la_data_out[2]
port 295 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 la_data_out[30]
port 296 nsew signal tristate
flabel metal2 s 25686 0 25742 800 0 FreeSans 224 90 0 0 la_data_out[31]
port 297 nsew signal tristate
flabel metal2 s 25962 0 26018 800 0 FreeSans 224 90 0 0 la_data_out[32]
port 298 nsew signal tristate
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 la_data_out[33]
port 299 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 la_data_out[34]
port 300 nsew signal tristate
flabel metal2 s 26790 0 26846 800 0 FreeSans 224 90 0 0 la_data_out[35]
port 301 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 la_data_out[36]
port 302 nsew signal tristate
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 la_data_out[37]
port 303 nsew signal tristate
flabel metal2 s 27618 0 27674 800 0 FreeSans 224 90 0 0 la_data_out[38]
port 304 nsew signal tristate
flabel metal2 s 27894 0 27950 800 0 FreeSans 224 90 0 0 la_data_out[39]
port 305 nsew signal tristate
flabel metal2 s 17958 0 18014 800 0 FreeSans 224 90 0 0 la_data_out[3]
port 306 nsew signal tristate
flabel metal2 s 28170 0 28226 800 0 FreeSans 224 90 0 0 la_data_out[40]
port 307 nsew signal tristate
flabel metal2 s 28446 0 28502 800 0 FreeSans 224 90 0 0 la_data_out[41]
port 308 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 la_data_out[42]
port 309 nsew signal tristate
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 la_data_out[43]
port 310 nsew signal tristate
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 la_data_out[44]
port 311 nsew signal tristate
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 la_data_out[45]
port 312 nsew signal tristate
flabel metal2 s 29826 0 29882 800 0 FreeSans 224 90 0 0 la_data_out[46]
port 313 nsew signal tristate
flabel metal2 s 30102 0 30158 800 0 FreeSans 224 90 0 0 la_data_out[47]
port 314 nsew signal tristate
flabel metal2 s 30378 0 30434 800 0 FreeSans 224 90 0 0 la_data_out[48]
port 315 nsew signal tristate
flabel metal2 s 30654 0 30710 800 0 FreeSans 224 90 0 0 la_data_out[49]
port 316 nsew signal tristate
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 la_data_out[4]
port 317 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_data_out[50]
port 318 nsew signal tristate
flabel metal2 s 31206 0 31262 800 0 FreeSans 224 90 0 0 la_data_out[51]
port 319 nsew signal tristate
flabel metal2 s 31482 0 31538 800 0 FreeSans 224 90 0 0 la_data_out[52]
port 320 nsew signal tristate
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 la_data_out[53]
port 321 nsew signal tristate
flabel metal2 s 32034 0 32090 800 0 FreeSans 224 90 0 0 la_data_out[54]
port 322 nsew signal tristate
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 la_data_out[55]
port 323 nsew signal tristate
flabel metal2 s 32586 0 32642 800 0 FreeSans 224 90 0 0 la_data_out[56]
port 324 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 la_data_out[57]
port 325 nsew signal tristate
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 la_data_out[58]
port 326 nsew signal tristate
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 la_data_out[59]
port 327 nsew signal tristate
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 la_data_out[5]
port 328 nsew signal tristate
flabel metal2 s 33690 0 33746 800 0 FreeSans 224 90 0 0 la_data_out[60]
port 329 nsew signal tristate
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 la_data_out[61]
port 330 nsew signal tristate
flabel metal2 s 34242 0 34298 800 0 FreeSans 224 90 0 0 la_data_out[62]
port 331 nsew signal tristate
flabel metal2 s 34518 0 34574 800 0 FreeSans 224 90 0 0 la_data_out[63]
port 332 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 la_data_out[64]
port 333 nsew signal tristate
flabel metal2 s 35070 0 35126 800 0 FreeSans 224 90 0 0 la_data_out[65]
port 334 nsew signal tristate
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 la_data_out[66]
port 335 nsew signal tristate
flabel metal2 s 35622 0 35678 800 0 FreeSans 224 90 0 0 la_data_out[67]
port 336 nsew signal tristate
flabel metal2 s 35898 0 35954 800 0 FreeSans 224 90 0 0 la_data_out[68]
port 337 nsew signal tristate
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 la_data_out[69]
port 338 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 la_data_out[6]
port 339 nsew signal tristate
flabel metal2 s 36450 0 36506 800 0 FreeSans 224 90 0 0 la_data_out[70]
port 340 nsew signal tristate
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 la_data_out[71]
port 341 nsew signal tristate
flabel metal2 s 37002 0 37058 800 0 FreeSans 224 90 0 0 la_data_out[72]
port 342 nsew signal tristate
flabel metal2 s 37278 0 37334 800 0 FreeSans 224 90 0 0 la_data_out[73]
port 343 nsew signal tristate
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 la_data_out[74]
port 344 nsew signal tristate
flabel metal2 s 37830 0 37886 800 0 FreeSans 224 90 0 0 la_data_out[75]
port 345 nsew signal tristate
flabel metal2 s 38106 0 38162 800 0 FreeSans 224 90 0 0 la_data_out[76]
port 346 nsew signal tristate
flabel metal2 s 38382 0 38438 800 0 FreeSans 224 90 0 0 la_data_out[77]
port 347 nsew signal tristate
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 la_data_out[78]
port 348 nsew signal tristate
flabel metal2 s 38934 0 38990 800 0 FreeSans 224 90 0 0 la_data_out[79]
port 349 nsew signal tristate
flabel metal2 s 19062 0 19118 800 0 FreeSans 224 90 0 0 la_data_out[7]
port 350 nsew signal tristate
flabel metal2 s 39210 0 39266 800 0 FreeSans 224 90 0 0 la_data_out[80]
port 351 nsew signal tristate
flabel metal2 s 39486 0 39542 800 0 FreeSans 224 90 0 0 la_data_out[81]
port 352 nsew signal tristate
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 la_data_out[82]
port 353 nsew signal tristate
flabel metal2 s 40038 0 40094 800 0 FreeSans 224 90 0 0 la_data_out[83]
port 354 nsew signal tristate
flabel metal2 s 40314 0 40370 800 0 FreeSans 224 90 0 0 la_data_out[84]
port 355 nsew signal tristate
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 la_data_out[85]
port 356 nsew signal tristate
flabel metal2 s 40866 0 40922 800 0 FreeSans 224 90 0 0 la_data_out[86]
port 357 nsew signal tristate
flabel metal2 s 41142 0 41198 800 0 FreeSans 224 90 0 0 la_data_out[87]
port 358 nsew signal tristate
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 la_data_out[88]
port 359 nsew signal tristate
flabel metal2 s 41694 0 41750 800 0 FreeSans 224 90 0 0 la_data_out[89]
port 360 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 la_data_out[8]
port 361 nsew signal tristate
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 la_data_out[90]
port 362 nsew signal tristate
flabel metal2 s 42246 0 42302 800 0 FreeSans 224 90 0 0 la_data_out[91]
port 363 nsew signal tristate
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 la_data_out[92]
port 364 nsew signal tristate
flabel metal2 s 42798 0 42854 800 0 FreeSans 224 90 0 0 la_data_out[93]
port 365 nsew signal tristate
flabel metal2 s 43074 0 43130 800 0 FreeSans 224 90 0 0 la_data_out[94]
port 366 nsew signal tristate
flabel metal2 s 43350 0 43406 800 0 FreeSans 224 90 0 0 la_data_out[95]
port 367 nsew signal tristate
flabel metal2 s 43626 0 43682 800 0 FreeSans 224 90 0 0 la_data_out[96]
port 368 nsew signal tristate
flabel metal2 s 43902 0 43958 800 0 FreeSans 224 90 0 0 la_data_out[97]
port 369 nsew signal tristate
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 la_data_out[98]
port 370 nsew signal tristate
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 la_data_out[99]
port 371 nsew signal tristate
flabel metal2 s 19614 0 19670 800 0 FreeSans 224 90 0 0 la_data_out[9]
port 372 nsew signal tristate
flabel metal2 s 17222 0 17278 800 0 FreeSans 224 90 0 0 la_oenb[0]
port 373 nsew signal input
flabel metal2 s 44822 0 44878 800 0 FreeSans 224 90 0 0 la_oenb[100]
port 374 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 la_oenb[101]
port 375 nsew signal input
flabel metal2 s 45374 0 45430 800 0 FreeSans 224 90 0 0 la_oenb[102]
port 376 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 la_oenb[103]
port 377 nsew signal input
flabel metal2 s 45926 0 45982 800 0 FreeSans 224 90 0 0 la_oenb[104]
port 378 nsew signal input
flabel metal2 s 46202 0 46258 800 0 FreeSans 224 90 0 0 la_oenb[105]
port 379 nsew signal input
flabel metal2 s 46478 0 46534 800 0 FreeSans 224 90 0 0 la_oenb[106]
port 380 nsew signal input
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 la_oenb[107]
port 381 nsew signal input
flabel metal2 s 47030 0 47086 800 0 FreeSans 224 90 0 0 la_oenb[108]
port 382 nsew signal input
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 la_oenb[109]
port 383 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 la_oenb[10]
port 384 nsew signal input
flabel metal2 s 47582 0 47638 800 0 FreeSans 224 90 0 0 la_oenb[110]
port 385 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 la_oenb[111]
port 386 nsew signal input
flabel metal2 s 48134 0 48190 800 0 FreeSans 224 90 0 0 la_oenb[112]
port 387 nsew signal input
flabel metal2 s 48410 0 48466 800 0 FreeSans 224 90 0 0 la_oenb[113]
port 388 nsew signal input
flabel metal2 s 48686 0 48742 800 0 FreeSans 224 90 0 0 la_oenb[114]
port 389 nsew signal input
flabel metal2 s 48962 0 49018 800 0 FreeSans 224 90 0 0 la_oenb[115]
port 390 nsew signal input
flabel metal2 s 49238 0 49294 800 0 FreeSans 224 90 0 0 la_oenb[116]
port 391 nsew signal input
flabel metal2 s 49514 0 49570 800 0 FreeSans 224 90 0 0 la_oenb[117]
port 392 nsew signal input
flabel metal2 s 49790 0 49846 800 0 FreeSans 224 90 0 0 la_oenb[118]
port 393 nsew signal input
flabel metal2 s 50066 0 50122 800 0 FreeSans 224 90 0 0 la_oenb[119]
port 394 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 la_oenb[11]
port 395 nsew signal input
flabel metal2 s 50342 0 50398 800 0 FreeSans 224 90 0 0 la_oenb[120]
port 396 nsew signal input
flabel metal2 s 50618 0 50674 800 0 FreeSans 224 90 0 0 la_oenb[121]
port 397 nsew signal input
flabel metal2 s 50894 0 50950 800 0 FreeSans 224 90 0 0 la_oenb[122]
port 398 nsew signal input
flabel metal2 s 51170 0 51226 800 0 FreeSans 224 90 0 0 la_oenb[123]
port 399 nsew signal input
flabel metal2 s 51446 0 51502 800 0 FreeSans 224 90 0 0 la_oenb[124]
port 400 nsew signal input
flabel metal2 s 51722 0 51778 800 0 FreeSans 224 90 0 0 la_oenb[125]
port 401 nsew signal input
flabel metal2 s 51998 0 52054 800 0 FreeSans 224 90 0 0 la_oenb[126]
port 402 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 la_oenb[127]
port 403 nsew signal input
flabel metal2 s 20534 0 20590 800 0 FreeSans 224 90 0 0 la_oenb[12]
port 404 nsew signal input
flabel metal2 s 20810 0 20866 800 0 FreeSans 224 90 0 0 la_oenb[13]
port 405 nsew signal input
flabel metal2 s 21086 0 21142 800 0 FreeSans 224 90 0 0 la_oenb[14]
port 406 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 la_oenb[15]
port 407 nsew signal input
flabel metal2 s 21638 0 21694 800 0 FreeSans 224 90 0 0 la_oenb[16]
port 408 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 la_oenb[17]
port 409 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 la_oenb[18]
port 410 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 la_oenb[19]
port 411 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 la_oenb[1]
port 412 nsew signal input
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 la_oenb[20]
port 413 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 la_oenb[21]
port 414 nsew signal input
flabel metal2 s 23294 0 23350 800 0 FreeSans 224 90 0 0 la_oenb[22]
port 415 nsew signal input
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 la_oenb[23]
port 416 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 la_oenb[24]
port 417 nsew signal input
flabel metal2 s 24122 0 24178 800 0 FreeSans 224 90 0 0 la_oenb[25]
port 418 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 la_oenb[26]
port 419 nsew signal input
flabel metal2 s 24674 0 24730 800 0 FreeSans 224 90 0 0 la_oenb[27]
port 420 nsew signal input
flabel metal2 s 24950 0 25006 800 0 FreeSans 224 90 0 0 la_oenb[28]
port 421 nsew signal input
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 la_oenb[29]
port 422 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 la_oenb[2]
port 423 nsew signal input
flabel metal2 s 25502 0 25558 800 0 FreeSans 224 90 0 0 la_oenb[30]
port 424 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 la_oenb[31]
port 425 nsew signal input
flabel metal2 s 26054 0 26110 800 0 FreeSans 224 90 0 0 la_oenb[32]
port 426 nsew signal input
flabel metal2 s 26330 0 26386 800 0 FreeSans 224 90 0 0 la_oenb[33]
port 427 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 la_oenb[34]
port 428 nsew signal input
flabel metal2 s 26882 0 26938 800 0 FreeSans 224 90 0 0 la_oenb[35]
port 429 nsew signal input
flabel metal2 s 27158 0 27214 800 0 FreeSans 224 90 0 0 la_oenb[36]
port 430 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 la_oenb[37]
port 431 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 la_oenb[38]
port 432 nsew signal input
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 la_oenb[39]
port 433 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 la_oenb[3]
port 434 nsew signal input
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 la_oenb[40]
port 435 nsew signal input
flabel metal2 s 28538 0 28594 800 0 FreeSans 224 90 0 0 la_oenb[41]
port 436 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 la_oenb[42]
port 437 nsew signal input
flabel metal2 s 29090 0 29146 800 0 FreeSans 224 90 0 0 la_oenb[43]
port 438 nsew signal input
flabel metal2 s 29366 0 29422 800 0 FreeSans 224 90 0 0 la_oenb[44]
port 439 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 la_oenb[45]
port 440 nsew signal input
flabel metal2 s 29918 0 29974 800 0 FreeSans 224 90 0 0 la_oenb[46]
port 441 nsew signal input
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 la_oenb[47]
port 442 nsew signal input
flabel metal2 s 30470 0 30526 800 0 FreeSans 224 90 0 0 la_oenb[48]
port 443 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 la_oenb[49]
port 444 nsew signal input
flabel metal2 s 18326 0 18382 800 0 FreeSans 224 90 0 0 la_oenb[4]
port 445 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 la_oenb[50]
port 446 nsew signal input
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 la_oenb[51]
port 447 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 la_oenb[52]
port 448 nsew signal input
flabel metal2 s 31850 0 31906 800 0 FreeSans 224 90 0 0 la_oenb[53]
port 449 nsew signal input
flabel metal2 s 32126 0 32182 800 0 FreeSans 224 90 0 0 la_oenb[54]
port 450 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 la_oenb[55]
port 451 nsew signal input
flabel metal2 s 32678 0 32734 800 0 FreeSans 224 90 0 0 la_oenb[56]
port 452 nsew signal input
flabel metal2 s 32954 0 33010 800 0 FreeSans 224 90 0 0 la_oenb[57]
port 453 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 la_oenb[58]
port 454 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 la_oenb[59]
port 455 nsew signal input
flabel metal2 s 18602 0 18658 800 0 FreeSans 224 90 0 0 la_oenb[5]
port 456 nsew signal input
flabel metal2 s 33782 0 33838 800 0 FreeSans 224 90 0 0 la_oenb[60]
port 457 nsew signal input
flabel metal2 s 34058 0 34114 800 0 FreeSans 224 90 0 0 la_oenb[61]
port 458 nsew signal input
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 la_oenb[62]
port 459 nsew signal input
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 la_oenb[63]
port 460 nsew signal input
flabel metal2 s 34886 0 34942 800 0 FreeSans 224 90 0 0 la_oenb[64]
port 461 nsew signal input
flabel metal2 s 35162 0 35218 800 0 FreeSans 224 90 0 0 la_oenb[65]
port 462 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 la_oenb[66]
port 463 nsew signal input
flabel metal2 s 35714 0 35770 800 0 FreeSans 224 90 0 0 la_oenb[67]
port 464 nsew signal input
flabel metal2 s 35990 0 36046 800 0 FreeSans 224 90 0 0 la_oenb[68]
port 465 nsew signal input
flabel metal2 s 36266 0 36322 800 0 FreeSans 224 90 0 0 la_oenb[69]
port 466 nsew signal input
flabel metal2 s 18878 0 18934 800 0 FreeSans 224 90 0 0 la_oenb[6]
port 467 nsew signal input
flabel metal2 s 36542 0 36598 800 0 FreeSans 224 90 0 0 la_oenb[70]
port 468 nsew signal input
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 la_oenb[71]
port 469 nsew signal input
flabel metal2 s 37094 0 37150 800 0 FreeSans 224 90 0 0 la_oenb[72]
port 470 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 la_oenb[73]
port 471 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 la_oenb[74]
port 472 nsew signal input
flabel metal2 s 37922 0 37978 800 0 FreeSans 224 90 0 0 la_oenb[75]
port 473 nsew signal input
flabel metal2 s 38198 0 38254 800 0 FreeSans 224 90 0 0 la_oenb[76]
port 474 nsew signal input
flabel metal2 s 38474 0 38530 800 0 FreeSans 224 90 0 0 la_oenb[77]
port 475 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 la_oenb[78]
port 476 nsew signal input
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 la_oenb[79]
port 477 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 la_oenb[7]
port 478 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 la_oenb[80]
port 479 nsew signal input
flabel metal2 s 39578 0 39634 800 0 FreeSans 224 90 0 0 la_oenb[81]
port 480 nsew signal input
flabel metal2 s 39854 0 39910 800 0 FreeSans 224 90 0 0 la_oenb[82]
port 481 nsew signal input
flabel metal2 s 40130 0 40186 800 0 FreeSans 224 90 0 0 la_oenb[83]
port 482 nsew signal input
flabel metal2 s 40406 0 40462 800 0 FreeSans 224 90 0 0 la_oenb[84]
port 483 nsew signal input
flabel metal2 s 40682 0 40738 800 0 FreeSans 224 90 0 0 la_oenb[85]
port 484 nsew signal input
flabel metal2 s 40958 0 41014 800 0 FreeSans 224 90 0 0 la_oenb[86]
port 485 nsew signal input
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 la_oenb[87]
port 486 nsew signal input
flabel metal2 s 41510 0 41566 800 0 FreeSans 224 90 0 0 la_oenb[88]
port 487 nsew signal input
flabel metal2 s 41786 0 41842 800 0 FreeSans 224 90 0 0 la_oenb[89]
port 488 nsew signal input
flabel metal2 s 19430 0 19486 800 0 FreeSans 224 90 0 0 la_oenb[8]
port 489 nsew signal input
flabel metal2 s 42062 0 42118 800 0 FreeSans 224 90 0 0 la_oenb[90]
port 490 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 la_oenb[91]
port 491 nsew signal input
flabel metal2 s 42614 0 42670 800 0 FreeSans 224 90 0 0 la_oenb[92]
port 492 nsew signal input
flabel metal2 s 42890 0 42946 800 0 FreeSans 224 90 0 0 la_oenb[93]
port 493 nsew signal input
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 la_oenb[94]
port 494 nsew signal input
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 la_oenb[95]
port 495 nsew signal input
flabel metal2 s 43718 0 43774 800 0 FreeSans 224 90 0 0 la_oenb[96]
port 496 nsew signal input
flabel metal2 s 43994 0 44050 800 0 FreeSans 224 90 0 0 la_oenb[97]
port 497 nsew signal input
flabel metal2 s 44270 0 44326 800 0 FreeSans 224 90 0 0 la_oenb[98]
port 498 nsew signal input
flabel metal2 s 44546 0 44602 800 0 FreeSans 224 90 0 0 la_oenb[99]
port 499 nsew signal input
flabel metal2 s 19706 0 19762 800 0 FreeSans 224 90 0 0 la_oenb[9]
port 500 nsew signal input
flabel metal4 s 8168 2128 8488 7664 0 FreeSans 1920 90 0 0 vccd1
port 501 nsew power bidirectional
flabel metal4 s 22616 2128 22936 7664 0 FreeSans 1920 90 0 0 vccd1
port 501 nsew power bidirectional
flabel metal4 s 37064 2128 37384 7664 0 FreeSans 1920 90 0 0 vccd1
port 501 nsew power bidirectional
flabel metal4 s 51512 2128 51832 7664 0 FreeSans 1920 90 0 0 vccd1
port 501 nsew power bidirectional
flabel metal4 s 15392 2128 15712 7664 0 FreeSans 1920 90 0 0 vssd1
port 502 nsew ground bidirectional
flabel metal4 s 29840 2128 30160 7664 0 FreeSans 1920 90 0 0 vssd1
port 502 nsew ground bidirectional
flabel metal4 s 44288 2128 44608 7664 0 FreeSans 1920 90 0 0 vssd1
port 502 nsew ground bidirectional
flabel metal2 s 7286 0 7342 800 0 FreeSans 224 90 0 0 wb_clk_i
port 503 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 wb_rst_i
port 504 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wbs_ack_o
port 505 nsew signal tristate
flabel metal2 s 7838 0 7894 800 0 FreeSans 224 90 0 0 wbs_adr_i[0]
port 506 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wbs_adr_i[10]
port 507 nsew signal input
flabel metal2 s 11242 0 11298 800 0 FreeSans 224 90 0 0 wbs_adr_i[11]
port 508 nsew signal input
flabel metal2 s 11518 0 11574 800 0 FreeSans 224 90 0 0 wbs_adr_i[12]
port 509 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 wbs_adr_i[13]
port 510 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 wbs_adr_i[14]
port 511 nsew signal input
flabel metal2 s 12346 0 12402 800 0 FreeSans 224 90 0 0 wbs_adr_i[15]
port 512 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wbs_adr_i[16]
port 513 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 wbs_adr_i[17]
port 514 nsew signal input
flabel metal2 s 13174 0 13230 800 0 FreeSans 224 90 0 0 wbs_adr_i[18]
port 515 nsew signal input
flabel metal2 s 13450 0 13506 800 0 FreeSans 224 90 0 0 wbs_adr_i[19]
port 516 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wbs_adr_i[1]
port 517 nsew signal input
flabel metal2 s 13726 0 13782 800 0 FreeSans 224 90 0 0 wbs_adr_i[20]
port 518 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 wbs_adr_i[21]
port 519 nsew signal input
flabel metal2 s 14278 0 14334 800 0 FreeSans 224 90 0 0 wbs_adr_i[22]
port 520 nsew signal input
flabel metal2 s 14554 0 14610 800 0 FreeSans 224 90 0 0 wbs_adr_i[23]
port 521 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wbs_adr_i[24]
port 522 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 wbs_adr_i[25]
port 523 nsew signal input
flabel metal2 s 15382 0 15438 800 0 FreeSans 224 90 0 0 wbs_adr_i[26]
port 524 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 wbs_adr_i[27]
port 525 nsew signal input
flabel metal2 s 15934 0 15990 800 0 FreeSans 224 90 0 0 wbs_adr_i[28]
port 526 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 wbs_adr_i[29]
port 527 nsew signal input
flabel metal2 s 8574 0 8630 800 0 FreeSans 224 90 0 0 wbs_adr_i[2]
port 528 nsew signal input
flabel metal2 s 16486 0 16542 800 0 FreeSans 224 90 0 0 wbs_adr_i[30]
port 529 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wbs_adr_i[31]
port 530 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wbs_adr_i[3]
port 531 nsew signal input
flabel metal2 s 9310 0 9366 800 0 FreeSans 224 90 0 0 wbs_adr_i[4]
port 532 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 wbs_adr_i[5]
port 533 nsew signal input
flabel metal2 s 9862 0 9918 800 0 FreeSans 224 90 0 0 wbs_adr_i[6]
port 534 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 wbs_adr_i[7]
port 535 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wbs_adr_i[8]
port 536 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 wbs_adr_i[9]
port 537 nsew signal input
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 wbs_cyc_i
port 538 nsew signal input
flabel metal2 s 7930 0 7986 800 0 FreeSans 224 90 0 0 wbs_dat_i[0]
port 539 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 wbs_dat_i[10]
port 540 nsew signal input
flabel metal2 s 11334 0 11390 800 0 FreeSans 224 90 0 0 wbs_dat_i[11]
port 541 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 wbs_dat_i[12]
port 542 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wbs_dat_i[13]
port 543 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 wbs_dat_i[14]
port 544 nsew signal input
flabel metal2 s 12438 0 12494 800 0 FreeSans 224 90 0 0 wbs_dat_i[15]
port 545 nsew signal input
flabel metal2 s 12714 0 12770 800 0 FreeSans 224 90 0 0 wbs_dat_i[16]
port 546 nsew signal input
flabel metal2 s 12990 0 13046 800 0 FreeSans 224 90 0 0 wbs_dat_i[17]
port 547 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 wbs_dat_i[18]
port 548 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wbs_dat_i[19]
port 549 nsew signal input
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 wbs_dat_i[1]
port 550 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 wbs_dat_i[20]
port 551 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wbs_dat_i[21]
port 552 nsew signal input
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 wbs_dat_i[22]
port 553 nsew signal input
flabel metal2 s 14646 0 14702 800 0 FreeSans 224 90 0 0 wbs_dat_i[23]
port 554 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wbs_dat_i[24]
port 555 nsew signal input
flabel metal2 s 15198 0 15254 800 0 FreeSans 224 90 0 0 wbs_dat_i[25]
port 556 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 wbs_dat_i[26]
port 557 nsew signal input
flabel metal2 s 15750 0 15806 800 0 FreeSans 224 90 0 0 wbs_dat_i[27]
port 558 nsew signal input
flabel metal2 s 16026 0 16082 800 0 FreeSans 224 90 0 0 wbs_dat_i[28]
port 559 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wbs_dat_i[29]
port 560 nsew signal input
flabel metal2 s 8666 0 8722 800 0 FreeSans 224 90 0 0 wbs_dat_i[2]
port 561 nsew signal input
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 wbs_dat_i[30]
port 562 nsew signal input
flabel metal2 s 16854 0 16910 800 0 FreeSans 224 90 0 0 wbs_dat_i[31]
port 563 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wbs_dat_i[3]
port 564 nsew signal input
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 wbs_dat_i[4]
port 565 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wbs_dat_i[5]
port 566 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 wbs_dat_i[6]
port 567 nsew signal input
flabel metal2 s 10230 0 10286 800 0 FreeSans 224 90 0 0 wbs_dat_i[7]
port 568 nsew signal input
flabel metal2 s 10506 0 10562 800 0 FreeSans 224 90 0 0 wbs_dat_i[8]
port 569 nsew signal input
flabel metal2 s 10782 0 10838 800 0 FreeSans 224 90 0 0 wbs_dat_i[9]
port 570 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 wbs_dat_o[0]
port 571 nsew signal tristate
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wbs_dat_o[10]
port 572 nsew signal tristate
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 wbs_dat_o[11]
port 573 nsew signal tristate
flabel metal2 s 11702 0 11758 800 0 FreeSans 224 90 0 0 wbs_dat_o[12]
port 574 nsew signal tristate
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 wbs_dat_o[13]
port 575 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wbs_dat_o[14]
port 576 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 wbs_dat_o[15]
port 577 nsew signal tristate
flabel metal2 s 12806 0 12862 800 0 FreeSans 224 90 0 0 wbs_dat_o[16]
port 578 nsew signal tristate
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 wbs_dat_o[17]
port 579 nsew signal tristate
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wbs_dat_o[18]
port 580 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 wbs_dat_o[19]
port 581 nsew signal tristate
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 wbs_dat_o[1]
port 582 nsew signal tristate
flabel metal2 s 13910 0 13966 800 0 FreeSans 224 90 0 0 wbs_dat_o[20]
port 583 nsew signal tristate
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 wbs_dat_o[21]
port 584 nsew signal tristate
flabel metal2 s 14462 0 14518 800 0 FreeSans 224 90 0 0 wbs_dat_o[22]
port 585 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 wbs_dat_o[23]
port 586 nsew signal tristate
flabel metal2 s 15014 0 15070 800 0 FreeSans 224 90 0 0 wbs_dat_o[24]
port 587 nsew signal tristate
flabel metal2 s 15290 0 15346 800 0 FreeSans 224 90 0 0 wbs_dat_o[25]
port 588 nsew signal tristate
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wbs_dat_o[26]
port 589 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 wbs_dat_o[27]
port 590 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wbs_dat_o[28]
port 591 nsew signal tristate
flabel metal2 s 16394 0 16450 800 0 FreeSans 224 90 0 0 wbs_dat_o[29]
port 592 nsew signal tristate
flabel metal2 s 8758 0 8814 800 0 FreeSans 224 90 0 0 wbs_dat_o[2]
port 593 nsew signal tristate
flabel metal2 s 16670 0 16726 800 0 FreeSans 224 90 0 0 wbs_dat_o[30]
port 594 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 wbs_dat_o[31]
port 595 nsew signal tristate
flabel metal2 s 9126 0 9182 800 0 FreeSans 224 90 0 0 wbs_dat_o[3]
port 596 nsew signal tristate
flabel metal2 s 9494 0 9550 800 0 FreeSans 224 90 0 0 wbs_dat_o[4]
port 597 nsew signal tristate
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 wbs_dat_o[5]
port 598 nsew signal tristate
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 wbs_dat_o[6]
port 599 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wbs_dat_o[7]
port 600 nsew signal tristate
flabel metal2 s 10598 0 10654 800 0 FreeSans 224 90 0 0 wbs_dat_o[8]
port 601 nsew signal tristate
flabel metal2 s 10874 0 10930 800 0 FreeSans 224 90 0 0 wbs_dat_o[9]
port 602 nsew signal tristate
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 wbs_sel_i[0]
port 603 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 wbs_sel_i[1]
port 604 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 wbs_sel_i[2]
port 605 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 wbs_sel_i[3]
port 606 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 wbs_stb_i
port 607 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wbs_we_i
port 608 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 10000
<< end >>
